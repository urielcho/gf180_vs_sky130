* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for Top_Module_4_ALU abstract view
.subckt Top_Module_4_ALU ALU_Output[0] ALU_Output[100] ALU_Output[101] ALU_Output[102]
+ ALU_Output[103] ALU_Output[104] ALU_Output[105] ALU_Output[106] ALU_Output[107]
+ ALU_Output[108] ALU_Output[109] ALU_Output[10] ALU_Output[110] ALU_Output[111] ALU_Output[112]
+ ALU_Output[113] ALU_Output[114] ALU_Output[115] ALU_Output[116] ALU_Output[117]
+ ALU_Output[118] ALU_Output[119] ALU_Output[11] ALU_Output[120] ALU_Output[121] ALU_Output[122]
+ ALU_Output[123] ALU_Output[124] ALU_Output[125] ALU_Output[126] ALU_Output[127]
+ ALU_Output[12] ALU_Output[13] ALU_Output[14] ALU_Output[15] ALU_Output[16] ALU_Output[17]
+ ALU_Output[18] ALU_Output[19] ALU_Output[1] ALU_Output[20] ALU_Output[21] ALU_Output[22]
+ ALU_Output[23] ALU_Output[24] ALU_Output[25] ALU_Output[26] ALU_Output[27] ALU_Output[28]
+ ALU_Output[29] ALU_Output[2] ALU_Output[30] ALU_Output[31] ALU_Output[32] ALU_Output[33]
+ ALU_Output[34] ALU_Output[35] ALU_Output[36] ALU_Output[37] ALU_Output[38] ALU_Output[39]
+ ALU_Output[3] ALU_Output[40] ALU_Output[41] ALU_Output[42] ALU_Output[43] ALU_Output[44]
+ ALU_Output[45] ALU_Output[46] ALU_Output[47] ALU_Output[48] ALU_Output[49] ALU_Output[4]
+ ALU_Output[50] ALU_Output[51] ALU_Output[52] ALU_Output[53] ALU_Output[54] ALU_Output[55]
+ ALU_Output[56] ALU_Output[57] ALU_Output[58] ALU_Output[59] ALU_Output[5] ALU_Output[60]
+ ALU_Output[61] ALU_Output[62] ALU_Output[63] ALU_Output[64] ALU_Output[65] ALU_Output[66]
+ ALU_Output[67] ALU_Output[68] ALU_Output[69] ALU_Output[6] ALU_Output[70] ALU_Output[71]
+ ALU_Output[72] ALU_Output[73] ALU_Output[74] ALU_Output[75] ALU_Output[76] ALU_Output[77]
+ ALU_Output[78] ALU_Output[79] ALU_Output[7] ALU_Output[80] ALU_Output[81] ALU_Output[82]
+ ALU_Output[83] ALU_Output[84] ALU_Output[85] ALU_Output[86] ALU_Output[87] ALU_Output[88]
+ ALU_Output[89] ALU_Output[8] ALU_Output[90] ALU_Output[91] ALU_Output[92] ALU_Output[93]
+ ALU_Output[94] ALU_Output[95] ALU_Output[96] ALU_Output[97] ALU_Output[98] ALU_Output[99]
+ ALU_Output[9] Exception[0] Exception[1] Exception[2] Exception[3] Operation[0] Operation[1]
+ Operation[2] Operation[3] Overflow[0] Overflow[1] Overflow[2] Overflow[3] Underflow[0]
+ Underflow[1] Underflow[2] Underflow[3] a_operand[0] a_operand[100] a_operand[101]
+ a_operand[102] a_operand[103] a_operand[104] a_operand[105] a_operand[106] a_operand[107]
+ a_operand[108] a_operand[109] a_operand[10] a_operand[110] a_operand[111] a_operand[112]
+ a_operand[113] a_operand[114] a_operand[115] a_operand[116] a_operand[117] a_operand[118]
+ a_operand[119] a_operand[11] a_operand[120] a_operand[121] a_operand[122] a_operand[123]
+ a_operand[124] a_operand[125] a_operand[126] a_operand[127] a_operand[12] a_operand[13]
+ a_operand[14] a_operand[15] a_operand[16] a_operand[17] a_operand[18] a_operand[19]
+ a_operand[1] a_operand[20] a_operand[21] a_operand[22] a_operand[23] a_operand[24]
+ a_operand[25] a_operand[26] a_operand[27] a_operand[28] a_operand[29] a_operand[2]
+ a_operand[30] a_operand[31] a_operand[32] a_operand[33] a_operand[34] a_operand[35]
+ a_operand[36] a_operand[37] a_operand[38] a_operand[39] a_operand[3] a_operand[40]
+ a_operand[41] a_operand[42] a_operand[43] a_operand[44] a_operand[45] a_operand[46]
+ a_operand[47] a_operand[48] a_operand[49] a_operand[4] a_operand[50] a_operand[51]
+ a_operand[52] a_operand[53] a_operand[54] a_operand[55] a_operand[56] a_operand[57]
+ a_operand[58] a_operand[59] a_operand[5] a_operand[60] a_operand[61] a_operand[62]
+ a_operand[63] a_operand[64] a_operand[65] a_operand[66] a_operand[67] a_operand[68]
+ a_operand[69] a_operand[6] a_operand[70] a_operand[71] a_operand[72] a_operand[73]
+ a_operand[74] a_operand[75] a_operand[76] a_operand[77] a_operand[78] a_operand[79]
+ a_operand[7] a_operand[80] a_operand[81] a_operand[82] a_operand[83] a_operand[84]
+ a_operand[85] a_operand[86] a_operand[87] a_operand[88] a_operand[89] a_operand[8]
+ a_operand[90] a_operand[91] a_operand[92] a_operand[93] a_operand[94] a_operand[95]
+ a_operand[96] a_operand[97] a_operand[98] a_operand[99] a_operand[9] b_operand[0]
+ b_operand[100] b_operand[101] b_operand[102] b_operand[103] b_operand[104] b_operand[105]
+ b_operand[106] b_operand[107] b_operand[108] b_operand[109] b_operand[10] b_operand[110]
+ b_operand[111] b_operand[112] b_operand[113] b_operand[114] b_operand[115] b_operand[116]
+ b_operand[117] b_operand[118] b_operand[119] b_operand[11] b_operand[120] b_operand[121]
+ b_operand[122] b_operand[123] b_operand[124] b_operand[125] b_operand[126] b_operand[127]
+ b_operand[12] b_operand[13] b_operand[14] b_operand[15] b_operand[16] b_operand[17]
+ b_operand[18] b_operand[19] b_operand[1] b_operand[20] b_operand[21] b_operand[22]
+ b_operand[23] b_operand[24] b_operand[25] b_operand[26] b_operand[27] b_operand[28]
+ b_operand[29] b_operand[2] b_operand[30] b_operand[31] b_operand[32] b_operand[33]
+ b_operand[34] b_operand[35] b_operand[36] b_operand[37] b_operand[38] b_operand[39]
+ b_operand[3] b_operand[40] b_operand[41] b_operand[42] b_operand[43] b_operand[44]
+ b_operand[45] b_operand[46] b_operand[47] b_operand[48] b_operand[49] b_operand[4]
+ b_operand[50] b_operand[51] b_operand[52] b_operand[53] b_operand[54] b_operand[55]
+ b_operand[56] b_operand[57] b_operand[58] b_operand[59] b_operand[5] b_operand[60]
+ b_operand[61] b_operand[62] b_operand[63] b_operand[64] b_operand[65] b_operand[66]
+ b_operand[67] b_operand[68] b_operand[69] b_operand[6] b_operand[70] b_operand[71]
+ b_operand[72] b_operand[73] b_operand[74] b_operand[75] b_operand[76] b_operand[77]
+ b_operand[78] b_operand[79] b_operand[7] b_operand[80] b_operand[81] b_operand[82]
+ b_operand[83] b_operand[84] b_operand[85] b_operand[86] b_operand[87] b_operand[88]
+ b_operand[89] b_operand[8] b_operand[90] b_operand[91] b_operand[92] b_operand[93]
+ b_operand[94] b_operand[95] b_operand[96] b_operand[97] b_operand[98] b_operand[99]
+ b_operand[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for OQPSK_PS_RCOSINE2 abstract view
.subckt OQPSK_PS_RCOSINE2 BitIn CLK EN I[0] I[10] I[11] I[12] I[1] I[2] I[3] I[4]
+ I[5] I[6] I[7] I[8] I[9] Q[0] Q[10] Q[11] Q[12] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] RST addI[0] addI[1] addI[2] addI[3] addI[4] addI[5] addQ[0] addQ[1] addQ[2]
+ addQ[3] addQ[4] addQ[5] vccd1 vssd1
.ends

* Black-box entry subcircuit for OQPSK_RCOSINE_ALL abstract view
.subckt OQPSK_RCOSINE_ALL ACK Bit_In EN I[0] I[10] I[11] I[12] I[1] I[2] I[3] I[4]
+ I[5] I[6] I[7] I[8] I[9] Q[0] Q[10] Q[11] Q[12] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] REQ_SAMPLE RST addI[0] addI[1] addI[2] addI[3] addI[4] addI[5] addQ[0]
+ addQ[1] addQ[2] addQ[3] addQ[4] addQ[5] vccd1 vssd1
.ends

* Black-box entry subcircuit for divider abstract view
.subckt divider clk cout1 cout10 cout2 cout3 cout4 cout5 cout6 cout7 cout8 cout9 vccd1
+ vssd1
.ends

* Black-box entry subcircuit for posoco2000 abstract view
.subckt posoco2000 clk segm[0] segm[1] segm[2] segm[3] segm[4] segm[5] segm[6] segm[7]
+ sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XTop_Module_4_ALU la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] Top_Module_4_ALU/Exception[0] Top_Module_4_ALU/Exception[1] Top_Module_4_ALU/Exception[2]
+ Top_Module_4_ALU/Exception[3] io_in[5] io_in[6] io_in[7] io_in[8] Top_Module_4_ALU/Overflow[0]
+ Top_Module_4_ALU/Overflow[1] Top_Module_4_ALU/Overflow[2] Top_Module_4_ALU/Overflow[3]
+ Top_Module_4_ALU/Underflow[0] Top_Module_4_ALU/Underflow[1] Top_Module_4_ALU/Underflow[2]
+ Top_Module_4_ALU/Underflow[3] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 Top_Module_4_ALU
XOQPSK_PS_RCOSINE2 OQPSK_PS_RCOSINE2/BitIn OQPSK_PS_RCOSINE2/CLK OQPSK_PS_RCOSINE2/EN
+ OQPSK_PS_RCOSINE2/I[0] OQPSK_PS_RCOSINE2/I[10] OQPSK_PS_RCOSINE2/I[11] OQPSK_PS_RCOSINE2/I[12]
+ OQPSK_PS_RCOSINE2/I[1] OQPSK_PS_RCOSINE2/I[2] OQPSK_PS_RCOSINE2/I[3] OQPSK_PS_RCOSINE2/I[4]
+ OQPSK_PS_RCOSINE2/I[5] OQPSK_PS_RCOSINE2/I[6] OQPSK_PS_RCOSINE2/I[7] OQPSK_PS_RCOSINE2/I[8]
+ OQPSK_PS_RCOSINE2/I[9] OQPSK_PS_RCOSINE2/Q[0] OQPSK_PS_RCOSINE2/Q[10] OQPSK_PS_RCOSINE2/Q[11]
+ OQPSK_PS_RCOSINE2/Q[12] OQPSK_PS_RCOSINE2/Q[1] OQPSK_PS_RCOSINE2/Q[2] OQPSK_PS_RCOSINE2/Q[3]
+ OQPSK_PS_RCOSINE2/Q[4] OQPSK_PS_RCOSINE2/Q[5] OQPSK_PS_RCOSINE2/Q[6] OQPSK_PS_RCOSINE2/Q[7]
+ OQPSK_PS_RCOSINE2/Q[8] OQPSK_PS_RCOSINE2/Q[9] OQPSK_PS_RCOSINE2/RST OQPSK_PS_RCOSINE2/addI[0]
+ OQPSK_PS_RCOSINE2/addI[1] OQPSK_PS_RCOSINE2/addI[2] OQPSK_PS_RCOSINE2/addI[3] OQPSK_PS_RCOSINE2/addI[4]
+ OQPSK_PS_RCOSINE2/addI[5] OQPSK_PS_RCOSINE2/addQ[0] OQPSK_PS_RCOSINE2/addQ[1] OQPSK_PS_RCOSINE2/addQ[2]
+ OQPSK_PS_RCOSINE2/addQ[3] OQPSK_PS_RCOSINE2/addQ[4] OQPSK_PS_RCOSINE2/addQ[5] vccd1
+ vssd1 OQPSK_PS_RCOSINE2
XOQPSK_RCOSINE_ALL OQPSK_RCOSINE_ALL/ACK OQPSK_RCOSINE_ALL/Bit_In OQPSK_RCOSINE_ALL/EN
+ OQPSK_RCOSINE_ALL/I[0] OQPSK_RCOSINE_ALL/I[10] OQPSK_RCOSINE_ALL/I[11] OQPSK_RCOSINE_ALL/I[12]
+ OQPSK_RCOSINE_ALL/I[1] OQPSK_RCOSINE_ALL/I[2] OQPSK_RCOSINE_ALL/I[3] OQPSK_RCOSINE_ALL/I[4]
+ OQPSK_RCOSINE_ALL/I[5] OQPSK_RCOSINE_ALL/I[6] OQPSK_RCOSINE_ALL/I[7] OQPSK_RCOSINE_ALL/I[8]
+ OQPSK_RCOSINE_ALL/I[9] OQPSK_RCOSINE_ALL/Q[0] OQPSK_RCOSINE_ALL/Q[10] OQPSK_RCOSINE_ALL/Q[11]
+ OQPSK_RCOSINE_ALL/Q[12] OQPSK_RCOSINE_ALL/Q[1] OQPSK_RCOSINE_ALL/Q[2] OQPSK_RCOSINE_ALL/Q[3]
+ OQPSK_RCOSINE_ALL/Q[4] OQPSK_RCOSINE_ALL/Q[5] OQPSK_RCOSINE_ALL/Q[6] OQPSK_RCOSINE_ALL/Q[7]
+ OQPSK_RCOSINE_ALL/Q[8] OQPSK_RCOSINE_ALL/Q[9] OQPSK_RCOSINE_ALL/REQ_SAMPLE OQPSK_RCOSINE_ALL/RST
+ OQPSK_RCOSINE_ALL/addI[0] OQPSK_RCOSINE_ALL/addI[1] OQPSK_RCOSINE_ALL/addI[2] OQPSK_RCOSINE_ALL/addI[3]
+ OQPSK_RCOSINE_ALL/addI[4] OQPSK_RCOSINE_ALL/addI[5] OQPSK_RCOSINE_ALL/addQ[0] OQPSK_RCOSINE_ALL/addQ[1]
+ OQPSK_RCOSINE_ALL/addQ[2] OQPSK_RCOSINE_ALL/addQ[3] OQPSK_RCOSINE_ALL/addQ[4] OQPSK_RCOSINE_ALL/addQ[5]
+ vccd1 vssd1 OQPSK_RCOSINE_ALL
Xdivider wb_clk_i io_out[10] io_out[19] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] vccd1 vssd1 divider
Xposoco2000 wb_clk_i io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] vccd1 vssd1 posoco2000
.ends

