VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OQPSK_PS_RCOSINE2
  CLASS BLOCK ;
  FOREIGN OQPSK_PS_RCOSINE2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN BitIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 88.440 4.000 89.040 ;
    END
  END BitIn
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1.000 222.550 4.000 ;
    END
  END CLK
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 296.000 161.370 299.000 ;
    END
  END EN
  PIN I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 234.640 4.000 235.240 ;
    END
  END I[0]
  PIN I[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1.000 280.510 4.000 ;
    END
  END I[10]
  PIN I[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 3.440 299.000 4.040 ;
    END
  END I[11]
  PIN I[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 183.640 299.000 184.240 ;
    END
  END I[12]
  PIN I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 296.000 19.690 299.000 ;
    END
  END I[1]
  PIN I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 265.240 4.000 265.840 ;
    END
  END I[2]
  PIN I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 296.000 245.090 299.000 ;
    END
  END I[3]
  PIN I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1.000 167.810 4.000 ;
    END
  END I[4]
  PIN I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.840 299.000 211.440 ;
    END
  END I[5]
  PIN I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 299.000 34.640 ;
    END
  END I[6]
  PIN I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1.000 55.110 4.000 ;
    END
  END I[7]
  PIN I[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 204.040 4.000 204.640 ;
    END
  END I[8]
  PIN I[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 146.240 4.000 146.840 ;
    END
  END I[9]
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 296.000 190.350 299.000 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 296.000 274.070 299.000 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 176.840 4.000 177.440 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.440 299.000 242.040 ;
    END
  END Q[12]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 296.000 77.650 299.000 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 57.840 4.000 58.440 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 153.040 299.000 153.640 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 296.000 48.670 299.000 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 27.240 4.000 27.840 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1.000 251.530 4.000 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 296.000 216.110 299.000 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.640 299.000 65.240 ;
    END
  END Q[9]
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1.000 26.130 4.000 ;
    END
  END RST
  PIN addI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 1.000 84.090 4.000 ;
    END
  END addI[0]
  PIN addI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1.000 109.850 4.000 ;
    END
  END addI[1]
  PIN addI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.840 299.000 92.440 ;
    END
  END addI[2]
  PIN addI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1.000 138.830 4.000 ;
    END
  END addI[3]
  PIN addI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.040 299.000 272.640 ;
    END
  END addI[4]
  PIN addI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 299.240 299.000 299.840 ;
    END
  END addI[5]
  PIN addQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 296.000 106.630 299.000 ;
    END
  END addQ[0]
  PIN addQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 296.000 132.390 299.000 ;
    END
  END addQ[1]
  PIN addQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1.000 193.570 4.000 ;
    END
  END addQ[2]
  PIN addQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 115.640 4.000 116.240 ;
    END
  END addQ[3]
  PIN addQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 295.840 4.000 296.440 ;
    END
  END addQ[4]
  PIN addQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 299.000 123.040 ;
    END
  END addQ[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 0.070 9.900 299.850 288.560 ;
      LAYER met2 ;
        RECT 0.100 299.280 299.830 299.725 ;
        RECT 0.100 295.720 19.130 299.280 ;
        RECT 19.970 295.720 48.110 299.280 ;
        RECT 48.950 295.720 77.090 299.280 ;
        RECT 77.930 295.720 106.070 299.280 ;
        RECT 106.910 295.720 131.830 299.280 ;
        RECT 132.670 295.720 160.810 299.280 ;
        RECT 161.650 295.720 189.790 299.280 ;
        RECT 190.630 295.720 215.550 299.280 ;
        RECT 216.390 295.720 244.530 299.280 ;
        RECT 245.370 295.720 273.510 299.280 ;
        RECT 274.350 295.720 299.830 299.280 ;
        RECT 0.100 4.280 299.830 295.720 ;
        RECT 0.650 3.555 25.570 4.280 ;
        RECT 26.410 3.555 54.550 4.280 ;
        RECT 55.390 3.555 83.530 4.280 ;
        RECT 84.370 3.555 109.290 4.280 ;
        RECT 110.130 3.555 138.270 4.280 ;
        RECT 139.110 3.555 167.250 4.280 ;
        RECT 168.090 3.555 193.010 4.280 ;
        RECT 193.850 3.555 221.990 4.280 ;
        RECT 222.830 3.555 250.970 4.280 ;
        RECT 251.810 3.555 279.950 4.280 ;
        RECT 280.790 3.555 299.830 4.280 ;
      LAYER met3 ;
        RECT 4.000 298.840 295.600 299.705 ;
        RECT 299.400 298.840 299.855 299.705 ;
        RECT 4.000 296.840 299.855 298.840 ;
        RECT 4.400 295.440 299.855 296.840 ;
        RECT 4.000 273.040 299.855 295.440 ;
        RECT 4.000 271.640 295.600 273.040 ;
        RECT 299.400 271.640 299.855 273.040 ;
        RECT 4.000 266.240 299.855 271.640 ;
        RECT 4.400 264.840 299.855 266.240 ;
        RECT 4.000 242.440 299.855 264.840 ;
        RECT 4.000 241.040 295.600 242.440 ;
        RECT 299.400 241.040 299.855 242.440 ;
        RECT 4.000 235.640 299.855 241.040 ;
        RECT 4.400 234.240 299.855 235.640 ;
        RECT 4.000 211.840 299.855 234.240 ;
        RECT 4.000 210.440 295.600 211.840 ;
        RECT 299.400 210.440 299.855 211.840 ;
        RECT 4.000 205.040 299.855 210.440 ;
        RECT 4.400 203.640 299.855 205.040 ;
        RECT 4.000 184.640 299.855 203.640 ;
        RECT 4.000 183.240 295.600 184.640 ;
        RECT 299.400 183.240 299.855 184.640 ;
        RECT 4.000 177.840 299.855 183.240 ;
        RECT 4.400 176.440 299.855 177.840 ;
        RECT 4.000 154.040 299.855 176.440 ;
        RECT 4.000 152.640 295.600 154.040 ;
        RECT 299.400 152.640 299.855 154.040 ;
        RECT 4.000 147.240 299.855 152.640 ;
        RECT 4.400 145.840 299.855 147.240 ;
        RECT 4.000 123.440 299.855 145.840 ;
        RECT 4.000 122.040 295.600 123.440 ;
        RECT 299.400 122.040 299.855 123.440 ;
        RECT 4.000 116.640 299.855 122.040 ;
        RECT 4.400 115.240 299.855 116.640 ;
        RECT 4.000 92.840 299.855 115.240 ;
        RECT 4.000 91.440 295.600 92.840 ;
        RECT 299.400 91.440 299.855 92.840 ;
        RECT 4.000 89.440 299.855 91.440 ;
        RECT 4.400 88.040 299.855 89.440 ;
        RECT 4.000 65.640 299.855 88.040 ;
        RECT 4.000 64.240 295.600 65.640 ;
        RECT 299.400 64.240 299.855 65.640 ;
        RECT 4.000 58.840 299.855 64.240 ;
        RECT 4.400 57.440 299.855 58.840 ;
        RECT 4.000 35.040 299.855 57.440 ;
        RECT 4.000 33.640 295.600 35.040 ;
        RECT 299.400 33.640 299.855 35.040 ;
        RECT 4.000 28.240 299.855 33.640 ;
        RECT 4.400 26.840 299.855 28.240 ;
        RECT 4.000 4.440 299.855 26.840 ;
        RECT 4.000 3.575 295.600 4.440 ;
        RECT 299.400 3.575 299.855 4.440 ;
      LAYER met4 ;
        RECT 133.695 13.095 174.240 286.105 ;
        RECT 176.640 13.095 251.040 286.105 ;
        RECT 253.440 13.095 275.705 286.105 ;
  END
END OQPSK_PS_RCOSINE2
END LIBRARY

