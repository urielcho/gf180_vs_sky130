magic
tech sky130A
magscale 1 2
timestamp 1671750862
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 14 2128 58880 57712
<< metal2 >>
rect 4526 59200 4582 59800
rect 16762 59200 16818 59800
rect 28998 59200 29054 59800
rect 41878 59200 41934 59800
rect 54114 59200 54170 59800
rect 18 200 74 800
rect 12254 200 12310 800
rect 24490 200 24546 800
rect 36726 200 36782 800
rect 49606 200 49662 800
<< obsm2 >>
rect 20 59144 4470 59200
rect 4638 59144 16706 59200
rect 16874 59144 28942 59200
rect 29110 59144 41822 59200
rect 41990 59144 54058 59200
rect 54226 59144 58402 59200
rect 20 856 58402 59144
rect 130 800 12198 856
rect 12366 800 24434 856
rect 24602 800 36670 856
rect 36838 800 49550 856
rect 49718 800 58402 856
<< metal3 >>
rect 59200 53728 59800 53848
rect 200 52368 800 52488
rect 59200 40808 59800 40928
rect 200 38768 800 38888
rect 59200 27208 59800 27328
rect 200 25848 800 25968
rect 59200 14288 59800 14408
rect 200 12928 800 13048
rect 59200 1368 59800 1488
<< obsm3 >>
rect 800 53928 59200 57697
rect 800 53648 59120 53928
rect 800 52568 59200 53648
rect 880 52288 59200 52568
rect 800 41008 59200 52288
rect 800 40728 59120 41008
rect 800 38968 59200 40728
rect 880 38688 59200 38968
rect 800 27408 59200 38688
rect 800 27128 59120 27408
rect 800 26048 59200 27128
rect 880 25768 59200 26048
rect 800 14488 59200 25768
rect 800 14208 59120 14488
rect 800 13128 59200 14208
rect 880 12848 59200 13128
rect 800 1568 59200 12848
rect 800 1395 59120 1568
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal3 s 59200 1368 59800 1488 6 clk
port 1 nsew signal input
rlabel metal3 s 59200 14288 59800 14408 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 36726 200 36782 800 6 segm[1]
port 3 nsew signal output
rlabel metal3 s 59200 40808 59800 40928 6 segm[2]
port 4 nsew signal output
rlabel metal3 s 59200 53728 59800 53848 6 segm[3]
port 5 nsew signal output
rlabel metal3 s 200 52368 800 52488 6 segm[4]
port 6 nsew signal output
rlabel metal2 s 41878 59200 41934 59800 6 segm[5]
port 7 nsew signal output
rlabel metal2 s 18 200 74 800 6 segm[6]
port 8 nsew signal output
rlabel metal2 s 16762 59200 16818 59800 6 segm[7]
port 9 nsew signal output
rlabel metal2 s 49606 200 49662 800 6 sel[0]
port 10 nsew signal output
rlabel metal2 s 12254 200 12310 800 6 sel[1]
port 11 nsew signal output
rlabel metal2 s 28998 59200 29054 59800 6 sel[2]
port 12 nsew signal output
rlabel metal3 s 200 12928 800 13048 6 sel[3]
port 13 nsew signal output
rlabel metal3 s 200 25848 800 25968 6 sel[4]
port 14 nsew signal output
rlabel metal2 s 54114 59200 54170 59800 6 sel[5]
port 15 nsew signal output
rlabel metal2 s 24490 200 24546 800 6 sel[6]
port 16 nsew signal output
rlabel metal3 s 200 38768 800 38888 6 sel[7]
port 17 nsew signal output
rlabel metal2 s 4526 59200 4582 59800 6 sel[8]
port 18 nsew signal output
rlabel metal3 s 59200 27208 59800 27328 6 sel[9]
port 19 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 20 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 20 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 21 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 21 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1376900
string GDS_FILE /home/urielcho/Proyectos_caravel/MPW8/gf180_vs_sky130/openlane/posoco2000/runs/22_12_22_17_13/results/signoff/posoco2000.magic.gds
string GDS_START 263486
<< end >>

