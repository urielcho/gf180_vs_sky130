magic
tech sky130A
magscale 1 2
timestamp 1671750299
<< viali >>
rect 6653 57545 6687 57579
rect 28549 57545 28583 57579
rect 50537 57545 50571 57579
rect 6837 57409 6871 57443
rect 28733 57409 28767 57443
rect 50353 57409 50387 57443
rect 58081 49181 58115 49215
rect 58265 49045 58299 49079
rect 6653 46121 6687 46155
rect 46581 46121 46615 46155
rect 5273 45917 5307 45951
rect 40509 45917 40543 45951
rect 45201 45917 45235 45951
rect 5540 45849 5574 45883
rect 45468 45849 45502 45883
rect 5825 45577 5859 45611
rect 8861 45577 8895 45611
rect 9505 45509 9539 45543
rect 40408 45509 40442 45543
rect 6009 45441 6043 45475
rect 6745 45441 6779 45475
rect 7748 45441 7782 45475
rect 9689 45441 9723 45475
rect 27169 45441 27203 45475
rect 27425 45441 27459 45475
rect 44189 45441 44223 45475
rect 44456 45441 44490 45475
rect 7481 45373 7515 45407
rect 40141 45373 40175 45407
rect 28549 45305 28583 45339
rect 45569 45305 45603 45339
rect 6561 45237 6595 45271
rect 9321 45237 9355 45271
rect 37657 45237 37691 45271
rect 41521 45237 41555 45271
rect 7665 45033 7699 45067
rect 8309 45033 8343 45067
rect 9873 45033 9907 45067
rect 45845 45033 45879 45067
rect 10793 44965 10827 44999
rect 43821 44965 43855 44999
rect 6745 44897 6779 44931
rect 43637 44897 43671 44931
rect 6478 44829 6512 44863
rect 7297 44829 7331 44863
rect 8493 44829 8527 44863
rect 10517 44829 10551 44863
rect 10793 44829 10827 44863
rect 36921 44829 36955 44863
rect 40233 44829 40267 44863
rect 42073 44829 42107 44863
rect 42993 44829 43027 44863
rect 45385 44829 45419 44863
rect 46029 44829 46063 44863
rect 10057 44761 10091 44795
rect 10609 44761 10643 44795
rect 37166 44761 37200 44795
rect 40500 44761 40534 44795
rect 44097 44761 44131 44795
rect 5365 44693 5399 44727
rect 7665 44693 7699 44727
rect 7849 44693 7883 44727
rect 9689 44693 9723 44727
rect 9857 44693 9891 44727
rect 38301 44693 38335 44727
rect 41613 44693 41647 44727
rect 43177 44693 43211 44727
rect 45201 44693 45235 44727
rect 7113 44489 7147 44523
rect 9137 44489 9171 44523
rect 11161 44489 11195 44523
rect 45477 44489 45511 44523
rect 6929 44421 6963 44455
rect 7941 44421 7975 44455
rect 8769 44421 8803 44455
rect 9045 44421 9079 44455
rect 5825 44353 5859 44387
rect 5917 44353 5951 44387
rect 7757 44353 7791 44387
rect 8953 44353 8987 44387
rect 10037 44353 10071 44387
rect 36277 44353 36311 44387
rect 37740 44353 37774 44387
rect 40049 44353 40083 44387
rect 40316 44353 40350 44387
rect 41889 44353 41923 44387
rect 44557 44353 44591 44387
rect 9781 44285 9815 44319
rect 37473 44285 37507 44319
rect 45017 44285 45051 44319
rect 5641 44217 5675 44251
rect 6561 44217 6595 44251
rect 7573 44217 7607 44251
rect 9321 44217 9355 44251
rect 45293 44217 45327 44251
rect 6929 44149 6963 44183
rect 24593 44149 24627 44183
rect 36921 44149 36955 44183
rect 38853 44149 38887 44183
rect 39589 44149 39623 44183
rect 41429 44149 41463 44183
rect 43269 44149 43303 44183
rect 6469 43945 6503 43979
rect 9413 43945 9447 43979
rect 38485 43945 38519 43979
rect 41889 43945 41923 43979
rect 44649 43945 44683 43979
rect 45385 43945 45419 43979
rect 45569 43945 45603 43979
rect 9137 43809 9171 43843
rect 38669 43809 38703 43843
rect 41981 43809 42015 43843
rect 9321 43741 9355 43775
rect 9413 43741 9447 43775
rect 11253 43741 11287 43775
rect 12081 43741 12115 43775
rect 24593 43741 24627 43775
rect 24860 43741 24894 43775
rect 36185 43741 36219 43775
rect 36645 43741 36679 43775
rect 38761 43741 38795 43775
rect 40049 43741 40083 43775
rect 40316 43741 40350 43775
rect 42165 43741 42199 43775
rect 43269 43741 43303 43775
rect 6285 43673 6319 43707
rect 6501 43673 6535 43707
rect 10986 43673 11020 43707
rect 12348 43673 12382 43707
rect 36890 43673 36924 43707
rect 38485 43673 38519 43707
rect 41889 43673 41923 43707
rect 43514 43673 43548 43707
rect 45201 43673 45235 43707
rect 6653 43605 6687 43639
rect 9873 43605 9907 43639
rect 13461 43605 13495 43639
rect 25973 43605 26007 43639
rect 38025 43605 38059 43639
rect 38945 43605 38979 43639
rect 41429 43605 41463 43639
rect 42349 43605 42383 43639
rect 45401 43605 45435 43639
rect 11069 43401 11103 43435
rect 38853 43401 38887 43435
rect 43269 43401 43303 43435
rect 43729 43401 43763 43435
rect 5641 43333 5675 43367
rect 6745 43333 6779 43367
rect 37740 43333 37774 43367
rect 40969 43333 41003 43367
rect 44864 43333 44898 43367
rect 5825 43265 5859 43299
rect 7113 43265 7147 43299
rect 8769 43265 8803 43299
rect 10977 43265 11011 43299
rect 11161 43265 11195 43299
rect 12357 43265 12391 43299
rect 41061 43265 41095 43299
rect 41337 43265 41371 43299
rect 43085 43265 43119 43299
rect 43269 43265 43303 43299
rect 45109 43265 45143 43299
rect 37473 43197 37507 43231
rect 6009 43129 6043 43163
rect 41153 43129 41187 43163
rect 6561 43061 6595 43095
rect 6745 43061 6779 43095
rect 10057 43061 10091 43095
rect 41337 43061 41371 43095
rect 6377 42857 6411 42891
rect 6837 42857 6871 42891
rect 44465 42857 44499 42891
rect 7941 42789 7975 42823
rect 9137 42721 9171 42755
rect 4997 42653 5031 42687
rect 7024 42631 7058 42665
rect 7113 42653 7147 42687
rect 7297 42653 7331 42687
rect 7389 42653 7423 42687
rect 24593 42653 24627 42687
rect 33885 42653 33919 42687
rect 35081 42653 35115 42687
rect 37473 42653 37507 42687
rect 44097 42653 44131 42687
rect 44281 42653 44315 42687
rect 5264 42585 5298 42619
rect 8309 42585 8343 42619
rect 9382 42585 9416 42619
rect 7849 42517 7883 42551
rect 10517 42517 10551 42551
rect 38117 42517 38151 42551
rect 5733 42313 5767 42347
rect 9045 42313 9079 42347
rect 10149 42313 10183 42347
rect 24216 42245 24250 42279
rect 28825 42245 28859 42279
rect 31125 42245 31159 42279
rect 37473 42245 37507 42279
rect 5917 42177 5951 42211
rect 6745 42177 6779 42211
rect 7021 42177 7055 42211
rect 7205 42177 7239 42211
rect 8953 42177 8987 42211
rect 9137 42177 9171 42211
rect 9781 42177 9815 42211
rect 22017 42177 22051 42211
rect 22273 42177 22307 42211
rect 33876 42177 33910 42211
rect 36562 42177 36596 42211
rect 44281 42177 44315 42211
rect 44373 42177 44407 42211
rect 44557 42177 44591 42211
rect 44649 42177 44683 42211
rect 9873 42109 9907 42143
rect 21465 42109 21499 42143
rect 23949 42109 23983 42143
rect 33609 42109 33643 42143
rect 36829 42109 36863 42143
rect 30113 42041 30147 42075
rect 38761 42041 38795 42075
rect 44097 42041 44131 42075
rect 6561 41973 6595 42007
rect 12081 41973 12115 42007
rect 15301 41973 15335 42007
rect 23397 41973 23431 42007
rect 25329 41973 25363 42007
rect 34989 41973 35023 42007
rect 35449 41973 35483 42007
rect 40693 41973 40727 42007
rect 43453 41973 43487 42007
rect 45109 41973 45143 42007
rect 7021 41769 7055 41803
rect 7665 41769 7699 41803
rect 13277 41769 13311 41803
rect 27261 41769 27295 41803
rect 35357 41769 35391 41803
rect 35541 41769 35575 41803
rect 39037 41769 39071 41803
rect 39497 41769 39531 41803
rect 44649 41769 44683 41803
rect 34345 41701 34379 41735
rect 11161 41633 11195 41667
rect 24593 41633 24627 41667
rect 32965 41633 32999 41667
rect 35173 41633 35207 41667
rect 39129 41633 39163 41667
rect 40417 41633 40451 41667
rect 5641 41565 5675 41599
rect 5908 41565 5942 41599
rect 7481 41565 7515 41599
rect 7665 41565 7699 41599
rect 9321 41565 9355 41599
rect 13185 41565 13219 41599
rect 13277 41565 13311 41599
rect 14933 41565 14967 41599
rect 15200 41565 15234 41599
rect 16773 41565 16807 41599
rect 20729 41565 20763 41599
rect 24041 41565 24075 41599
rect 27077 41565 27111 41599
rect 27169 41565 27203 41599
rect 35357 41565 35391 41599
rect 37105 41565 37139 41599
rect 37372 41565 37406 41599
rect 39313 41565 39347 41599
rect 40684 41565 40718 41599
rect 43269 41565 43303 41599
rect 43536 41565 43570 41599
rect 11406 41497 11440 41531
rect 13001 41497 13035 41531
rect 20996 41497 21030 41531
rect 24838 41497 24872 41531
rect 27353 41497 27387 41531
rect 33232 41497 33266 41531
rect 35081 41497 35115 41531
rect 39037 41497 39071 41531
rect 12541 41429 12575 41463
rect 13461 41429 13495 41463
rect 16313 41429 16347 41463
rect 22109 41429 22143 41463
rect 25973 41429 26007 41463
rect 38485 41429 38519 41463
rect 41797 41429 41831 41463
rect 12173 41225 12207 41259
rect 25053 41225 25087 41259
rect 27537 41225 27571 41259
rect 34621 41225 34655 41259
rect 43637 41225 43671 41259
rect 22753 41157 22787 41191
rect 25513 41157 25547 41191
rect 44772 41157 44806 41191
rect 9137 41089 9171 41123
rect 9393 41089 9427 41123
rect 11161 41089 11195 41123
rect 13297 41089 13331 41123
rect 14013 41089 14047 41123
rect 15200 41089 15234 41123
rect 21097 41089 21131 41123
rect 23029 41089 23063 41123
rect 23673 41089 23707 41123
rect 23940 41089 23974 41123
rect 25789 41089 25823 41123
rect 28650 41089 28684 41123
rect 28917 41089 28951 41123
rect 30297 41089 30331 41123
rect 33241 41089 33275 41123
rect 33508 41089 33542 41123
rect 35081 41089 35115 41123
rect 37740 41089 37774 41123
rect 40868 41089 40902 41123
rect 45017 41089 45051 41123
rect 13553 41021 13587 41055
rect 14933 41021 14967 41055
rect 22937 41021 22971 41055
rect 25605 41021 25639 41055
rect 37473 41021 37507 41055
rect 40601 41021 40635 41055
rect 5549 40885 5583 40919
rect 10517 40885 10551 40919
rect 16313 40885 16347 40919
rect 22201 40885 22235 40919
rect 23029 40885 23063 40919
rect 23213 40885 23247 40919
rect 25513 40885 25547 40919
rect 25973 40885 26007 40919
rect 30113 40885 30147 40919
rect 38853 40885 38887 40919
rect 40141 40885 40175 40919
rect 41981 40885 42015 40919
rect 8585 40681 8619 40715
rect 13185 40681 13219 40715
rect 16773 40681 16807 40715
rect 24593 40681 24627 40715
rect 26341 40681 26375 40715
rect 33517 40681 33551 40715
rect 38761 40681 38795 40715
rect 39221 40681 39255 40715
rect 42165 40681 42199 40715
rect 42625 40681 42659 40715
rect 16313 40613 16347 40647
rect 38301 40613 38335 40647
rect 5273 40545 5307 40579
rect 9137 40545 9171 40579
rect 14933 40545 14967 40579
rect 16865 40545 16899 40579
rect 22293 40545 22327 40579
rect 25881 40545 25915 40579
rect 38853 40545 38887 40579
rect 5540 40477 5574 40511
rect 9404 40477 9438 40511
rect 11805 40477 11839 40511
rect 12072 40477 12106 40511
rect 14473 40477 14507 40511
rect 15189 40477 15223 40511
rect 17049 40477 17083 40511
rect 21741 40477 21775 40511
rect 25513 40477 25547 40511
rect 25697 40477 25731 40511
rect 26341 40477 26375 40511
rect 26525 40477 26559 40511
rect 27445 40477 27479 40511
rect 27905 40477 27939 40511
rect 27997 40477 28031 40511
rect 29837 40477 29871 40511
rect 30104 40477 30138 40511
rect 36461 40477 36495 40511
rect 36921 40477 36955 40511
rect 39037 40477 39071 40511
rect 40325 40477 40359 40511
rect 42349 40477 42383 40511
rect 42441 40477 42475 40511
rect 16773 40409 16807 40443
rect 24041 40409 24075 40443
rect 37166 40409 37200 40443
rect 38761 40409 38795 40443
rect 40592 40409 40626 40443
rect 42165 40409 42199 40443
rect 6653 40341 6687 40375
rect 10517 40341 10551 40375
rect 17233 40341 17267 40375
rect 26709 40341 26743 40375
rect 27788 40341 27822 40375
rect 31217 40341 31251 40375
rect 41705 40341 41739 40375
rect 7205 40137 7239 40171
rect 12725 40137 12759 40171
rect 23397 40137 23431 40171
rect 26617 40137 26651 40171
rect 28273 40137 28307 40171
rect 30389 40137 30423 40171
rect 38853 40137 38887 40171
rect 41797 40137 41831 40171
rect 10517 40069 10551 40103
rect 13829 40069 13863 40103
rect 40662 40069 40696 40103
rect 6837 40001 6871 40035
rect 8769 40001 8803 40035
rect 12909 40001 12943 40035
rect 13185 40001 13219 40035
rect 15393 40001 15427 40035
rect 15853 40001 15887 40035
rect 22017 40001 22051 40035
rect 22284 40001 22318 40035
rect 25237 40001 25271 40035
rect 25504 40001 25538 40035
rect 27169 40001 27203 40035
rect 27353 40001 27387 40035
rect 27629 40001 27663 40035
rect 27813 40001 27847 40035
rect 28457 40001 28491 40035
rect 29929 40001 29963 40035
rect 36921 40001 36955 40035
rect 37729 40001 37763 40035
rect 6929 39933 6963 39967
rect 13093 39933 13127 39967
rect 28733 39933 28767 39967
rect 37473 39933 37507 39967
rect 40417 39933 40451 39967
rect 11069 39865 11103 39899
rect 28641 39865 28675 39899
rect 30205 39865 30239 39899
rect 5641 39797 5675 39831
rect 6929 39797 6963 39831
rect 8309 39797 8343 39831
rect 13185 39797 13219 39831
rect 24225 39797 24259 39831
rect 6653 39593 6687 39627
rect 7297 39593 7331 39627
rect 7665 39593 7699 39627
rect 11161 39593 11195 39627
rect 11345 39593 11379 39627
rect 14473 39593 14507 39627
rect 16405 39593 16439 39627
rect 23581 39593 23615 39627
rect 37657 39593 37691 39627
rect 40693 39593 40727 39627
rect 41337 39593 41371 39627
rect 5273 39457 5307 39491
rect 7389 39457 7423 39491
rect 15025 39457 15059 39491
rect 22201 39457 22235 39491
rect 5540 39389 5574 39423
rect 7481 39389 7515 39423
rect 8309 39389 8343 39423
rect 9137 39389 9171 39423
rect 9393 39389 9427 39423
rect 10977 39389 11011 39423
rect 11161 39389 11195 39423
rect 15292 39389 15326 39423
rect 22468 39389 22502 39423
rect 7205 39321 7239 39355
rect 10517 39253 10551 39287
rect 9597 39049 9631 39083
rect 27169 39049 27203 39083
rect 7297 38981 7331 39015
rect 27353 38981 27387 39015
rect 27721 38981 27755 39015
rect 23213 38913 23247 38947
rect 23480 38913 23514 38947
rect 27445 38913 27479 38947
rect 27537 38913 27571 38947
rect 30573 38913 30607 38947
rect 30757 38913 30791 38947
rect 40785 38913 40819 38947
rect 40969 38913 41003 38947
rect 5733 38709 5767 38743
rect 6745 38709 6779 38743
rect 8769 38709 8803 38743
rect 11713 38709 11747 38743
rect 24593 38709 24627 38743
rect 30665 38709 30699 38743
rect 36737 38709 36771 38743
rect 41153 38709 41187 38743
rect 7113 38505 7147 38539
rect 12633 38505 12667 38539
rect 13093 38505 13127 38539
rect 13553 38505 13587 38539
rect 23121 38505 23155 38539
rect 26893 38505 26927 38539
rect 28825 38505 28859 38539
rect 30021 38505 30055 38539
rect 30941 38505 30975 38539
rect 39221 38505 39255 38539
rect 42625 38505 42659 38539
rect 43453 38505 43487 38539
rect 6653 38437 6687 38471
rect 26709 38437 26743 38471
rect 27261 38437 27295 38471
rect 28641 38437 28675 38471
rect 30205 38437 30239 38471
rect 5273 38369 5307 38403
rect 13185 38369 13219 38403
rect 5540 38301 5574 38335
rect 8237 38301 8271 38335
rect 8493 38301 8527 38335
rect 10609 38301 10643 38335
rect 11253 38301 11287 38335
rect 13369 38301 13403 38335
rect 23581 38301 23615 38335
rect 26065 38301 26099 38335
rect 27905 38301 27939 38335
rect 28181 38301 28215 38335
rect 31677 38301 31711 38335
rect 36093 38301 36127 38335
rect 36553 38301 36587 38335
rect 40049 38301 40083 38335
rect 40693 38301 40727 38335
rect 43269 38301 43303 38335
rect 11520 38233 11554 38267
rect 13093 38233 13127 38267
rect 29009 38233 29043 38267
rect 29837 38233 29871 38267
rect 30757 38233 30791 38267
rect 36798 38233 36832 38267
rect 40960 38233 40994 38267
rect 26249 38165 26283 38199
rect 26893 38165 26927 38199
rect 27721 38165 27755 38199
rect 28089 38165 28123 38199
rect 28799 38165 28833 38199
rect 30037 38165 30071 38199
rect 30957 38165 30991 38199
rect 31125 38165 31159 38199
rect 31861 38165 31895 38199
rect 37933 38165 37967 38199
rect 40233 38165 40267 38199
rect 42073 38165 42107 38199
rect 8125 37961 8159 37995
rect 11161 37961 11195 37995
rect 13921 37961 13955 37995
rect 27337 37961 27371 37995
rect 27997 37961 28031 37995
rect 30297 37961 30331 37995
rect 31125 37961 31159 37995
rect 42073 37961 42107 37995
rect 10048 37893 10082 37927
rect 12786 37893 12820 37927
rect 23572 37893 23606 37927
rect 27537 37893 27571 37927
rect 29377 37893 29411 37927
rect 29561 37893 29595 37927
rect 31309 37893 31343 37927
rect 32566 37893 32600 37927
rect 39405 37893 39439 37927
rect 42809 37893 42843 37927
rect 44557 37893 44591 37927
rect 6745 37825 6779 37859
rect 7012 37825 7046 37859
rect 12081 37825 12115 37859
rect 12541 37825 12575 37859
rect 23305 37825 23339 37859
rect 28181 37825 28215 37859
rect 28365 37825 28399 37859
rect 29653 37825 29687 37859
rect 30389 37825 30423 37859
rect 30481 37825 30515 37859
rect 31493 37825 31527 37859
rect 36654 37825 36688 37859
rect 36921 37825 36955 37859
rect 37740 37825 37774 37859
rect 9781 37757 9815 37791
rect 32321 37757 32355 37791
rect 37473 37757 37507 37791
rect 41613 37757 41647 37791
rect 30113 37689 30147 37723
rect 30665 37689 30699 37723
rect 41889 37689 41923 37723
rect 5825 37621 5859 37655
rect 24685 37621 24719 37655
rect 27169 37621 27203 37655
rect 27353 37621 27387 37655
rect 29653 37621 29687 37655
rect 33701 37621 33735 37655
rect 35541 37621 35575 37655
rect 38853 37621 38887 37655
rect 40693 37621 40727 37655
rect 13001 37417 13035 37451
rect 24593 37417 24627 37451
rect 27445 37417 27479 37451
rect 28825 37417 28859 37451
rect 31125 37417 31159 37451
rect 38209 37417 38243 37451
rect 39405 37417 39439 37451
rect 42073 37417 42107 37451
rect 42717 37417 42751 37451
rect 28641 37349 28675 37383
rect 29193 37349 29227 37383
rect 5549 37281 5583 37315
rect 24685 37281 24719 37315
rect 31861 37281 31895 37315
rect 38301 37281 38335 37315
rect 40049 37281 40083 37315
rect 5816 37213 5850 37247
rect 11621 37213 11655 37247
rect 22661 37213 22695 37247
rect 24869 37213 24903 37247
rect 26065 37213 26099 37247
rect 26332 37213 26366 37247
rect 27997 37213 28031 37247
rect 29745 37213 29779 37247
rect 30001 37213 30035 37247
rect 31769 37213 31803 37247
rect 31953 37213 31987 37247
rect 32045 37213 32079 37247
rect 36369 37213 36403 37247
rect 38485 37213 38519 37247
rect 39313 37213 39347 37247
rect 39497 37213 39531 37247
rect 40316 37213 40350 37247
rect 42901 37213 42935 37247
rect 11888 37145 11922 37179
rect 22928 37145 22962 37179
rect 24593 37145 24627 37179
rect 36636 37145 36670 37179
rect 38209 37145 38243 37179
rect 41889 37145 41923 37179
rect 42089 37145 42123 37179
rect 6929 37077 6963 37111
rect 24041 37077 24075 37111
rect 25053 37077 25087 37111
rect 28181 37077 28215 37111
rect 28825 37077 28859 37111
rect 31585 37077 31619 37111
rect 37749 37077 37783 37111
rect 38669 37077 38703 37111
rect 41429 37077 41463 37111
rect 42257 37077 42291 37111
rect 24869 36873 24903 36907
rect 26617 36873 26651 36907
rect 28549 36873 28583 36907
rect 31309 36873 31343 36907
rect 32413 36873 32447 36907
rect 40141 36873 40175 36907
rect 40325 36873 40359 36907
rect 30021 36805 30055 36839
rect 11897 36737 11931 36771
rect 22845 36737 22879 36771
rect 23756 36737 23790 36771
rect 26433 36737 26467 36771
rect 26617 36737 26651 36771
rect 27169 36737 27203 36771
rect 27425 36737 27459 36771
rect 36645 36737 36679 36771
rect 37657 36737 37691 36771
rect 39497 36737 39531 36771
rect 41153 36737 41187 36771
rect 41337 36737 41371 36771
rect 23489 36669 23523 36703
rect 39681 36669 39715 36703
rect 39313 36601 39347 36635
rect 40693 36601 40727 36635
rect 33333 36533 33367 36567
rect 40325 36533 40359 36567
rect 41521 36533 41555 36567
rect 23765 36329 23799 36363
rect 27261 36329 27295 36363
rect 29745 36329 29779 36363
rect 40325 36329 40359 36363
rect 31125 36193 31159 36227
rect 32965 36193 32999 36227
rect 36185 36193 36219 36227
rect 27077 36125 27111 36159
rect 31769 36125 31803 36159
rect 33232 36125 33266 36159
rect 40693 36125 40727 36159
rect 30880 36057 30914 36091
rect 36452 36057 36486 36091
rect 40325 36057 40359 36091
rect 31585 35989 31619 36023
rect 34345 35989 34379 36023
rect 37565 35989 37599 36023
rect 40141 35989 40175 36023
rect 25973 35785 26007 35819
rect 30021 35785 30055 35819
rect 30389 35785 30423 35819
rect 41153 35785 41187 35819
rect 33302 35717 33336 35751
rect 40040 35717 40074 35751
rect 25605 35649 25639 35683
rect 25789 35649 25823 35683
rect 30205 35649 30239 35683
rect 30481 35649 30515 35683
rect 32597 35649 32631 35683
rect 33057 35649 33091 35683
rect 39773 35581 39807 35615
rect 22017 35445 22051 35479
rect 25605 35445 25639 35479
rect 34437 35445 34471 35479
rect 34897 35445 34931 35479
rect 36553 35445 36587 35479
rect 23121 35241 23155 35275
rect 23581 35241 23615 35275
rect 34897 35241 34931 35275
rect 38117 35241 38151 35275
rect 40233 35241 40267 35275
rect 34345 35173 34379 35207
rect 25053 35105 25087 35139
rect 32965 35105 32999 35139
rect 34989 35105 35023 35139
rect 20821 35037 20855 35071
rect 21281 35037 21315 35071
rect 23305 35037 23339 35071
rect 23397 35037 23431 35071
rect 25320 35037 25354 35071
rect 26893 35037 26927 35071
rect 33232 35037 33266 35071
rect 34897 35037 34931 35071
rect 35173 35037 35207 35071
rect 36277 35037 36311 35071
rect 36544 35037 36578 35071
rect 40417 35037 40451 35071
rect 21526 34969 21560 35003
rect 23121 34969 23155 35003
rect 22661 34901 22695 34935
rect 26433 34901 26467 34935
rect 35357 34901 35391 34935
rect 37657 34901 37691 34935
rect 20085 34697 20119 34731
rect 23397 34697 23431 34731
rect 25973 34697 26007 34731
rect 34989 34697 35023 34731
rect 21220 34629 21254 34663
rect 37473 34629 37507 34663
rect 22284 34561 22318 34595
rect 24593 34561 24627 34595
rect 24860 34561 24894 34595
rect 33876 34561 33910 34595
rect 37749 34561 37783 34595
rect 39681 34561 39715 34595
rect 39773 34561 39807 34595
rect 39957 34561 39991 34595
rect 21465 34493 21499 34527
rect 22017 34493 22051 34527
rect 33609 34493 33643 34527
rect 37565 34493 37599 34527
rect 28181 34357 28215 34391
rect 28825 34357 28859 34391
rect 31309 34357 31343 34391
rect 36461 34357 36495 34391
rect 37657 34357 37691 34391
rect 37933 34357 37967 34391
rect 40141 34357 40175 34391
rect 21097 34153 21131 34187
rect 22937 34153 22971 34187
rect 26617 34153 26651 34187
rect 27077 34153 27111 34187
rect 33057 34153 33091 34187
rect 33977 34153 34011 34187
rect 37565 34153 37599 34187
rect 39313 34153 39347 34187
rect 39497 34153 39531 34187
rect 40233 34153 40267 34187
rect 26157 34085 26191 34119
rect 32321 34085 32355 34119
rect 40601 34085 40635 34119
rect 21557 34017 21591 34051
rect 24777 34017 24811 34051
rect 26709 34017 26743 34051
rect 27813 34017 27847 34051
rect 32873 34017 32907 34051
rect 24041 33949 24075 33983
rect 26893 33949 26927 33983
rect 28080 33949 28114 33983
rect 30481 33949 30515 33983
rect 30941 33949 30975 33983
rect 31208 33949 31242 33983
rect 33057 33949 33091 33983
rect 36185 33949 36219 33983
rect 38025 33949 38059 33983
rect 38209 33949 38243 33983
rect 41061 33949 41095 33983
rect 41245 33949 41279 33983
rect 43453 33949 43487 33983
rect 21824 33881 21858 33915
rect 25044 33881 25078 33915
rect 26617 33881 26651 33915
rect 32781 33881 32815 33915
rect 36452 33881 36486 33915
rect 39129 33881 39163 33915
rect 40233 33881 40267 33915
rect 29193 33813 29227 33847
rect 33241 33813 33275 33847
rect 38117 33813 38151 33847
rect 39329 33813 39363 33847
rect 40049 33813 40083 33847
rect 41153 33813 41187 33847
rect 43269 33813 43303 33847
rect 25237 33609 25271 33643
rect 31769 33609 31803 33643
rect 33701 33609 33735 33643
rect 40049 33609 40083 33643
rect 41889 33609 41923 33643
rect 28172 33541 28206 33575
rect 32566 33541 32600 33575
rect 43260 33541 43294 33575
rect 22017 33473 22051 33507
rect 23949 33473 23983 33507
rect 30389 33473 30423 33507
rect 30656 33473 30690 33507
rect 38936 33473 38970 33507
rect 40509 33473 40543 33507
rect 40776 33473 40810 33507
rect 26157 33405 26191 33439
rect 27905 33405 27939 33439
rect 32321 33405 32355 33439
rect 38669 33405 38703 33439
rect 42993 33405 43027 33439
rect 27445 33269 27479 33303
rect 29285 33269 29319 33303
rect 29929 33269 29963 33303
rect 44373 33269 44407 33303
rect 25973 33065 26007 33099
rect 26433 33065 26467 33099
rect 29745 33065 29779 33099
rect 32505 33065 32539 33099
rect 33057 33065 33091 33099
rect 33425 33065 33459 33099
rect 39221 33065 39255 33099
rect 40233 33065 40267 33099
rect 40877 33065 40911 33099
rect 42441 33065 42475 33099
rect 43545 33065 43579 33099
rect 45385 33065 45419 33099
rect 29193 32997 29227 33031
rect 40417 32997 40451 33031
rect 43361 32997 43395 33031
rect 24593 32929 24627 32963
rect 29837 32929 29871 32963
rect 27813 32861 27847 32895
rect 28069 32861 28103 32895
rect 30021 32861 30055 32895
rect 31125 32861 31159 32895
rect 33149 32861 33183 32895
rect 33241 32861 33275 32895
rect 35081 32861 35115 32895
rect 39405 32861 39439 32895
rect 41061 32861 41095 32895
rect 24860 32793 24894 32827
rect 29745 32793 29779 32827
rect 31392 32793 31426 32827
rect 32965 32793 32999 32827
rect 40049 32793 40083 32827
rect 42625 32793 42659 32827
rect 43085 32793 43119 32827
rect 45201 32793 45235 32827
rect 30205 32725 30239 32759
rect 40249 32725 40283 32759
rect 42257 32725 42291 32759
rect 42425 32725 42459 32759
rect 45401 32725 45435 32759
rect 45569 32725 45603 32759
rect 35633 32521 35667 32555
rect 40325 32521 40359 32555
rect 42073 32521 42107 32555
rect 42625 32521 42659 32555
rect 42993 32521 43027 32555
rect 43821 32521 43855 32555
rect 45109 32521 45143 32555
rect 36921 32453 36955 32487
rect 37473 32453 37507 32487
rect 24777 32385 24811 32419
rect 31125 32385 31159 32419
rect 35817 32385 35851 32419
rect 36093 32385 36127 32419
rect 39957 32385 39991 32419
rect 40141 32385 40175 32419
rect 41153 32385 41187 32419
rect 41797 32385 41831 32419
rect 41981 32385 42015 32419
rect 42073 32385 42107 32419
rect 42809 32385 42843 32419
rect 43085 32385 43119 32419
rect 43729 32385 43763 32419
rect 43913 32385 43947 32419
rect 46222 32385 46256 32419
rect 36001 32317 36035 32351
rect 46489 32317 46523 32351
rect 44097 32249 44131 32283
rect 27813 32181 27847 32215
rect 34989 32181 35023 32215
rect 36093 32181 36127 32215
rect 38761 32181 38795 32215
rect 41337 32181 41371 32215
rect 43545 32181 43579 32215
rect 28917 31977 28951 32011
rect 36277 31977 36311 32011
rect 42993 31977 43027 32011
rect 44557 31977 44591 32011
rect 45569 31977 45603 32011
rect 46213 31977 46247 32011
rect 27537 31841 27571 31875
rect 43453 31841 43487 31875
rect 43729 31841 43763 31875
rect 43821 31841 43855 31875
rect 43913 31841 43947 31875
rect 27793 31773 27827 31807
rect 34345 31773 34379 31807
rect 34897 31773 34931 31807
rect 35164 31773 35198 31807
rect 36737 31773 36771 31807
rect 41613 31773 41647 31807
rect 41880 31773 41914 31807
rect 43637 31773 43671 31807
rect 44465 31773 44499 31807
rect 44649 31773 44683 31807
rect 45385 31773 45419 31807
rect 46029 31773 46063 31807
rect 45201 31705 45235 31739
rect 36461 31433 36495 31467
rect 32413 31365 32447 31399
rect 32873 31365 32907 31399
rect 43729 31365 43763 31399
rect 44281 31365 44315 31399
rect 23213 31297 23247 31331
rect 23480 31297 23514 31331
rect 35337 31297 35371 31331
rect 41889 31297 41923 31331
rect 34621 31229 34655 31263
rect 35081 31229 35115 31263
rect 45569 31161 45603 31195
rect 24593 31093 24627 31127
rect 30849 31093 30883 31127
rect 31493 31093 31527 31127
rect 42073 31093 42107 31127
rect 43637 31093 43671 31127
rect 31953 30889 31987 30923
rect 32413 30889 32447 30923
rect 32873 30889 32907 30923
rect 36277 30889 36311 30923
rect 44005 30889 44039 30923
rect 44465 30889 44499 30923
rect 32505 30753 32539 30787
rect 23581 30685 23615 30719
rect 30573 30685 30607 30719
rect 32689 30685 32723 30719
rect 34897 30685 34931 30719
rect 42625 30685 42659 30719
rect 42881 30685 42915 30719
rect 30840 30617 30874 30651
rect 32413 30617 32447 30651
rect 35164 30617 35198 30651
rect 42717 30345 42751 30379
rect 23572 30277 23606 30311
rect 30656 30277 30690 30311
rect 35940 30277 35974 30311
rect 42901 30277 42935 30311
rect 25145 30209 25179 30243
rect 30389 30209 30423 30243
rect 43269 30209 43303 30243
rect 23305 30141 23339 30175
rect 36185 30141 36219 30175
rect 31769 30073 31803 30107
rect 22845 30005 22879 30039
rect 24685 30005 24719 30039
rect 32321 30005 32355 30039
rect 34805 30005 34839 30039
rect 42901 30005 42935 30039
rect 24685 29801 24719 29835
rect 32781 29801 32815 29835
rect 24685 29665 24719 29699
rect 31401 29665 31435 29699
rect 22109 29597 22143 29631
rect 22569 29597 22603 29631
rect 24869 29597 24903 29631
rect 30389 29597 30423 29631
rect 31668 29597 31702 29631
rect 44373 29597 44407 29631
rect 46581 29597 46615 29631
rect 22814 29529 22848 29563
rect 24593 29529 24627 29563
rect 46314 29529 46348 29563
rect 23949 29461 23983 29495
rect 25053 29461 25087 29495
rect 44557 29461 44591 29495
rect 45201 29461 45235 29495
rect 24685 29257 24719 29291
rect 31401 29257 31435 29291
rect 43913 29257 43947 29291
rect 23550 29189 23584 29223
rect 42993 29189 43027 29223
rect 43545 29189 43579 29223
rect 43761 29189 43795 29223
rect 44373 29189 44407 29223
rect 45293 29189 45327 29223
rect 45493 29189 45527 29223
rect 23305 29121 23339 29155
rect 30021 29121 30055 29155
rect 30288 29121 30322 29155
rect 42901 29121 42935 29155
rect 43085 29121 43119 29155
rect 44557 29121 44591 29155
rect 44741 29121 44775 29155
rect 44833 29121 44867 29155
rect 46121 29121 46155 29155
rect 35541 28985 35575 29019
rect 38669 28985 38703 29019
rect 45661 28985 45695 29019
rect 17325 28917 17359 28951
rect 18337 28917 18371 28951
rect 36185 28917 36219 28951
rect 43729 28917 43763 28951
rect 45477 28917 45511 28951
rect 46305 28917 46339 28951
rect 32505 28713 32539 28747
rect 44649 28577 44683 28611
rect 17049 28509 17083 28543
rect 17316 28509 17350 28543
rect 24777 28509 24811 28543
rect 35265 28509 35299 28543
rect 38761 28509 38795 28543
rect 42993 28509 43027 28543
rect 43269 28509 43303 28543
rect 44281 28509 44315 28543
rect 44465 28509 44499 28543
rect 46314 28509 46348 28543
rect 46581 28509 46615 28543
rect 31217 28441 31251 28475
rect 35532 28441 35566 28475
rect 43177 28441 43211 28475
rect 18429 28373 18463 28407
rect 30665 28373 30699 28407
rect 36645 28373 36679 28407
rect 42809 28373 42843 28407
rect 45201 28373 45235 28407
rect 19441 28169 19475 28203
rect 36461 28169 36495 28203
rect 42073 28169 42107 28203
rect 44005 28169 44039 28203
rect 45293 28169 45327 28203
rect 18328 28101 18362 28135
rect 35326 28101 35360 28135
rect 37473 28101 37507 28135
rect 38660 28101 38694 28135
rect 42870 28101 42904 28135
rect 44925 28101 44959 28135
rect 19901 28033 19935 28067
rect 20085 28033 20119 28067
rect 20177 28033 20211 28067
rect 23397 28033 23431 28067
rect 34621 28033 34655 28067
rect 35081 28033 35115 28067
rect 37657 28033 37691 28067
rect 37749 28033 37783 28067
rect 38393 28033 38427 28067
rect 41889 28033 41923 28067
rect 42625 28033 42659 28067
rect 45109 28033 45143 28067
rect 18061 27965 18095 27999
rect 22845 27897 22879 27931
rect 16313 27829 16347 27863
rect 17325 27829 17359 27863
rect 19901 27829 19935 27863
rect 20361 27829 20395 27863
rect 21097 27829 21131 27863
rect 24685 27829 24719 27863
rect 25605 27829 25639 27863
rect 28641 27829 28675 27863
rect 32321 27829 32355 27863
rect 32965 27829 32999 27863
rect 37473 27829 37507 27863
rect 37933 27829 37967 27863
rect 39773 27829 39807 27863
rect 40233 27829 40267 27863
rect 42533 27625 42567 27659
rect 42717 27625 42751 27659
rect 43729 27625 43763 27659
rect 18429 27557 18463 27591
rect 36553 27557 36587 27591
rect 43085 27557 43119 27591
rect 43545 27557 43579 27591
rect 45293 27557 45327 27591
rect 17049 27421 17083 27455
rect 17316 27421 17350 27455
rect 20729 27421 20763 27455
rect 20996 27421 21030 27455
rect 23213 27421 23247 27455
rect 24041 27421 24075 27455
rect 25706 27421 25740 27455
rect 25973 27421 26007 27455
rect 27721 27421 27755 27455
rect 31217 27421 31251 27455
rect 31677 27421 31711 27455
rect 35173 27421 35207 27455
rect 35440 27421 35474 27455
rect 37013 27421 37047 27455
rect 38117 27421 38151 27455
rect 40049 27421 40083 27455
rect 45201 27421 45235 27455
rect 45385 27421 45419 27455
rect 27966 27353 28000 27387
rect 31944 27353 31978 27387
rect 38384 27353 38418 27387
rect 40316 27353 40350 27387
rect 42717 27353 42751 27387
rect 43713 27353 43747 27387
rect 43913 27353 43947 27387
rect 22109 27285 22143 27319
rect 24593 27285 24627 27319
rect 29101 27285 29135 27319
rect 33057 27285 33091 27319
rect 39497 27285 39531 27319
rect 41429 27285 41463 27319
rect 18245 27081 18279 27115
rect 36737 27081 36771 27115
rect 44005 27081 44039 27115
rect 17110 27013 17144 27047
rect 23020 27013 23054 27047
rect 24860 27013 24894 27047
rect 28242 27013 28276 27047
rect 32566 27013 32600 27047
rect 38660 27013 38694 27047
rect 40233 27013 40267 27047
rect 44189 27013 44223 27047
rect 16865 26945 16899 26979
rect 27537 26945 27571 26979
rect 27997 26945 28031 26979
rect 30389 26945 30423 26979
rect 30656 26945 30690 26979
rect 35357 26945 35391 26979
rect 35624 26945 35658 26979
rect 38393 26945 38427 26979
rect 40509 26945 40543 26979
rect 42901 26945 42935 26979
rect 43085 26945 43119 26979
rect 44097 26945 44131 26979
rect 58081 26945 58115 26979
rect 22753 26877 22787 26911
rect 24593 26877 24627 26911
rect 32321 26877 32355 26911
rect 37933 26877 37967 26911
rect 40325 26877 40359 26911
rect 42993 26877 43027 26911
rect 43177 26877 43211 26911
rect 39773 26809 39807 26843
rect 43821 26809 43855 26843
rect 24133 26741 24167 26775
rect 25973 26741 26007 26775
rect 26617 26741 26651 26775
rect 29377 26741 29411 26775
rect 31769 26741 31803 26775
rect 33701 26741 33735 26775
rect 40233 26741 40267 26775
rect 40693 26741 40727 26775
rect 43361 26741 43395 26775
rect 44373 26741 44407 26775
rect 58265 26741 58299 26775
rect 20729 26537 20763 26571
rect 27353 26537 27387 26571
rect 38577 26537 38611 26571
rect 43453 26537 43487 26571
rect 44097 26537 44131 26571
rect 24593 26401 24627 26435
rect 27813 26401 27847 26435
rect 38577 26401 38611 26435
rect 13553 26333 13587 26367
rect 24860 26333 24894 26367
rect 28080 26333 28114 26367
rect 30113 26333 30147 26367
rect 31861 26333 31895 26367
rect 32321 26333 32355 26367
rect 38485 26333 38519 26367
rect 42073 26333 42107 26367
rect 43913 26333 43947 26367
rect 44005 26333 44039 26367
rect 18889 26265 18923 26299
rect 19441 26265 19475 26299
rect 32588 26265 32622 26299
rect 42318 26265 42352 26299
rect 44189 26265 44223 26299
rect 13369 26197 13403 26231
rect 25973 26197 26007 26231
rect 29193 26197 29227 26231
rect 33701 26197 33735 26231
rect 38853 26197 38887 26231
rect 24133 25993 24167 26027
rect 41889 25993 41923 26027
rect 13176 25925 13210 25959
rect 25053 25925 25087 25959
rect 33701 25925 33735 25959
rect 45560 25925 45594 25959
rect 18889 25857 18923 25891
rect 19073 25857 19107 25891
rect 19257 25857 19291 25891
rect 22017 25857 22051 25891
rect 22293 25857 22327 25891
rect 24317 25857 24351 25891
rect 24593 25857 24627 25891
rect 25329 25857 25363 25891
rect 27813 25857 27847 25891
rect 28069 25857 28103 25891
rect 29745 25857 29779 25891
rect 30021 25857 30055 25891
rect 32505 25857 32539 25891
rect 33425 25857 33459 25891
rect 42073 25857 42107 25891
rect 43453 25857 43487 25891
rect 44097 25857 44131 25891
rect 44373 25857 44407 25891
rect 45293 25857 45327 25891
rect 12909 25789 12943 25823
rect 18705 25789 18739 25823
rect 22109 25789 22143 25823
rect 24409 25789 24443 25823
rect 25237 25789 25271 25823
rect 29837 25789 29871 25823
rect 33609 25789 33643 25823
rect 22477 25721 22511 25755
rect 25513 25721 25547 25755
rect 43085 25721 43119 25755
rect 14289 25653 14323 25687
rect 17325 25653 17359 25687
rect 20729 25653 20763 25687
rect 21189 25653 21223 25687
rect 22293 25653 22327 25687
rect 24593 25653 24627 25687
rect 25053 25653 25087 25687
rect 29193 25653 29227 25687
rect 29745 25653 29779 25687
rect 30205 25653 30239 25687
rect 31769 25653 31803 25687
rect 33241 25653 33275 25687
rect 33425 25653 33459 25687
rect 40325 25653 40359 25687
rect 46673 25653 46707 25687
rect 13277 25449 13311 25483
rect 22201 25449 22235 25483
rect 33241 25449 33275 25483
rect 44097 25449 44131 25483
rect 13461 25381 13495 25415
rect 20821 25313 20855 25347
rect 33149 25313 33183 25347
rect 13737 25245 13771 25279
rect 14473 25245 14507 25279
rect 17049 25245 17083 25279
rect 17316 25245 17350 25279
rect 20361 25245 20395 25279
rect 21088 25245 21122 25279
rect 24777 25245 24811 25279
rect 30665 25245 30699 25279
rect 33057 25245 33091 25279
rect 33333 25245 33367 25279
rect 33977 25245 34011 25279
rect 36277 25245 36311 25279
rect 36921 25245 36955 25279
rect 38577 25245 38611 25279
rect 39497 25245 39531 25279
rect 40049 25245 40083 25279
rect 40316 25245 40350 25279
rect 42717 25245 42751 25279
rect 14289 25177 14323 25211
rect 42984 25177 43018 25211
rect 14657 25109 14691 25143
rect 18429 25109 18463 25143
rect 33517 25109 33551 25143
rect 41429 25109 41463 25143
rect 14581 24905 14615 24939
rect 21465 24905 21499 24939
rect 42717 24905 42751 24939
rect 43821 24905 43855 24939
rect 13645 24837 13679 24871
rect 14381 24837 14415 24871
rect 38568 24837 38602 24871
rect 12817 24769 12851 24803
rect 13553 24769 13587 24803
rect 13829 24769 13863 24803
rect 15209 24769 15243 24803
rect 17601 24769 17635 24803
rect 17868 24769 17902 24803
rect 19441 24769 19475 24803
rect 20085 24769 20119 24803
rect 20352 24769 20386 24803
rect 23121 24769 23155 24803
rect 23673 24769 23707 24803
rect 30369 24769 30403 24803
rect 32965 24769 32999 24803
rect 33681 24769 33715 24803
rect 35808 24769 35842 24803
rect 37473 24769 37507 24803
rect 38301 24769 38335 24803
rect 40141 24769 40175 24803
rect 40397 24769 40431 24803
rect 42901 24769 42935 24803
rect 43361 24769 43395 24803
rect 44005 24769 44039 24803
rect 44281 24769 44315 24803
rect 30113 24701 30147 24735
rect 33425 24701 33459 24735
rect 35541 24701 35575 24735
rect 37565 24701 37599 24735
rect 43085 24701 43119 24735
rect 14749 24633 14783 24667
rect 24961 24633 24995 24667
rect 37841 24633 37875 24667
rect 44189 24633 44223 24667
rect 13001 24565 13035 24599
rect 13553 24565 13587 24599
rect 14565 24565 14599 24599
rect 15393 24565 15427 24599
rect 17141 24565 17175 24599
rect 18981 24565 19015 24599
rect 29653 24565 29687 24599
rect 31493 24565 31527 24599
rect 34805 24565 34839 24599
rect 36921 24565 36955 24599
rect 37473 24565 37507 24599
rect 39681 24565 39715 24599
rect 41521 24565 41555 24599
rect 43177 24565 43211 24599
rect 22109 24361 22143 24395
rect 31309 24361 31343 24395
rect 31769 24361 31803 24395
rect 32229 24361 32263 24395
rect 34345 24361 34379 24395
rect 34897 24361 34931 24395
rect 42809 24361 42843 24395
rect 12541 24293 12575 24327
rect 35265 24293 35299 24327
rect 17325 24225 17359 24259
rect 24593 24225 24627 24259
rect 29929 24225 29963 24259
rect 31861 24225 31895 24259
rect 34989 24225 35023 24259
rect 37841 24225 37875 24259
rect 13461 24157 13495 24191
rect 13737 24157 13771 24191
rect 16037 24157 16071 24191
rect 16865 24157 16899 24191
rect 17581 24157 17615 24191
rect 20729 24157 20763 24191
rect 23029 24157 23063 24191
rect 24041 24157 24075 24191
rect 29193 24157 29227 24191
rect 30185 24157 30219 24191
rect 32045 24157 32079 24191
rect 32965 24157 32999 24191
rect 33232 24157 33266 24191
rect 34897 24157 34931 24191
rect 12817 24089 12851 24123
rect 15770 24089 15804 24123
rect 20996 24089 21030 24123
rect 24860 24089 24894 24123
rect 31769 24089 31803 24123
rect 36093 24089 36127 24123
rect 41521 24089 41555 24123
rect 12357 24021 12391 24055
rect 13277 24021 13311 24055
rect 13645 24021 13679 24055
rect 14657 24021 14691 24055
rect 18705 24021 18739 24055
rect 25973 24021 26007 24055
rect 38393 24021 38427 24055
rect 41061 24021 41095 24055
rect 18429 23817 18463 23851
rect 19349 23817 19383 23851
rect 26065 23817 26099 23851
rect 31677 23817 31711 23851
rect 34621 23817 34655 23851
rect 36921 23817 36955 23851
rect 39221 23817 39255 23851
rect 42993 23817 43027 23851
rect 14749 23749 14783 23783
rect 17294 23749 17328 23783
rect 18889 23749 18923 23783
rect 30564 23749 30598 23783
rect 11897 23681 11931 23715
rect 12081 23681 12115 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 15669 23681 15703 23715
rect 15853 23681 15887 23715
rect 17049 23681 17083 23715
rect 19165 23681 19199 23715
rect 23305 23681 23339 23715
rect 23765 23681 23799 23715
rect 24032 23681 24066 23715
rect 25605 23681 25639 23715
rect 25881 23681 25915 23715
rect 29837 23681 29871 23715
rect 30297 23681 30331 23715
rect 33241 23681 33275 23715
rect 33508 23681 33542 23715
rect 35541 23681 35575 23715
rect 35808 23681 35842 23715
rect 37841 23681 37875 23715
rect 38097 23681 38131 23715
rect 40049 23681 40083 23715
rect 40316 23681 40350 23715
rect 42625 23681 42659 23715
rect 42809 23681 42843 23715
rect 11989 23613 12023 23647
rect 18981 23613 19015 23647
rect 25789 23613 25823 23647
rect 13461 23477 13495 23511
rect 15209 23477 15243 23511
rect 18889 23477 18923 23511
rect 25145 23477 25179 23511
rect 25605 23477 25639 23511
rect 41429 23477 41463 23511
rect 12357 23273 12391 23307
rect 14841 23273 14875 23307
rect 16221 23273 16255 23307
rect 24041 23273 24075 23307
rect 25973 23273 26007 23307
rect 31125 23273 31159 23307
rect 33609 23273 33643 23307
rect 36553 23273 36587 23307
rect 40233 23273 40267 23307
rect 41153 23273 41187 23307
rect 15577 23205 15611 23239
rect 41337 23205 41371 23239
rect 13737 23137 13771 23171
rect 14381 23137 14415 23171
rect 14657 23137 14691 23171
rect 24593 23137 24627 23171
rect 41061 23137 41095 23171
rect 3065 23069 3099 23103
rect 14473 23069 14507 23103
rect 14565 23069 14599 23103
rect 15485 23069 15519 23103
rect 15669 23069 15703 23103
rect 22661 23069 22695 23103
rect 24860 23069 24894 23103
rect 29745 23069 29779 23103
rect 40877 23069 40911 23103
rect 41153 23069 41187 23103
rect 13492 23001 13526 23035
rect 22928 23001 22962 23035
rect 29990 23001 30024 23035
rect 2881 22933 2915 22967
rect 12173 22729 12207 22763
rect 15301 22729 15335 22763
rect 2728 22661 2762 22695
rect 13286 22661 13320 22695
rect 13553 22593 13587 22627
rect 14013 22593 14047 22627
rect 37841 22593 37875 22627
rect 38025 22593 38059 22627
rect 2973 22525 3007 22559
rect 1593 22389 1627 22423
rect 16865 22389 16899 22423
rect 37933 22389 37967 22423
rect 41613 22389 41647 22423
rect 42625 22389 42659 22423
rect 1777 22185 1811 22219
rect 13369 22185 13403 22219
rect 40877 22185 40911 22219
rect 42717 22185 42751 22219
rect 43177 22185 43211 22219
rect 2881 22117 2915 22151
rect 32873 22117 32907 22151
rect 36185 22049 36219 22083
rect 1593 21981 1627 22015
rect 16957 21981 16991 22015
rect 17601 21981 17635 22015
rect 20361 21981 20395 22015
rect 21005 21981 21039 22015
rect 33885 21981 33919 22015
rect 34069 21981 34103 22015
rect 38853 21981 38887 22015
rect 39037 21981 39071 22015
rect 41337 21981 41371 22015
rect 41604 21981 41638 22015
rect 43361 21981 43395 22015
rect 43453 21981 43487 22015
rect 13323 21947 13357 21981
rect 13553 21913 13587 21947
rect 36452 21913 36486 21947
rect 38025 21913 38059 21947
rect 38209 21913 38243 21947
rect 43177 21913 43211 21947
rect 4537 21845 4571 21879
rect 13185 21845 13219 21879
rect 14381 21845 14415 21879
rect 33977 21845 34011 21879
rect 37565 21845 37599 21879
rect 38393 21845 38427 21879
rect 39221 21845 39255 21879
rect 43637 21845 43671 21879
rect 2881 21641 2915 21675
rect 38853 21641 38887 21675
rect 44005 21641 44039 21675
rect 17132 21573 17166 21607
rect 20352 21573 20386 21607
rect 36921 21573 36955 21607
rect 4353 21505 4387 21539
rect 16865 21505 16899 21539
rect 18705 21505 18739 21539
rect 18981 21505 19015 21539
rect 28457 21505 28491 21539
rect 29173 21505 29207 21539
rect 30757 21505 30791 21539
rect 31033 21505 31067 21539
rect 33425 21505 33459 21539
rect 33692 21505 33726 21539
rect 35449 21505 35483 21539
rect 35725 21505 35759 21539
rect 37473 21505 37507 21539
rect 37740 21505 37774 21539
rect 40426 21505 40460 21539
rect 40693 21505 40727 21539
rect 42625 21505 42659 21539
rect 42892 21505 42926 21539
rect 18797 21437 18831 21471
rect 20085 21437 20119 21471
rect 28917 21437 28951 21471
rect 30849 21437 30883 21471
rect 35633 21437 35667 21471
rect 18245 21369 18279 21403
rect 31217 21369 31251 21403
rect 34805 21369 34839 21403
rect 36645 21369 36679 21403
rect 2145 21301 2179 21335
rect 4997 21301 5031 21335
rect 16313 21301 16347 21335
rect 18705 21301 18739 21335
rect 19165 21301 19199 21335
rect 21465 21301 21499 21335
rect 22017 21301 22051 21335
rect 30297 21301 30331 21335
rect 30757 21301 30791 21335
rect 31769 21301 31803 21335
rect 32505 21301 32539 21335
rect 35265 21301 35299 21335
rect 35449 21301 35483 21335
rect 36461 21301 36495 21335
rect 39313 21301 39347 21335
rect 41153 21301 41187 21335
rect 3985 21097 4019 21131
rect 18061 21097 18095 21131
rect 22109 21097 22143 21131
rect 29193 21097 29227 21131
rect 34161 21097 34195 21131
rect 36277 21097 36311 21131
rect 37565 21097 37599 21131
rect 38669 21097 38703 21131
rect 39405 21097 39439 21131
rect 41889 21097 41923 21131
rect 43729 21097 43763 21131
rect 3433 21029 3467 21063
rect 21649 21029 21683 21063
rect 4077 20961 4111 20995
rect 22201 20961 22235 20995
rect 38301 20961 38335 20995
rect 40509 20961 40543 20995
rect 42349 20961 42383 20995
rect 2053 20893 2087 20927
rect 4261 20893 4295 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 16681 20893 16715 20927
rect 19809 20893 19843 20927
rect 20269 20893 20303 20927
rect 20536 20893 20570 20927
rect 22385 20893 22419 20927
rect 27813 20893 27847 20927
rect 31861 20893 31895 20927
rect 32321 20893 32355 20927
rect 32588 20893 32622 20927
rect 34897 20893 34931 20927
rect 36737 20893 36771 20927
rect 38393 20893 38427 20927
rect 39221 20893 39255 20927
rect 40776 20893 40810 20927
rect 42616 20893 42650 20927
rect 2298 20825 2332 20859
rect 3985 20825 4019 20859
rect 16948 20825 16982 20859
rect 22109 20825 22143 20859
rect 28080 20825 28114 20859
rect 30113 20825 30147 20859
rect 35164 20825 35198 20859
rect 37381 20825 37415 20859
rect 37597 20825 37631 20859
rect 4445 20757 4479 20791
rect 22569 20757 22603 20791
rect 33701 20757 33735 20791
rect 37749 20757 37783 20791
rect 3985 20553 4019 20587
rect 4445 20553 4479 20587
rect 15669 20553 15703 20587
rect 21465 20553 21499 20587
rect 29377 20553 29411 20587
rect 31309 20553 31343 20587
rect 33977 20553 34011 20587
rect 34621 20553 34655 20587
rect 36645 20553 36679 20587
rect 37749 20553 37783 20587
rect 2872 20485 2906 20519
rect 5558 20485 5592 20519
rect 17110 20485 17144 20519
rect 18797 20485 18831 20519
rect 32864 20485 32898 20519
rect 35756 20485 35790 20519
rect 39129 20485 39163 20519
rect 2145 20417 2179 20451
rect 2605 20417 2639 20451
rect 13369 20417 13403 20451
rect 13636 20417 13670 20451
rect 15209 20417 15243 20451
rect 15485 20417 15519 20451
rect 16865 20417 16899 20451
rect 19073 20417 19107 20451
rect 20341 20417 20375 20451
rect 27997 20417 28031 20451
rect 28264 20417 28298 20451
rect 29929 20417 29963 20451
rect 30185 20417 30219 20451
rect 36001 20417 36035 20451
rect 36829 20417 36863 20451
rect 37933 20417 37967 20451
rect 5825 20349 5859 20383
rect 15301 20349 15335 20383
rect 18981 20349 19015 20383
rect 20085 20349 20119 20383
rect 32597 20349 32631 20383
rect 18245 20281 18279 20315
rect 39405 20281 39439 20315
rect 12725 20213 12759 20247
rect 14749 20213 14783 20247
rect 15209 20213 15243 20247
rect 19073 20213 19107 20247
rect 19257 20213 19291 20247
rect 39589 20213 39623 20247
rect 3433 20009 3467 20043
rect 13737 20009 13771 20043
rect 15669 20009 15703 20043
rect 17969 20009 18003 20043
rect 21557 20009 21591 20043
rect 28273 20009 28307 20043
rect 30021 20009 30055 20043
rect 30481 20009 30515 20043
rect 33517 20009 33551 20043
rect 33701 20009 33735 20043
rect 35081 20009 35115 20043
rect 14289 19873 14323 19907
rect 33425 19873 33459 19907
rect 2053 19805 2087 19839
rect 2320 19805 2354 19839
rect 12357 19805 12391 19839
rect 16589 19805 16623 19839
rect 20177 19805 20211 19839
rect 20444 19805 20478 19839
rect 32137 19805 32171 19839
rect 33241 19805 33275 19839
rect 33517 19805 33551 19839
rect 12624 19737 12658 19771
rect 14556 19737 14590 19771
rect 16834 19737 16868 19771
rect 18429 19669 18463 19703
rect 14749 19465 14783 19499
rect 33701 19465 33735 19499
rect 32566 19397 32600 19431
rect 6561 19329 6595 19363
rect 6817 19329 6851 19363
rect 13369 19329 13403 19363
rect 13636 19329 13670 19363
rect 18521 19329 18555 19363
rect 32321 19329 32355 19363
rect 6009 19261 6043 19295
rect 2513 19125 2547 19159
rect 7941 19125 7975 19159
rect 17417 19125 17451 19159
rect 19993 19125 20027 19159
rect 37841 19125 37875 19159
rect 40969 19125 41003 19159
rect 41797 19125 41831 19159
rect 3433 18921 3467 18955
rect 3985 18921 4019 18955
rect 7389 18921 7423 18955
rect 14473 18921 14507 18955
rect 2053 18785 2087 18819
rect 4077 18785 4111 18819
rect 2320 18717 2354 18751
rect 4261 18717 4295 18751
rect 5641 18717 5675 18751
rect 7113 18717 7147 18751
rect 7205 18717 7239 18751
rect 16773 18717 16807 18751
rect 18613 18717 18647 18751
rect 20913 18717 20947 18751
rect 21097 18717 21131 18751
rect 37105 18717 37139 18751
rect 37565 18717 37599 18751
rect 40693 18717 40727 18751
rect 40960 18717 40994 18751
rect 44465 18717 44499 18751
rect 3985 18649 4019 18683
rect 7389 18649 7423 18683
rect 17018 18649 17052 18683
rect 37832 18649 37866 18683
rect 4445 18581 4479 18615
rect 6929 18581 6963 18615
rect 18153 18581 18187 18615
rect 21005 18581 21039 18615
rect 38945 18581 38979 18615
rect 42073 18581 42107 18615
rect 3525 18377 3559 18411
rect 7941 18377 7975 18411
rect 19257 18377 19291 18411
rect 18797 18309 18831 18343
rect 44456 18309 44490 18343
rect 2145 18241 2179 18275
rect 2401 18241 2435 18275
rect 4629 18241 4663 18275
rect 4813 18241 4847 18275
rect 6561 18241 6595 18275
rect 6817 18241 6851 18275
rect 16313 18241 16347 18275
rect 17213 18241 17247 18275
rect 19073 18241 19107 18275
rect 20352 18241 20386 18275
rect 22017 18241 22051 18275
rect 22109 18241 22143 18275
rect 22293 18241 22327 18275
rect 37740 18241 37774 18275
rect 39313 18241 39347 18275
rect 40693 18241 40727 18275
rect 40960 18241 40994 18275
rect 42625 18241 42659 18275
rect 42901 18241 42935 18275
rect 6009 18173 6043 18207
rect 16957 18173 16991 18207
rect 18889 18173 18923 18207
rect 20085 18173 20119 18207
rect 37473 18173 37507 18207
rect 42717 18173 42751 18207
rect 44189 18173 44223 18207
rect 42073 18105 42107 18139
rect 3985 18037 4019 18071
rect 4629 18037 4663 18071
rect 4997 18037 5031 18071
rect 8401 18037 8435 18071
rect 18337 18037 18371 18071
rect 18797 18037 18831 18071
rect 21465 18037 21499 18071
rect 22293 18037 22327 18071
rect 36921 18037 36955 18071
rect 38853 18037 38887 18071
rect 40233 18037 40267 18071
rect 42625 18037 42659 18071
rect 43085 18037 43119 18071
rect 45569 18037 45603 18071
rect 3433 17833 3467 17867
rect 6561 17833 6595 17867
rect 17049 17833 17083 17867
rect 18889 17833 18923 17867
rect 38761 17833 38795 17867
rect 43361 17833 43395 17867
rect 22937 17765 22971 17799
rect 2053 17697 2087 17731
rect 38853 17697 38887 17731
rect 43453 17697 43487 17731
rect 2320 17629 2354 17663
rect 4169 17629 4203 17663
rect 7941 17629 7975 17663
rect 14657 17629 14691 17663
rect 17509 17629 17543 17663
rect 19717 17629 19751 17663
rect 21557 17629 21591 17663
rect 36645 17629 36679 17663
rect 38945 17629 38979 17663
rect 43637 17629 43671 17663
rect 44649 17629 44683 17663
rect 45201 17629 45235 17663
rect 7696 17561 7730 17595
rect 17776 17561 17810 17595
rect 19984 17561 20018 17595
rect 21802 17561 21836 17595
rect 36912 17561 36946 17595
rect 38669 17561 38703 17595
rect 40693 17561 40727 17595
rect 41153 17561 41187 17595
rect 42901 17561 42935 17595
rect 43361 17561 43395 17595
rect 5457 17493 5491 17527
rect 21097 17493 21131 17527
rect 38025 17493 38059 17527
rect 39129 17493 39163 17527
rect 43821 17493 43855 17527
rect 3985 17289 4019 17323
rect 18429 17289 18463 17323
rect 20821 17289 20855 17323
rect 22227 17289 22261 17323
rect 38853 17289 38887 17323
rect 41613 17289 41647 17323
rect 46765 17289 46799 17323
rect 4896 17221 4930 17255
rect 14648 17221 14682 17255
rect 17316 17221 17350 17255
rect 22017 17221 22051 17255
rect 37718 17221 37752 17255
rect 42892 17221 42926 17255
rect 44732 17221 44766 17255
rect 2605 17153 2639 17187
rect 2872 17153 2906 17187
rect 4629 17153 4663 17187
rect 17049 17153 17083 17187
rect 21189 17153 21223 17187
rect 37473 17153 37507 17187
rect 40233 17153 40267 17187
rect 40489 17153 40523 17187
rect 44465 17153 44499 17187
rect 46305 17153 46339 17187
rect 46581 17153 46615 17187
rect 2145 17085 2179 17119
rect 14381 17085 14415 17119
rect 21097 17085 21131 17119
rect 42625 17085 42659 17119
rect 46397 17085 46431 17119
rect 6009 17017 6043 17051
rect 44005 17017 44039 17051
rect 45845 17017 45879 17051
rect 6561 16949 6595 16983
rect 15761 16949 15795 16983
rect 22201 16949 22235 16983
rect 22385 16949 22419 16983
rect 46305 16949 46339 16983
rect 3985 16745 4019 16779
rect 16129 16745 16163 16779
rect 20729 16745 20763 16779
rect 21557 16745 21591 16779
rect 40969 16745 41003 16779
rect 46581 16745 46615 16779
rect 21465 16677 21499 16711
rect 13737 16609 13771 16643
rect 16221 16609 16255 16643
rect 43177 16609 43211 16643
rect 45201 16609 45235 16643
rect 14289 16541 14323 16575
rect 16405 16541 16439 16575
rect 20729 16541 20763 16575
rect 20913 16541 20947 16575
rect 21373 16541 21407 16575
rect 41429 16541 41463 16575
rect 44465 16541 44499 16575
rect 45457 16541 45491 16575
rect 14534 16473 14568 16507
rect 16129 16473 16163 16507
rect 21649 16473 21683 16507
rect 15669 16405 15703 16439
rect 16589 16405 16623 16439
rect 15945 16201 15979 16235
rect 41245 16201 41279 16235
rect 45477 16201 45511 16235
rect 14810 16133 14844 16167
rect 19441 16133 19475 16167
rect 19625 16133 19659 16167
rect 44364 16133 44398 16167
rect 8769 16065 8803 16099
rect 14105 16065 14139 16099
rect 19717 16065 19751 16099
rect 20177 16065 20211 16099
rect 20361 16065 20395 16099
rect 44097 16065 44131 16099
rect 14565 15997 14599 16031
rect 8953 15861 8987 15895
rect 16865 15861 16899 15895
rect 19441 15861 19475 15895
rect 20269 15861 20303 15895
rect 40141 15861 40175 15895
rect 40601 15861 40635 15895
rect 7849 15657 7883 15691
rect 16497 15657 16531 15691
rect 20085 15657 20119 15691
rect 41429 15657 41463 15691
rect 41889 15657 41923 15691
rect 42349 15657 42383 15691
rect 40049 15521 40083 15555
rect 41981 15521 42015 15555
rect 10250 15453 10284 15487
rect 10517 15453 10551 15487
rect 15117 15453 15151 15487
rect 15384 15453 15418 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 19901 15453 19935 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 22845 15453 22879 15487
rect 39497 15453 39531 15487
rect 40316 15453 40350 15487
rect 42165 15453 42199 15487
rect 43729 15453 43763 15487
rect 8033 15385 8067 15419
rect 19717 15385 19751 15419
rect 19809 15385 19843 15419
rect 20729 15385 20763 15419
rect 20913 15385 20947 15419
rect 21833 15385 21867 15419
rect 41889 15385 41923 15419
rect 7665 15317 7699 15351
rect 7833 15317 7867 15351
rect 9137 15317 9171 15351
rect 20545 15317 20579 15351
rect 22661 15317 22695 15351
rect 8953 15113 8987 15147
rect 18705 15113 18739 15147
rect 21465 15113 21499 15147
rect 23397 15113 23431 15147
rect 40693 15113 40727 15147
rect 9321 15045 9355 15079
rect 10057 15045 10091 15079
rect 11713 15045 11747 15079
rect 11913 15045 11947 15079
rect 19818 15045 19852 15079
rect 21281 15045 21315 15079
rect 22284 15045 22318 15079
rect 3525 14977 3559 15011
rect 3781 14977 3815 15011
rect 7113 14977 7147 15011
rect 7380 14977 7414 15011
rect 9137 14977 9171 15011
rect 9413 14977 9447 15011
rect 10241 14977 10275 15011
rect 12541 14977 12575 15011
rect 18245 14977 18279 15011
rect 20913 14977 20947 15011
rect 39580 14977 39614 15011
rect 43821 14977 43855 15011
rect 44088 14977 44122 15011
rect 20085 14909 20119 14943
rect 22017 14909 22051 14943
rect 39313 14909 39347 14943
rect 8493 14841 8527 14875
rect 12081 14841 12115 14875
rect 4905 14773 4939 14807
rect 9873 14773 9907 14807
rect 11897 14773 11931 14807
rect 13829 14773 13863 14807
rect 14841 14773 14875 14807
rect 18153 14773 18187 14807
rect 21281 14773 21315 14807
rect 41153 14773 41187 14807
rect 45201 14773 45235 14807
rect 3433 14569 3467 14603
rect 7573 14569 7607 14603
rect 9321 14569 9355 14603
rect 10793 14569 10827 14603
rect 17785 14569 17819 14603
rect 18889 14569 18923 14603
rect 21925 14569 21959 14603
rect 41429 14569 41463 14603
rect 45845 14569 45879 14603
rect 9137 14501 9171 14535
rect 17325 14501 17359 14535
rect 18153 14501 18187 14535
rect 19441 14501 19475 14535
rect 8585 14433 8619 14467
rect 17877 14433 17911 14467
rect 20821 14433 20855 14467
rect 3249 14365 3283 14399
rect 4445 14365 4479 14399
rect 4721 14365 4755 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 5733 14365 5767 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 10977 14365 11011 14399
rect 11253 14365 11287 14399
rect 13093 14365 13127 14399
rect 13737 14365 13771 14399
rect 14473 14365 14507 14399
rect 15485 14365 15519 14399
rect 15945 14365 15979 14399
rect 17785 14365 17819 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 21465 14365 21499 14399
rect 22109 14365 22143 14399
rect 22293 14365 22327 14399
rect 40049 14365 40083 14399
rect 40316 14365 40350 14399
rect 43269 14365 43303 14399
rect 45201 14365 45235 14399
rect 5365 14297 5399 14331
rect 9305 14297 9339 14331
rect 9505 14297 9539 14331
rect 12848 14297 12882 14331
rect 16190 14297 16224 14331
rect 20576 14297 20610 14331
rect 43536 14297 43570 14331
rect 4261 14229 4295 14263
rect 8217 14229 8251 14263
rect 11161 14229 11195 14263
rect 11713 14229 11747 14263
rect 13553 14229 13587 14263
rect 14289 14229 14323 14263
rect 21281 14229 21315 14263
rect 44649 14229 44683 14263
rect 4813 14025 4847 14059
rect 5365 14025 5399 14059
rect 5733 14025 5767 14059
rect 8033 14025 8067 14059
rect 8861 14025 8895 14059
rect 11161 14025 11195 14059
rect 12081 14025 12115 14059
rect 41429 14025 41463 14059
rect 45753 14025 45787 14059
rect 11069 13957 11103 13991
rect 11713 13957 11747 13991
rect 11929 13957 11963 13991
rect 13676 13957 13710 13991
rect 17693 13957 17727 13991
rect 18153 13957 18187 13991
rect 19901 13957 19935 13991
rect 40316 13957 40350 13991
rect 43720 13957 43754 13991
rect 3433 13889 3467 13923
rect 3700 13889 3734 13923
rect 5273 13889 5307 13923
rect 5549 13889 5583 13923
rect 7941 13889 7975 13923
rect 8125 13889 8159 13923
rect 8677 13889 8711 13923
rect 8861 13889 8895 13923
rect 10885 13889 10919 13923
rect 11161 13889 11195 13923
rect 13921 13889 13955 13923
rect 20821 13889 20855 13923
rect 20913 13889 20947 13923
rect 43453 13889 43487 13923
rect 45293 13889 45327 13923
rect 45569 13889 45603 13923
rect 20637 13821 20671 13855
rect 40049 13821 40083 13855
rect 45385 13821 45419 13855
rect 44833 13753 44867 13787
rect 11897 13685 11931 13719
rect 12541 13685 12575 13719
rect 16037 13685 16071 13719
rect 45293 13685 45327 13719
rect 12633 13481 12667 13515
rect 17141 13481 17175 13515
rect 19993 13481 20027 13515
rect 20177 13481 20211 13515
rect 44373 13481 44407 13515
rect 4169 13413 4203 13447
rect 12173 13413 12207 13447
rect 3985 13345 4019 13379
rect 15761 13345 15795 13379
rect 42993 13345 43027 13379
rect 4261 13277 4295 13311
rect 4813 13277 4847 13311
rect 5089 13277 5123 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 6561 13277 6595 13311
rect 7941 13277 7975 13311
rect 8217 13277 8251 13311
rect 10977 13277 11011 13311
rect 13001 13277 13035 13311
rect 16028 13277 16062 13311
rect 40049 13277 40083 13311
rect 8033 13209 8067 13243
rect 11989 13209 12023 13243
rect 12817 13209 12851 13243
rect 19809 13209 19843 13243
rect 20025 13209 20059 13243
rect 43260 13209 43294 13243
rect 4261 13141 4295 13175
rect 6561 13141 6595 13175
rect 8401 13141 8435 13175
rect 10793 13141 10827 13175
rect 11621 13141 11655 13175
rect 11805 13141 11839 13175
rect 11897 13141 11931 13175
rect 4629 12937 4663 12971
rect 7415 12937 7449 12971
rect 8309 12937 8343 12971
rect 11069 12937 11103 12971
rect 11713 12937 11747 12971
rect 12817 12937 12851 12971
rect 43269 12937 43303 12971
rect 43913 12937 43947 12971
rect 7205 12869 7239 12903
rect 8677 12869 8711 12903
rect 9321 12869 9355 12903
rect 10885 12869 10919 12903
rect 39396 12869 39430 12903
rect 43361 12869 43395 12903
rect 43821 12869 43855 12903
rect 44189 12869 44223 12903
rect 4813 12801 4847 12835
rect 4905 12801 4939 12835
rect 5089 12801 5123 12835
rect 5181 12807 5215 12841
rect 8401 12801 8435 12835
rect 8493 12801 8527 12835
rect 9137 12801 9171 12835
rect 10517 12801 10551 12835
rect 12173 12801 12207 12835
rect 12725 12801 12759 12835
rect 12909 12801 12943 12835
rect 42993 12801 43027 12835
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 39129 12733 39163 12767
rect 7573 12665 7607 12699
rect 44097 12665 44131 12699
rect 7389 12597 7423 12631
rect 8125 12597 8159 12631
rect 9505 12597 9539 12631
rect 10885 12597 10919 12631
rect 40509 12597 40543 12631
rect 43085 12597 43119 12631
rect 43177 12597 43211 12631
rect 44005 12597 44039 12631
rect 8585 12393 8619 12427
rect 9321 12393 9355 12427
rect 11897 12393 11931 12427
rect 9689 12325 9723 12359
rect 3985 12189 4019 12223
rect 7205 12189 7239 12223
rect 10517 12189 10551 12223
rect 10784 12189 10818 12223
rect 38853 12189 38887 12223
rect 39313 12189 39347 12223
rect 42901 12189 42935 12223
rect 7450 12121 7484 12155
rect 9321 12121 9355 12155
rect 9137 12053 9171 12087
rect 41613 12053 41647 12087
rect 6561 11849 6595 11883
rect 7297 11849 7331 11883
rect 9137 11849 9171 11883
rect 9597 11849 9631 11883
rect 41337 11849 41371 11883
rect 8024 11781 8058 11815
rect 12173 11781 12207 11815
rect 39304 11781 39338 11815
rect 2964 11713 2998 11747
rect 4629 11713 4663 11747
rect 7113 11713 7147 11747
rect 7757 11713 7791 11747
rect 9781 11713 9815 11747
rect 39037 11713 39071 11747
rect 40877 11713 40911 11747
rect 41153 11713 41187 11747
rect 2697 11645 2731 11679
rect 40969 11645 41003 11679
rect 4077 11577 4111 11611
rect 11805 11577 11839 11611
rect 40417 11577 40451 11611
rect 2237 11509 2271 11543
rect 11713 11509 11747 11543
rect 38393 11509 38427 11543
rect 40877 11509 40911 11543
rect 42625 11509 42659 11543
rect 43453 11509 43487 11543
rect 12725 11305 12759 11339
rect 39497 11305 39531 11339
rect 41429 11305 41463 11339
rect 43545 11305 43579 11339
rect 44005 11305 44039 11339
rect 44465 11305 44499 11339
rect 6561 11169 6595 11203
rect 11345 11169 11379 11203
rect 1961 11101 1995 11135
rect 6101 11101 6135 11135
rect 20361 11101 20395 11135
rect 38117 11101 38151 11135
rect 40049 11101 40083 11135
rect 42165 11101 42199 11135
rect 44189 11101 44223 11135
rect 44281 11101 44315 11135
rect 2228 11033 2262 11067
rect 4353 11033 4387 11067
rect 6806 11033 6840 11067
rect 11612 11033 11646 11067
rect 38384 11033 38418 11067
rect 40294 11033 40328 11067
rect 42432 11033 42466 11067
rect 44005 11033 44039 11067
rect 3341 10965 3375 10999
rect 7941 10965 7975 10999
rect 20177 10965 20211 10999
rect 6653 10761 6687 10795
rect 8309 10761 8343 10795
rect 11713 10761 11747 10795
rect 44005 10761 44039 10795
rect 45845 10761 45879 10795
rect 8125 10693 8159 10727
rect 44732 10693 44766 10727
rect 1593 10625 1627 10659
rect 1860 10625 1894 10659
rect 3433 10625 3467 10659
rect 3700 10625 3734 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 7757 10625 7791 10659
rect 11897 10625 11931 10659
rect 40141 10625 40175 10659
rect 42625 10625 42659 10659
rect 42881 10625 42915 10659
rect 42073 10557 42107 10591
rect 44465 10557 44499 10591
rect 2973 10421 3007 10455
rect 4813 10421 4847 10455
rect 5733 10421 5767 10455
rect 6837 10421 6871 10455
rect 8125 10421 8159 10455
rect 40325 10421 40359 10455
rect 4077 10217 4111 10251
rect 4537 10217 4571 10251
rect 6837 10217 6871 10251
rect 43913 10217 43947 10251
rect 2973 10081 3007 10115
rect 4261 10081 4295 10115
rect 5457 10081 5491 10115
rect 19993 10081 20027 10115
rect 42533 10081 42567 10115
rect 45201 10081 45235 10115
rect 4077 10013 4111 10047
rect 4353 10013 4387 10047
rect 5724 10013 5758 10047
rect 20260 10013 20294 10047
rect 45457 10013 45491 10047
rect 2728 9945 2762 9979
rect 42800 9945 42834 9979
rect 1593 9877 1627 9911
rect 21373 9877 21407 9911
rect 46581 9877 46615 9911
rect 2789 9537 2823 9571
rect 5733 9537 5767 9571
rect 40509 9537 40543 9571
rect 40765 9537 40799 9571
rect 42809 9537 42843 9571
rect 41889 9333 41923 9367
rect 57529 3689 57563 3723
rect 58081 3485 58115 3519
rect 58265 3349 58299 3383
rect 1869 2397 1903 2431
rect 22017 2397 22051 2431
rect 42625 2397 42659 2431
rect 1685 2261 1719 2295
rect 22201 2261 22235 2295
rect 42809 2261 42843 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 6454 57536 6460 57588
rect 6512 57576 6518 57588
rect 6641 57579 6699 57585
rect 6641 57576 6653 57579
rect 6512 57548 6653 57576
rect 6512 57536 6518 57548
rect 6641 57545 6653 57548
rect 6687 57545 6699 57579
rect 6641 57539 6699 57545
rect 28350 57536 28356 57588
rect 28408 57576 28414 57588
rect 28537 57579 28595 57585
rect 28537 57576 28549 57579
rect 28408 57548 28549 57576
rect 28408 57536 28414 57548
rect 28537 57545 28549 57548
rect 28583 57545 28595 57579
rect 28537 57539 28595 57545
rect 49694 57536 49700 57588
rect 49752 57576 49758 57588
rect 50525 57579 50583 57585
rect 50525 57576 50537 57579
rect 49752 57548 50537 57576
rect 49752 57536 49758 57548
rect 50525 57545 50537 57548
rect 50571 57545 50583 57579
rect 50525 57539 50583 57545
rect 6638 57400 6644 57452
rect 6696 57440 6702 57452
rect 6825 57443 6883 57449
rect 6825 57440 6837 57443
rect 6696 57412 6837 57440
rect 6696 57400 6702 57412
rect 6825 57409 6837 57412
rect 6871 57409 6883 57443
rect 6825 57403 6883 57409
rect 28534 57400 28540 57452
rect 28592 57440 28598 57452
rect 28721 57443 28779 57449
rect 28721 57440 28733 57443
rect 28592 57412 28733 57440
rect 28592 57400 28598 57412
rect 28721 57409 28733 57412
rect 28767 57409 28779 57443
rect 28721 57403 28779 57409
rect 46566 57400 46572 57452
rect 46624 57440 46630 57452
rect 50341 57443 50399 57449
rect 50341 57440 50353 57443
rect 46624 57412 50353 57440
rect 46624 57400 46630 57412
rect 50341 57409 50353 57412
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 45554 49172 45560 49224
rect 45612 49212 45618 49224
rect 58069 49215 58127 49221
rect 58069 49212 58081 49215
rect 45612 49184 58081 49212
rect 45612 49172 45618 49184
rect 58069 49181 58081 49184
rect 58115 49181 58127 49215
rect 58069 49175 58127 49181
rect 58250 49076 58256 49088
rect 58211 49048 58256 49076
rect 58250 49036 58256 49048
rect 58308 49036 58314 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 6638 46152 6644 46164
rect 6599 46124 6644 46152
rect 6638 46112 6644 46124
rect 6696 46112 6702 46164
rect 46566 46152 46572 46164
rect 46527 46124 46572 46152
rect 46566 46112 46572 46124
rect 46624 46112 46630 46164
rect 5261 45951 5319 45957
rect 5261 45917 5273 45951
rect 5307 45948 5319 45951
rect 6730 45948 6736 45960
rect 5307 45920 6736 45948
rect 5307 45917 5319 45920
rect 5261 45911 5319 45917
rect 6730 45908 6736 45920
rect 6788 45908 6794 45960
rect 40494 45948 40500 45960
rect 40455 45920 40500 45948
rect 40494 45908 40500 45920
rect 40552 45908 40558 45960
rect 44266 45908 44272 45960
rect 44324 45948 44330 45960
rect 45189 45951 45247 45957
rect 45189 45948 45201 45951
rect 44324 45920 45201 45948
rect 44324 45908 44330 45920
rect 45189 45917 45201 45920
rect 45235 45917 45247 45951
rect 45189 45911 45247 45917
rect 5528 45883 5586 45889
rect 5528 45849 5540 45883
rect 5574 45880 5586 45883
rect 5810 45880 5816 45892
rect 5574 45852 5816 45880
rect 5574 45849 5586 45852
rect 5528 45843 5586 45849
rect 5810 45840 5816 45852
rect 5868 45840 5874 45892
rect 45456 45883 45514 45889
rect 45456 45849 45468 45883
rect 45502 45880 45514 45883
rect 45830 45880 45836 45892
rect 45502 45852 45836 45880
rect 45502 45849 45514 45852
rect 45456 45843 45514 45849
rect 45830 45840 45836 45852
rect 45888 45840 45894 45892
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 5810 45608 5816 45620
rect 5771 45580 5816 45608
rect 5810 45568 5816 45580
rect 5868 45568 5874 45620
rect 8849 45611 8907 45617
rect 8849 45577 8861 45611
rect 8895 45608 8907 45611
rect 8895 45580 8929 45608
rect 8895 45577 8907 45580
rect 8849 45571 8907 45577
rect 8864 45540 8892 45571
rect 9122 45540 9128 45552
rect 8864 45512 9128 45540
rect 9122 45500 9128 45512
rect 9180 45540 9186 45552
rect 9493 45543 9551 45549
rect 9493 45540 9505 45543
rect 9180 45512 9505 45540
rect 9180 45500 9186 45512
rect 9493 45509 9505 45512
rect 9539 45509 9551 45543
rect 28994 45540 29000 45552
rect 9493 45503 9551 45509
rect 27172 45512 29000 45540
rect 5997 45475 6055 45481
rect 5997 45441 6009 45475
rect 6043 45441 6055 45475
rect 5997 45435 6055 45441
rect 6733 45475 6791 45481
rect 6733 45441 6745 45475
rect 6779 45472 6791 45475
rect 7098 45472 7104 45484
rect 6779 45444 7104 45472
rect 6779 45441 6791 45444
rect 6733 45435 6791 45441
rect 6012 45404 6040 45435
rect 7098 45432 7104 45444
rect 7156 45432 7162 45484
rect 7736 45475 7794 45481
rect 7736 45441 7748 45475
rect 7782 45472 7794 45475
rect 8294 45472 8300 45484
rect 7782 45444 8300 45472
rect 7782 45441 7794 45444
rect 7736 45435 7794 45441
rect 8294 45432 8300 45444
rect 8352 45432 8358 45484
rect 9674 45472 9680 45484
rect 9635 45444 9680 45472
rect 9674 45432 9680 45444
rect 9732 45432 9738 45484
rect 27172 45481 27200 45512
rect 28994 45500 29000 45512
rect 29052 45500 29058 45552
rect 40396 45543 40454 45549
rect 40396 45509 40408 45543
rect 40442 45540 40454 45543
rect 40494 45540 40500 45552
rect 40442 45512 40500 45540
rect 40442 45509 40454 45512
rect 40396 45503 40454 45509
rect 40494 45500 40500 45512
rect 40552 45500 40558 45552
rect 27157 45475 27215 45481
rect 27157 45441 27169 45475
rect 27203 45441 27215 45475
rect 27157 45435 27215 45441
rect 27246 45432 27252 45484
rect 27304 45472 27310 45484
rect 27413 45475 27471 45481
rect 27413 45472 27425 45475
rect 27304 45444 27425 45472
rect 27304 45432 27310 45444
rect 27413 45441 27425 45444
rect 27459 45441 27471 45475
rect 27413 45435 27471 45441
rect 44177 45475 44235 45481
rect 44177 45441 44189 45475
rect 44223 45472 44235 45475
rect 44266 45472 44272 45484
rect 44223 45444 44272 45472
rect 44223 45441 44235 45444
rect 44177 45435 44235 45441
rect 44266 45432 44272 45444
rect 44324 45432 44330 45484
rect 44450 45481 44456 45484
rect 44444 45435 44456 45481
rect 44508 45472 44514 45484
rect 44508 45444 44544 45472
rect 44450 45432 44456 45435
rect 44508 45432 44514 45444
rect 7374 45404 7380 45416
rect 6012 45376 7380 45404
rect 7374 45364 7380 45376
rect 7432 45364 7438 45416
rect 7469 45407 7527 45413
rect 7469 45373 7481 45407
rect 7515 45373 7527 45407
rect 40126 45404 40132 45416
rect 40087 45376 40132 45404
rect 7469 45367 7527 45373
rect 6730 45296 6736 45348
rect 6788 45336 6794 45348
rect 6914 45336 6920 45348
rect 6788 45308 6920 45336
rect 6788 45296 6794 45308
rect 6914 45296 6920 45308
rect 6972 45336 6978 45348
rect 7484 45336 7512 45367
rect 40126 45364 40132 45376
rect 40184 45364 40190 45416
rect 28534 45336 28540 45348
rect 6972 45308 7512 45336
rect 28495 45308 28540 45336
rect 6972 45296 6978 45308
rect 28534 45296 28540 45308
rect 28592 45296 28598 45348
rect 45554 45296 45560 45348
rect 45612 45336 45618 45348
rect 45612 45308 45657 45336
rect 45612 45296 45618 45308
rect 6454 45228 6460 45280
rect 6512 45268 6518 45280
rect 6549 45271 6607 45277
rect 6549 45268 6561 45271
rect 6512 45240 6561 45268
rect 6512 45228 6518 45240
rect 6549 45237 6561 45240
rect 6595 45237 6607 45271
rect 6549 45231 6607 45237
rect 7650 45228 7656 45280
rect 7708 45268 7714 45280
rect 9309 45271 9367 45277
rect 9309 45268 9321 45271
rect 7708 45240 9321 45268
rect 7708 45228 7714 45240
rect 9309 45237 9321 45240
rect 9355 45237 9367 45271
rect 9309 45231 9367 45237
rect 37645 45271 37703 45277
rect 37645 45237 37657 45271
rect 37691 45268 37703 45271
rect 37734 45268 37740 45280
rect 37691 45240 37740 45268
rect 37691 45237 37703 45240
rect 37645 45231 37703 45237
rect 37734 45228 37740 45240
rect 37792 45228 37798 45280
rect 41506 45268 41512 45280
rect 41467 45240 41512 45268
rect 41506 45228 41512 45240
rect 41564 45228 41570 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 7650 45064 7656 45076
rect 7611 45036 7656 45064
rect 7650 45024 7656 45036
rect 7708 45024 7714 45076
rect 8294 45064 8300 45076
rect 8255 45036 8300 45064
rect 8294 45024 8300 45036
rect 8352 45024 8358 45076
rect 9030 45024 9036 45076
rect 9088 45064 9094 45076
rect 9861 45067 9919 45073
rect 9861 45064 9873 45067
rect 9088 45036 9873 45064
rect 9088 45024 9094 45036
rect 9861 45033 9873 45036
rect 9907 45033 9919 45067
rect 45830 45064 45836 45076
rect 45791 45036 45836 45064
rect 9861 45027 9919 45033
rect 6730 44928 6736 44940
rect 6691 44900 6736 44928
rect 6730 44888 6736 44900
rect 6788 44888 6794 44940
rect 9876 44928 9904 45027
rect 45830 45024 45836 45036
rect 45888 45024 45894 45076
rect 10778 44996 10784 45008
rect 10739 44968 10784 44996
rect 10778 44956 10784 44968
rect 10836 44956 10842 45008
rect 43809 44999 43867 45005
rect 43809 44965 43821 44999
rect 43855 44996 43867 44999
rect 44358 44996 44364 45008
rect 43855 44968 44364 44996
rect 43855 44965 43867 44968
rect 43809 44959 43867 44965
rect 44358 44956 44364 44968
rect 44416 44956 44422 45008
rect 43625 44931 43683 44937
rect 9876 44900 10824 44928
rect 6454 44820 6460 44872
rect 6512 44869 6518 44872
rect 6512 44860 6524 44869
rect 6512 44832 6557 44860
rect 6512 44823 6524 44832
rect 6512 44820 6518 44823
rect 6822 44820 6828 44872
rect 6880 44860 6886 44872
rect 7282 44860 7288 44872
rect 6880 44832 7288 44860
rect 6880 44820 6886 44832
rect 7282 44820 7288 44832
rect 7340 44820 7346 44872
rect 10796 44869 10824 44900
rect 43625 44897 43637 44931
rect 43671 44897 43683 44931
rect 43625 44891 43683 44897
rect 8481 44863 8539 44869
rect 8481 44860 8493 44863
rect 7852 44832 8493 44860
rect 5353 44727 5411 44733
rect 5353 44693 5365 44727
rect 5399 44724 5411 44727
rect 5902 44724 5908 44736
rect 5399 44696 5908 44724
rect 5399 44693 5411 44696
rect 5353 44687 5411 44693
rect 5902 44684 5908 44696
rect 5960 44684 5966 44736
rect 7006 44684 7012 44736
rect 7064 44724 7070 44736
rect 7852 44733 7880 44832
rect 8481 44829 8493 44832
rect 8527 44829 8539 44863
rect 10505 44863 10563 44869
rect 10505 44860 10517 44863
rect 8481 44823 8539 44829
rect 9876 44832 10517 44860
rect 7653 44727 7711 44733
rect 7653 44724 7665 44727
rect 7064 44696 7665 44724
rect 7064 44684 7070 44696
rect 7653 44693 7665 44696
rect 7699 44693 7711 44727
rect 7653 44687 7711 44693
rect 7837 44727 7895 44733
rect 7837 44693 7849 44727
rect 7883 44693 7895 44727
rect 9674 44724 9680 44736
rect 9635 44696 9680 44724
rect 7837 44687 7895 44693
rect 9674 44684 9680 44696
rect 9732 44684 9738 44736
rect 9876 44733 9904 44832
rect 10505 44829 10517 44832
rect 10551 44829 10563 44863
rect 10505 44823 10563 44829
rect 10781 44863 10839 44869
rect 10781 44829 10793 44863
rect 10827 44860 10839 44863
rect 11146 44860 11152 44872
rect 10827 44832 11152 44860
rect 10827 44829 10839 44832
rect 10781 44823 10839 44829
rect 11146 44820 11152 44832
rect 11204 44820 11210 44872
rect 36909 44863 36967 44869
rect 36909 44829 36921 44863
rect 36955 44860 36967 44863
rect 36955 44832 37320 44860
rect 36955 44829 36967 44832
rect 36909 44823 36967 44829
rect 37292 44804 37320 44832
rect 40126 44820 40132 44872
rect 40184 44860 40190 44872
rect 40221 44863 40279 44869
rect 40221 44860 40233 44863
rect 40184 44832 40233 44860
rect 40184 44820 40190 44832
rect 40221 44829 40233 44832
rect 40267 44860 40279 44863
rect 41046 44860 41052 44872
rect 40267 44832 41052 44860
rect 40267 44829 40279 44832
rect 40221 44823 40279 44829
rect 41046 44820 41052 44832
rect 41104 44820 41110 44872
rect 42061 44863 42119 44869
rect 42061 44829 42073 44863
rect 42107 44829 42119 44863
rect 42061 44823 42119 44829
rect 42981 44863 43039 44869
rect 42981 44829 42993 44863
rect 43027 44860 43039 44863
rect 43640 44860 43668 44891
rect 43027 44832 43668 44860
rect 45373 44863 45431 44869
rect 43027 44829 43039 44832
rect 42981 44823 43039 44829
rect 45373 44829 45385 44863
rect 45419 44829 45431 44863
rect 45373 44823 45431 44829
rect 10042 44792 10048 44804
rect 10003 44764 10048 44792
rect 10042 44752 10048 44764
rect 10100 44792 10106 44804
rect 10597 44795 10655 44801
rect 10597 44792 10609 44795
rect 10100 44764 10609 44792
rect 10100 44752 10106 44764
rect 10597 44761 10609 44764
rect 10643 44761 10655 44795
rect 10597 44755 10655 44761
rect 36262 44752 36268 44804
rect 36320 44792 36326 44804
rect 37154 44795 37212 44801
rect 37154 44792 37166 44795
rect 36320 44764 37166 44792
rect 36320 44752 36326 44764
rect 37154 44761 37166 44764
rect 37200 44761 37212 44795
rect 37154 44755 37212 44761
rect 37274 44752 37280 44804
rect 37332 44752 37338 44804
rect 40488 44795 40546 44801
rect 40488 44761 40500 44795
rect 40534 44792 40546 44795
rect 42076 44792 42104 44823
rect 40534 44764 42104 44792
rect 40534 44761 40546 44764
rect 40488 44755 40546 44761
rect 43990 44752 43996 44804
rect 44048 44792 44054 44804
rect 44085 44795 44143 44801
rect 44085 44792 44097 44795
rect 44048 44764 44097 44792
rect 44048 44752 44054 44764
rect 44085 44761 44097 44764
rect 44131 44761 44143 44795
rect 45388 44792 45416 44823
rect 45462 44820 45468 44872
rect 45520 44860 45526 44872
rect 46017 44863 46075 44869
rect 46017 44860 46029 44863
rect 45520 44832 46029 44860
rect 45520 44820 45526 44832
rect 46017 44829 46029 44832
rect 46063 44829 46075 44863
rect 46017 44823 46075 44829
rect 45554 44792 45560 44804
rect 45388 44764 45560 44792
rect 44085 44755 44143 44761
rect 45554 44752 45560 44764
rect 45612 44752 45618 44804
rect 9845 44727 9904 44733
rect 9845 44693 9857 44727
rect 9891 44724 9904 44727
rect 9950 44724 9956 44736
rect 9891 44696 9956 44724
rect 9891 44693 9903 44696
rect 9845 44687 9903 44693
rect 9950 44684 9956 44696
rect 10008 44684 10014 44736
rect 38289 44727 38347 44733
rect 38289 44693 38301 44727
rect 38335 44724 38347 44727
rect 38470 44724 38476 44736
rect 38335 44696 38476 44724
rect 38335 44693 38347 44696
rect 38289 44687 38347 44693
rect 38470 44684 38476 44696
rect 38528 44684 38534 44736
rect 41601 44727 41659 44733
rect 41601 44693 41613 44727
rect 41647 44724 41659 44727
rect 42150 44724 42156 44736
rect 41647 44696 42156 44724
rect 41647 44693 41659 44696
rect 41601 44687 41659 44693
rect 42150 44684 42156 44696
rect 42208 44684 42214 44736
rect 43162 44724 43168 44736
rect 43123 44696 43168 44724
rect 43162 44684 43168 44696
rect 43220 44684 43226 44736
rect 45186 44724 45192 44736
rect 45147 44696 45192 44724
rect 45186 44684 45192 44696
rect 45244 44684 45250 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 7098 44520 7104 44532
rect 7059 44492 7104 44520
rect 7098 44480 7104 44492
rect 7156 44480 7162 44532
rect 9122 44520 9128 44532
rect 9083 44492 9128 44520
rect 9122 44480 9128 44492
rect 9180 44480 9186 44532
rect 9950 44480 9956 44532
rect 10008 44480 10014 44532
rect 11146 44520 11152 44532
rect 11107 44492 11152 44520
rect 11146 44480 11152 44492
rect 11204 44480 11210 44532
rect 45462 44520 45468 44532
rect 45423 44492 45468 44520
rect 45462 44480 45468 44492
rect 45520 44480 45526 44532
rect 6917 44455 6975 44461
rect 6917 44421 6929 44455
rect 6963 44452 6975 44455
rect 7006 44452 7012 44464
rect 6963 44424 7012 44452
rect 6963 44421 6975 44424
rect 6917 44415 6975 44421
rect 7006 44412 7012 44424
rect 7064 44412 7070 44464
rect 7282 44412 7288 44464
rect 7340 44452 7346 44464
rect 7929 44455 7987 44461
rect 7929 44452 7941 44455
rect 7340 44424 7941 44452
rect 7340 44412 7346 44424
rect 7929 44421 7941 44424
rect 7975 44452 7987 44455
rect 8757 44455 8815 44461
rect 8757 44452 8769 44455
rect 7975 44424 8769 44452
rect 7975 44421 7987 44424
rect 7929 44415 7987 44421
rect 8757 44421 8769 44424
rect 8803 44421 8815 44455
rect 9030 44452 9036 44464
rect 8991 44424 9036 44452
rect 8757 44415 8815 44421
rect 9030 44412 9036 44424
rect 9088 44412 9094 44464
rect 9968 44452 9996 44480
rect 9600 44424 9996 44452
rect 5813 44387 5871 44393
rect 5813 44353 5825 44387
rect 5859 44353 5871 44387
rect 5813 44347 5871 44353
rect 5828 44316 5856 44347
rect 5902 44344 5908 44396
rect 5960 44384 5966 44396
rect 7745 44387 7803 44393
rect 7745 44384 7757 44387
rect 5960 44356 7757 44384
rect 5960 44344 5966 44356
rect 7745 44353 7757 44356
rect 7791 44353 7803 44387
rect 7745 44347 7803 44353
rect 8941 44387 8999 44393
rect 8941 44353 8953 44387
rect 8987 44384 8999 44387
rect 9600 44384 9628 44424
rect 8987 44356 9628 44384
rect 8987 44353 8999 44356
rect 8941 44347 8999 44353
rect 9674 44344 9680 44396
rect 9732 44384 9738 44396
rect 10025 44387 10083 44393
rect 10025 44384 10037 44387
rect 9732 44356 10037 44384
rect 9732 44344 9738 44356
rect 10025 44353 10037 44356
rect 10071 44353 10083 44387
rect 36262 44384 36268 44396
rect 36223 44356 36268 44384
rect 10025 44347 10083 44353
rect 36262 44344 36268 44356
rect 36320 44344 36326 44396
rect 37734 44393 37740 44396
rect 37728 44384 37740 44393
rect 37695 44356 37740 44384
rect 37728 44347 37740 44356
rect 37734 44344 37740 44347
rect 37792 44344 37798 44396
rect 40037 44387 40095 44393
rect 40037 44353 40049 44387
rect 40083 44384 40095 44387
rect 40126 44384 40132 44396
rect 40083 44356 40132 44384
rect 40083 44353 40095 44356
rect 40037 44347 40095 44353
rect 40126 44344 40132 44356
rect 40184 44344 40190 44396
rect 40304 44387 40362 44393
rect 40304 44353 40316 44387
rect 40350 44384 40362 44387
rect 41877 44387 41935 44393
rect 41877 44384 41889 44387
rect 40350 44356 41889 44384
rect 40350 44353 40362 44356
rect 40304 44347 40362 44353
rect 41877 44353 41889 44356
rect 41923 44353 41935 44387
rect 44542 44384 44548 44396
rect 44503 44356 44548 44384
rect 41877 44347 41935 44353
rect 44542 44344 44548 44356
rect 44600 44344 44606 44396
rect 6822 44316 6828 44328
rect 5828 44288 6828 44316
rect 6822 44276 6828 44288
rect 6880 44276 6886 44328
rect 9766 44316 9772 44328
rect 9727 44288 9772 44316
rect 9766 44276 9772 44288
rect 9824 44276 9830 44328
rect 37274 44276 37280 44328
rect 37332 44316 37338 44328
rect 37461 44319 37519 44325
rect 37461 44316 37473 44319
rect 37332 44288 37473 44316
rect 37332 44276 37338 44288
rect 37461 44285 37473 44288
rect 37507 44285 37519 44319
rect 37461 44279 37519 44285
rect 44174 44276 44180 44328
rect 44232 44316 44238 44328
rect 45005 44319 45063 44325
rect 45005 44316 45017 44319
rect 44232 44288 45017 44316
rect 44232 44276 44238 44288
rect 45005 44285 45017 44288
rect 45051 44285 45063 44319
rect 45005 44279 45063 44285
rect 5626 44248 5632 44260
rect 5539 44220 5632 44248
rect 5626 44208 5632 44220
rect 5684 44248 5690 44260
rect 6549 44251 6607 44257
rect 6549 44248 6561 44251
rect 5684 44220 6561 44248
rect 5684 44208 5690 44220
rect 6549 44217 6561 44220
rect 6595 44217 6607 44251
rect 7561 44251 7619 44257
rect 7561 44248 7573 44251
rect 6549 44211 6607 44217
rect 6932 44220 7573 44248
rect 6932 44189 6960 44220
rect 7561 44217 7573 44220
rect 7607 44217 7619 44251
rect 7561 44211 7619 44217
rect 9309 44251 9367 44257
rect 9309 44217 9321 44251
rect 9355 44217 9367 44251
rect 9309 44211 9367 44217
rect 6917 44183 6975 44189
rect 6917 44149 6929 44183
rect 6963 44149 6975 44183
rect 9324 44180 9352 44211
rect 41046 44208 41052 44260
rect 41104 44248 41110 44260
rect 41104 44220 43300 44248
rect 41104 44208 41110 44220
rect 43272 44192 43300 44220
rect 44358 44208 44364 44260
rect 44416 44248 44422 44260
rect 45281 44251 45339 44257
rect 45281 44248 45293 44251
rect 44416 44220 45293 44248
rect 44416 44208 44422 44220
rect 45281 44217 45293 44220
rect 45327 44248 45339 44251
rect 45370 44248 45376 44260
rect 45327 44220 45376 44248
rect 45327 44217 45339 44220
rect 45281 44211 45339 44217
rect 45370 44208 45376 44220
rect 45428 44208 45434 44260
rect 10042 44180 10048 44192
rect 9324 44152 10048 44180
rect 6917 44143 6975 44149
rect 10042 44140 10048 44152
rect 10100 44180 10106 44192
rect 10502 44180 10508 44192
rect 10100 44152 10508 44180
rect 10100 44140 10106 44152
rect 10502 44140 10508 44152
rect 10560 44140 10566 44192
rect 24581 44183 24639 44189
rect 24581 44149 24593 44183
rect 24627 44180 24639 44183
rect 24854 44180 24860 44192
rect 24627 44152 24860 44180
rect 24627 44149 24639 44152
rect 24581 44143 24639 44149
rect 24854 44140 24860 44152
rect 24912 44140 24918 44192
rect 36909 44183 36967 44189
rect 36909 44149 36921 44183
rect 36955 44180 36967 44183
rect 37734 44180 37740 44192
rect 36955 44152 37740 44180
rect 36955 44149 36967 44152
rect 36909 44143 36967 44149
rect 37734 44140 37740 44152
rect 37792 44140 37798 44192
rect 38746 44140 38752 44192
rect 38804 44180 38810 44192
rect 38841 44183 38899 44189
rect 38841 44180 38853 44183
rect 38804 44152 38853 44180
rect 38804 44140 38810 44152
rect 38841 44149 38853 44152
rect 38887 44149 38899 44183
rect 38841 44143 38899 44149
rect 39577 44183 39635 44189
rect 39577 44149 39589 44183
rect 39623 44180 39635 44183
rect 40310 44180 40316 44192
rect 39623 44152 40316 44180
rect 39623 44149 39635 44152
rect 39577 44143 39635 44149
rect 40310 44140 40316 44152
rect 40368 44140 40374 44192
rect 41417 44183 41475 44189
rect 41417 44149 41429 44183
rect 41463 44180 41475 44183
rect 41966 44180 41972 44192
rect 41463 44152 41972 44180
rect 41463 44149 41475 44152
rect 41417 44143 41475 44149
rect 41966 44140 41972 44152
rect 42024 44140 42030 44192
rect 43254 44180 43260 44192
rect 43215 44152 43260 44180
rect 43254 44140 43260 44152
rect 43312 44140 43318 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 5902 43936 5908 43988
rect 5960 43976 5966 43988
rect 6457 43979 6515 43985
rect 6457 43976 6469 43979
rect 5960 43948 6469 43976
rect 5960 43936 5966 43948
rect 6457 43945 6469 43948
rect 6503 43945 6515 43979
rect 6457 43939 6515 43945
rect 9401 43979 9459 43985
rect 9401 43945 9413 43979
rect 9447 43976 9459 43979
rect 9674 43976 9680 43988
rect 9447 43948 9680 43976
rect 9447 43945 9459 43948
rect 9401 43939 9459 43945
rect 9674 43936 9680 43948
rect 9732 43936 9738 43988
rect 38470 43976 38476 43988
rect 38431 43948 38476 43976
rect 38470 43936 38476 43948
rect 38528 43936 38534 43988
rect 41506 43936 41512 43988
rect 41564 43976 41570 43988
rect 41877 43979 41935 43985
rect 41877 43976 41889 43979
rect 41564 43948 41889 43976
rect 41564 43936 41570 43948
rect 41877 43945 41889 43948
rect 41923 43945 41935 43979
rect 41877 43939 41935 43945
rect 43990 43936 43996 43988
rect 44048 43976 44054 43988
rect 44637 43979 44695 43985
rect 44637 43976 44649 43979
rect 44048 43948 44649 43976
rect 44048 43936 44054 43948
rect 44637 43945 44649 43948
rect 44683 43945 44695 43979
rect 45370 43976 45376 43988
rect 45331 43948 45376 43976
rect 44637 43939 44695 43945
rect 45370 43936 45376 43948
rect 45428 43936 45434 43988
rect 45554 43936 45560 43988
rect 45612 43976 45618 43988
rect 45612 43948 45657 43976
rect 45612 43936 45618 43948
rect 9125 43843 9183 43849
rect 9125 43809 9137 43843
rect 9171 43840 9183 43843
rect 9858 43840 9864 43852
rect 9171 43812 9864 43840
rect 9171 43809 9183 43812
rect 9125 43803 9183 43809
rect 9858 43800 9864 43812
rect 9916 43800 9922 43852
rect 38654 43840 38660 43852
rect 38615 43812 38660 43840
rect 38654 43800 38660 43812
rect 38712 43800 38718 43852
rect 41966 43840 41972 43852
rect 41927 43812 41972 43840
rect 41966 43800 41972 43812
rect 42024 43800 42030 43852
rect 9309 43775 9367 43781
rect 9309 43741 9321 43775
rect 9355 43741 9367 43775
rect 9309 43735 9367 43741
rect 9401 43775 9459 43781
rect 9401 43741 9413 43775
rect 9447 43741 9459 43775
rect 9401 43735 9459 43741
rect 6270 43704 6276 43716
rect 6231 43676 6276 43704
rect 6270 43664 6276 43676
rect 6328 43664 6334 43716
rect 6489 43707 6547 43713
rect 6489 43673 6501 43707
rect 6535 43704 6547 43707
rect 6822 43704 6828 43716
rect 6535 43676 6828 43704
rect 6535 43673 6547 43676
rect 6489 43667 6547 43673
rect 6822 43664 6828 43676
rect 6880 43664 6886 43716
rect 9122 43664 9128 43716
rect 9180 43704 9186 43716
rect 9324 43704 9352 43735
rect 9180 43676 9352 43704
rect 9416 43704 9444 43735
rect 9766 43732 9772 43784
rect 9824 43772 9830 43784
rect 11241 43775 11299 43781
rect 11241 43772 11253 43775
rect 9824 43744 11253 43772
rect 9824 43732 9830 43744
rect 11241 43741 11253 43744
rect 11287 43772 11299 43775
rect 12069 43775 12127 43781
rect 12069 43772 12081 43775
rect 11287 43744 12081 43772
rect 11287 43741 11299 43744
rect 11241 43735 11299 43741
rect 12069 43741 12081 43744
rect 12115 43741 12127 43775
rect 24578 43772 24584 43784
rect 24539 43744 24584 43772
rect 12069 43735 12127 43741
rect 24578 43732 24584 43744
rect 24636 43732 24642 43784
rect 24854 43781 24860 43784
rect 24848 43772 24860 43781
rect 24815 43744 24860 43772
rect 24848 43735 24860 43744
rect 24854 43732 24860 43735
rect 24912 43732 24918 43784
rect 36173 43775 36231 43781
rect 36173 43741 36185 43775
rect 36219 43741 36231 43775
rect 36173 43735 36231 43741
rect 36633 43775 36691 43781
rect 36633 43741 36645 43775
rect 36679 43772 36691 43775
rect 37274 43772 37280 43784
rect 36679 43744 37280 43772
rect 36679 43741 36691 43744
rect 36633 43735 36691 43741
rect 10778 43704 10784 43716
rect 9416 43676 10784 43704
rect 9180 43664 9186 43676
rect 10778 43664 10784 43676
rect 10836 43664 10842 43716
rect 10962 43704 10968 43716
rect 11020 43713 11026 43716
rect 12342 43713 12348 43716
rect 10932 43676 10968 43704
rect 10962 43664 10968 43676
rect 11020 43667 11032 43713
rect 12336 43667 12348 43713
rect 12400 43704 12406 43716
rect 36188 43704 36216 43735
rect 37274 43732 37280 43744
rect 37332 43732 37338 43784
rect 38746 43772 38752 43784
rect 38707 43744 38752 43772
rect 38746 43732 38752 43744
rect 38804 43732 38810 43784
rect 40037 43775 40095 43781
rect 40037 43741 40049 43775
rect 40083 43772 40095 43775
rect 40126 43772 40132 43784
rect 40083 43744 40132 43772
rect 40083 43741 40095 43744
rect 40037 43735 40095 43741
rect 40126 43732 40132 43744
rect 40184 43732 40190 43784
rect 40310 43781 40316 43784
rect 40304 43772 40316 43781
rect 40271 43744 40316 43772
rect 40304 43735 40316 43744
rect 40310 43732 40316 43735
rect 40368 43732 40374 43784
rect 42150 43772 42156 43784
rect 42111 43744 42156 43772
rect 42150 43732 42156 43744
rect 42208 43732 42214 43784
rect 43254 43772 43260 43784
rect 43167 43744 43260 43772
rect 43254 43732 43260 43744
rect 43312 43772 43318 43784
rect 44266 43772 44272 43784
rect 43312 43744 44272 43772
rect 43312 43732 43318 43744
rect 44266 43732 44272 43744
rect 44324 43772 44330 43784
rect 45002 43772 45008 43784
rect 44324 43744 45008 43772
rect 44324 43732 44330 43744
rect 45002 43732 45008 43744
rect 45060 43732 45066 43784
rect 36878 43707 36936 43713
rect 36878 43704 36890 43707
rect 12400 43676 12436 43704
rect 36188 43676 36890 43704
rect 11020 43664 11026 43667
rect 12342 43664 12348 43667
rect 12400 43664 12406 43676
rect 36878 43673 36890 43676
rect 36924 43673 36936 43707
rect 36878 43667 36936 43673
rect 38473 43707 38531 43713
rect 38473 43673 38485 43707
rect 38519 43673 38531 43707
rect 38473 43667 38531 43673
rect 41877 43707 41935 43713
rect 41877 43673 41889 43707
rect 41923 43673 41935 43707
rect 41877 43667 41935 43673
rect 6641 43639 6699 43645
rect 6641 43605 6653 43639
rect 6687 43636 6699 43639
rect 7098 43636 7104 43648
rect 6687 43608 7104 43636
rect 6687 43605 6699 43608
rect 6641 43599 6699 43605
rect 7098 43596 7104 43608
rect 7156 43596 7162 43648
rect 9858 43636 9864 43648
rect 9819 43608 9864 43636
rect 9858 43596 9864 43608
rect 9916 43596 9922 43648
rect 13262 43596 13268 43648
rect 13320 43636 13326 43648
rect 13449 43639 13507 43645
rect 13449 43636 13461 43639
rect 13320 43608 13461 43636
rect 13320 43596 13326 43608
rect 13449 43605 13461 43608
rect 13495 43605 13507 43639
rect 13449 43599 13507 43605
rect 25498 43596 25504 43648
rect 25556 43636 25562 43648
rect 25961 43639 26019 43645
rect 25961 43636 25973 43639
rect 25556 43608 25973 43636
rect 25556 43596 25562 43608
rect 25961 43605 25973 43608
rect 26007 43605 26019 43639
rect 25961 43599 26019 43605
rect 38013 43639 38071 43645
rect 38013 43605 38025 43639
rect 38059 43636 38071 43639
rect 38488 43636 38516 43667
rect 38059 43608 38516 43636
rect 38933 43639 38991 43645
rect 38059 43605 38071 43608
rect 38013 43599 38071 43605
rect 38933 43605 38945 43639
rect 38979 43636 38991 43639
rect 40954 43636 40960 43648
rect 38979 43608 40960 43636
rect 38979 43605 38991 43608
rect 38933 43599 38991 43605
rect 40954 43596 40960 43608
rect 41012 43596 41018 43648
rect 41417 43639 41475 43645
rect 41417 43605 41429 43639
rect 41463 43636 41475 43639
rect 41892 43636 41920 43667
rect 43162 43664 43168 43716
rect 43220 43704 43226 43716
rect 43502 43707 43560 43713
rect 43502 43704 43514 43707
rect 43220 43676 43514 43704
rect 43220 43664 43226 43676
rect 43502 43673 43514 43676
rect 43548 43673 43560 43707
rect 43502 43667 43560 43673
rect 43622 43664 43628 43716
rect 43680 43704 43686 43716
rect 45189 43707 45247 43713
rect 45189 43704 45201 43707
rect 43680 43676 45201 43704
rect 43680 43664 43686 43676
rect 45189 43673 45201 43676
rect 45235 43673 45247 43707
rect 45189 43667 45247 43673
rect 42334 43636 42340 43648
rect 41463 43608 41920 43636
rect 42295 43608 42340 43636
rect 41463 43605 41475 43608
rect 41417 43599 41475 43605
rect 42334 43596 42340 43608
rect 42392 43596 42398 43648
rect 44818 43596 44824 43648
rect 44876 43636 44882 43648
rect 45389 43639 45447 43645
rect 45389 43636 45401 43639
rect 44876 43608 45401 43636
rect 44876 43596 44882 43608
rect 45389 43605 45401 43608
rect 45435 43605 45447 43639
rect 45389 43599 45447 43605
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 10962 43392 10968 43444
rect 11020 43432 11026 43444
rect 11057 43435 11115 43441
rect 11057 43432 11069 43435
rect 11020 43404 11069 43432
rect 11020 43392 11026 43404
rect 11057 43401 11069 43404
rect 11103 43401 11115 43435
rect 11057 43395 11115 43401
rect 38654 43392 38660 43444
rect 38712 43432 38718 43444
rect 38841 43435 38899 43441
rect 38841 43432 38853 43435
rect 38712 43404 38853 43432
rect 38712 43392 38718 43404
rect 38841 43401 38853 43404
rect 38887 43401 38899 43435
rect 38841 43395 38899 43401
rect 43257 43435 43315 43441
rect 43257 43401 43269 43435
rect 43303 43432 43315 43435
rect 43622 43432 43628 43444
rect 43303 43404 43628 43432
rect 43303 43401 43315 43404
rect 43257 43395 43315 43401
rect 43622 43392 43628 43404
rect 43680 43392 43686 43444
rect 43717 43435 43775 43441
rect 43717 43401 43729 43435
rect 43763 43432 43775 43435
rect 44174 43432 44180 43444
rect 43763 43404 44180 43432
rect 43763 43401 43775 43404
rect 43717 43395 43775 43401
rect 5626 43364 5632 43376
rect 5587 43336 5632 43364
rect 5626 43324 5632 43336
rect 5684 43324 5690 43376
rect 6733 43367 6791 43373
rect 6733 43333 6745 43367
rect 6779 43364 6791 43367
rect 7006 43364 7012 43376
rect 6779 43336 7012 43364
rect 6779 43333 6791 43336
rect 6733 43327 6791 43333
rect 7006 43324 7012 43336
rect 7064 43364 7070 43376
rect 7650 43364 7656 43376
rect 7064 43336 7656 43364
rect 7064 43324 7070 43336
rect 7650 43324 7656 43336
rect 7708 43324 7714 43376
rect 9122 43324 9128 43376
rect 9180 43364 9186 43376
rect 37734 43373 37740 43376
rect 37728 43364 37740 43373
rect 9180 43336 11192 43364
rect 37695 43336 37740 43364
rect 9180 43324 9186 43336
rect 5813 43299 5871 43305
rect 5813 43265 5825 43299
rect 5859 43296 5871 43299
rect 6270 43296 6276 43308
rect 5859 43268 6276 43296
rect 5859 43265 5871 43268
rect 5813 43259 5871 43265
rect 6270 43256 6276 43268
rect 6328 43256 6334 43308
rect 7098 43296 7104 43308
rect 7059 43268 7104 43296
rect 7098 43256 7104 43268
rect 7156 43256 7162 43308
rect 8754 43296 8760 43308
rect 8715 43268 8760 43296
rect 8754 43256 8760 43268
rect 8812 43256 8818 43308
rect 10962 43296 10968 43308
rect 10923 43268 10968 43296
rect 10962 43256 10968 43268
rect 11020 43256 11026 43308
rect 11164 43305 11192 43336
rect 37728 43327 37740 43336
rect 37734 43324 37740 43327
rect 37792 43324 37798 43376
rect 40954 43364 40960 43376
rect 40915 43336 40960 43364
rect 40954 43324 40960 43336
rect 41012 43324 41018 43376
rect 42334 43364 42340 43376
rect 41064 43336 42340 43364
rect 11149 43299 11207 43305
rect 11149 43265 11161 43299
rect 11195 43265 11207 43299
rect 12342 43296 12348 43308
rect 12303 43268 12348 43296
rect 11149 43259 11207 43265
rect 12342 43256 12348 43268
rect 12400 43256 12406 43308
rect 41064 43305 41092 43336
rect 42334 43324 42340 43336
rect 42392 43324 42398 43376
rect 41049 43299 41107 43305
rect 41049 43265 41061 43299
rect 41095 43265 41107 43299
rect 41322 43296 41328 43308
rect 41283 43268 41328 43296
rect 41049 43259 41107 43265
rect 41322 43256 41328 43268
rect 41380 43256 41386 43308
rect 43073 43299 43131 43305
rect 43073 43265 43085 43299
rect 43119 43265 43131 43299
rect 43073 43259 43131 43265
rect 43257 43299 43315 43305
rect 43257 43265 43269 43299
rect 43303 43296 43315 43299
rect 43732 43296 43760 43395
rect 44174 43392 44180 43404
rect 44232 43392 44238 43444
rect 44852 43367 44910 43373
rect 44852 43333 44864 43367
rect 44898 43364 44910 43367
rect 45186 43364 45192 43376
rect 44898 43336 45192 43364
rect 44898 43333 44910 43336
rect 44852 43327 44910 43333
rect 45186 43324 45192 43336
rect 45244 43324 45250 43376
rect 43303 43268 43760 43296
rect 43303 43265 43315 43268
rect 43257 43259 43315 43265
rect 37274 43188 37280 43240
rect 37332 43228 37338 43240
rect 37461 43231 37519 43237
rect 37461 43228 37473 43231
rect 37332 43200 37473 43228
rect 37332 43188 37338 43200
rect 37461 43197 37473 43200
rect 37507 43197 37519 43231
rect 43088 43228 43116 43259
rect 45002 43256 45008 43308
rect 45060 43296 45066 43308
rect 45097 43299 45155 43305
rect 45097 43296 45109 43299
rect 45060 43268 45109 43296
rect 45060 43256 45066 43268
rect 45097 43265 45109 43268
rect 45143 43265 45155 43299
rect 45097 43259 45155 43265
rect 43990 43228 43996 43240
rect 43088 43200 43996 43228
rect 37461 43191 37519 43197
rect 43990 43188 43996 43200
rect 44048 43188 44054 43240
rect 5997 43163 6055 43169
rect 5997 43129 6009 43163
rect 6043 43160 6055 43163
rect 41141 43163 41199 43169
rect 6043 43132 6776 43160
rect 6043 43129 6055 43132
rect 5997 43123 6055 43129
rect 5902 43052 5908 43104
rect 5960 43092 5966 43104
rect 6748 43101 6776 43132
rect 41141 43129 41153 43163
rect 41187 43160 41199 43163
rect 42610 43160 42616 43172
rect 41187 43132 42616 43160
rect 41187 43129 41199 43132
rect 41141 43123 41199 43129
rect 42610 43120 42616 43132
rect 42668 43120 42674 43172
rect 6549 43095 6607 43101
rect 6549 43092 6561 43095
rect 5960 43064 6561 43092
rect 5960 43052 5966 43064
rect 6549 43061 6561 43064
rect 6595 43061 6607 43095
rect 6549 43055 6607 43061
rect 6733 43095 6791 43101
rect 6733 43061 6745 43095
rect 6779 43061 6791 43095
rect 6733 43055 6791 43061
rect 9766 43052 9772 43104
rect 9824 43092 9830 43104
rect 10045 43095 10103 43101
rect 10045 43092 10057 43095
rect 9824 43064 10057 43092
rect 9824 43052 9830 43064
rect 10045 43061 10057 43064
rect 10091 43061 10103 43095
rect 10045 43055 10103 43061
rect 41325 43095 41383 43101
rect 41325 43061 41337 43095
rect 41371 43092 41383 43095
rect 44358 43092 44364 43104
rect 41371 43064 44364 43092
rect 41371 43061 41383 43064
rect 41325 43055 41383 43061
rect 44358 43052 44364 43064
rect 44416 43052 44422 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 6270 42848 6276 42900
rect 6328 42888 6334 42900
rect 6365 42891 6423 42897
rect 6365 42888 6377 42891
rect 6328 42860 6377 42888
rect 6328 42848 6334 42860
rect 6365 42857 6377 42860
rect 6411 42857 6423 42891
rect 6365 42851 6423 42857
rect 6730 42848 6736 42900
rect 6788 42888 6794 42900
rect 6825 42891 6883 42897
rect 6825 42888 6837 42891
rect 6788 42860 6837 42888
rect 6788 42848 6794 42860
rect 6825 42857 6837 42860
rect 6871 42888 6883 42891
rect 9122 42888 9128 42900
rect 6871 42860 9128 42888
rect 6871 42857 6883 42860
rect 6825 42851 6883 42857
rect 9122 42848 9128 42860
rect 9180 42848 9186 42900
rect 44453 42891 44511 42897
rect 44453 42857 44465 42891
rect 44499 42888 44511 42891
rect 44818 42888 44824 42900
rect 44499 42860 44824 42888
rect 44499 42857 44511 42860
rect 44453 42851 44511 42857
rect 44818 42848 44824 42860
rect 44876 42848 44882 42900
rect 7650 42780 7656 42832
rect 7708 42820 7714 42832
rect 7929 42823 7987 42829
rect 7929 42820 7941 42823
rect 7708 42792 7941 42820
rect 7708 42780 7714 42792
rect 7929 42789 7941 42792
rect 7975 42789 7987 42823
rect 7929 42783 7987 42789
rect 9125 42755 9183 42761
rect 9125 42752 9137 42755
rect 6932 42724 9137 42752
rect 6932 42696 6960 42724
rect 9125 42721 9137 42724
rect 9171 42721 9183 42755
rect 9125 42715 9183 42721
rect 4985 42687 5043 42693
rect 4985 42653 4997 42687
rect 5031 42684 5043 42687
rect 6914 42684 6920 42696
rect 5031 42656 6920 42684
rect 5031 42653 5043 42656
rect 4985 42647 5043 42653
rect 6914 42644 6920 42656
rect 6972 42644 6978 42696
rect 7012 42665 7070 42671
rect 7012 42631 7024 42665
rect 7058 42631 7070 42665
rect 7098 42644 7104 42696
rect 7156 42684 7162 42696
rect 7282 42684 7288 42696
rect 7156 42656 7201 42684
rect 7243 42656 7288 42684
rect 7156 42644 7162 42656
rect 7282 42644 7288 42656
rect 7340 42644 7346 42696
rect 7377 42687 7435 42693
rect 7377 42653 7389 42687
rect 7423 42653 7435 42687
rect 9140 42684 9168 42715
rect 9766 42684 9772 42696
rect 9140 42656 9772 42684
rect 7377 42647 7435 42653
rect 7012 42628 7070 42631
rect 5252 42619 5310 42625
rect 5252 42585 5264 42619
rect 5298 42616 5310 42619
rect 5718 42616 5724 42628
rect 5298 42588 5724 42616
rect 5298 42585 5310 42588
rect 5252 42579 5310 42585
rect 5718 42576 5724 42588
rect 5776 42576 5782 42628
rect 7006 42576 7012 42628
rect 7064 42576 7070 42628
rect 7392 42616 7420 42647
rect 9766 42644 9772 42656
rect 9824 42644 9830 42696
rect 24210 42644 24216 42696
rect 24268 42684 24274 42696
rect 24581 42687 24639 42693
rect 24581 42684 24593 42687
rect 24268 42656 24593 42684
rect 24268 42644 24274 42656
rect 24581 42653 24593 42656
rect 24627 42653 24639 42687
rect 33870 42684 33876 42696
rect 33831 42656 33876 42684
rect 24581 42647 24639 42653
rect 33870 42644 33876 42656
rect 33928 42644 33934 42696
rect 35066 42684 35072 42696
rect 35027 42656 35072 42684
rect 35066 42644 35072 42656
rect 35124 42644 35130 42696
rect 37366 42644 37372 42696
rect 37424 42684 37430 42696
rect 37461 42687 37519 42693
rect 37461 42684 37473 42687
rect 37424 42656 37473 42684
rect 37424 42644 37430 42656
rect 37461 42653 37473 42656
rect 37507 42653 37519 42687
rect 37461 42647 37519 42653
rect 43990 42644 43996 42696
rect 44048 42684 44054 42696
rect 44085 42687 44143 42693
rect 44085 42684 44097 42687
rect 44048 42656 44097 42684
rect 44048 42644 44054 42656
rect 44085 42653 44097 42656
rect 44131 42653 44143 42687
rect 44085 42647 44143 42653
rect 44174 42644 44180 42696
rect 44232 42684 44238 42696
rect 44269 42687 44327 42693
rect 44269 42684 44281 42687
rect 44232 42656 44281 42684
rect 44232 42644 44238 42656
rect 44269 42653 44281 42656
rect 44315 42684 44327 42687
rect 44358 42684 44364 42696
rect 44315 42656 44364 42684
rect 44315 42653 44327 42656
rect 44269 42647 44327 42653
rect 44358 42644 44364 42656
rect 44416 42644 44422 42696
rect 8294 42616 8300 42628
rect 7208 42588 7420 42616
rect 8255 42588 8300 42616
rect 7208 42560 7236 42588
rect 8294 42576 8300 42588
rect 8352 42576 8358 42628
rect 9030 42576 9036 42628
rect 9088 42616 9094 42628
rect 9370 42619 9428 42625
rect 9370 42616 9382 42619
rect 9088 42588 9382 42616
rect 9088 42576 9094 42588
rect 9370 42585 9382 42588
rect 9416 42585 9428 42619
rect 9370 42579 9428 42585
rect 7190 42508 7196 42560
rect 7248 42508 7254 42560
rect 7374 42508 7380 42560
rect 7432 42548 7438 42560
rect 7837 42551 7895 42557
rect 7837 42548 7849 42551
rect 7432 42520 7849 42548
rect 7432 42508 7438 42520
rect 7837 42517 7849 42520
rect 7883 42517 7895 42551
rect 10502 42548 10508 42560
rect 10463 42520 10508 42548
rect 7837 42511 7895 42517
rect 10502 42508 10508 42520
rect 10560 42508 10566 42560
rect 38102 42548 38108 42560
rect 38063 42520 38108 42548
rect 38102 42508 38108 42520
rect 38160 42508 38166 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 5718 42344 5724 42356
rect 5679 42316 5724 42344
rect 5718 42304 5724 42316
rect 5776 42304 5782 42356
rect 9030 42344 9036 42356
rect 8991 42316 9036 42344
rect 9030 42304 9036 42316
rect 9088 42304 9094 42356
rect 10137 42347 10195 42353
rect 10137 42313 10149 42347
rect 10183 42344 10195 42347
rect 10962 42344 10968 42356
rect 10183 42316 10968 42344
rect 10183 42313 10195 42316
rect 10137 42307 10195 42313
rect 10962 42304 10968 42316
rect 11020 42304 11026 42356
rect 10502 42276 10508 42288
rect 8956 42248 10508 42276
rect 5902 42208 5908 42220
rect 5863 42180 5908 42208
rect 5902 42168 5908 42180
rect 5960 42168 5966 42220
rect 6730 42208 6736 42220
rect 6691 42180 6736 42208
rect 6730 42168 6736 42180
rect 6788 42168 6794 42220
rect 7006 42208 7012 42220
rect 6967 42180 7012 42208
rect 7006 42168 7012 42180
rect 7064 42168 7070 42220
rect 7098 42168 7104 42220
rect 7156 42208 7162 42220
rect 7193 42211 7251 42217
rect 7193 42208 7205 42211
rect 7156 42180 7205 42208
rect 7156 42168 7162 42180
rect 7193 42177 7205 42180
rect 7239 42208 7251 42211
rect 8294 42208 8300 42220
rect 7239 42180 8300 42208
rect 7239 42177 7251 42180
rect 7193 42171 7251 42177
rect 8294 42168 8300 42180
rect 8352 42168 8358 42220
rect 8956 42217 8984 42248
rect 8941 42211 8999 42217
rect 8941 42177 8953 42211
rect 8987 42177 8999 42211
rect 9122 42208 9128 42220
rect 9083 42180 9128 42208
rect 8941 42171 8999 42177
rect 9122 42168 9128 42180
rect 9180 42168 9186 42220
rect 9784 42217 9812 42248
rect 10502 42236 10508 42248
rect 10560 42236 10566 42288
rect 24210 42285 24216 42288
rect 24204 42276 24216 42285
rect 22020 42248 23428 42276
rect 24171 42248 24216 42276
rect 22020 42217 22048 42248
rect 9769 42211 9827 42217
rect 9769 42177 9781 42211
rect 9815 42177 9827 42211
rect 9769 42171 9827 42177
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22261 42211 22319 42217
rect 22261 42208 22273 42211
rect 22005 42171 22063 42177
rect 22112 42180 22273 42208
rect 9858 42140 9864 42152
rect 9819 42112 9864 42140
rect 9858 42100 9864 42112
rect 9916 42100 9922 42152
rect 21453 42143 21511 42149
rect 21453 42109 21465 42143
rect 21499 42140 21511 42143
rect 22112 42140 22140 42180
rect 22261 42177 22273 42180
rect 22307 42177 22319 42211
rect 22261 42171 22319 42177
rect 23400 42152 23428 42248
rect 24204 42239 24216 42248
rect 24210 42236 24216 42239
rect 24268 42236 24274 42288
rect 28813 42279 28871 42285
rect 28813 42245 28825 42279
rect 28859 42276 28871 42279
rect 31113 42279 31171 42285
rect 31113 42276 31125 42279
rect 28859 42248 31125 42276
rect 28859 42245 28871 42248
rect 28813 42239 28871 42245
rect 31113 42245 31125 42248
rect 31159 42276 31171 42279
rect 32398 42276 32404 42288
rect 31159 42248 32404 42276
rect 31159 42245 31171 42248
rect 31113 42239 31171 42245
rect 24762 42168 24768 42220
rect 24820 42208 24826 42220
rect 28828 42208 28856 42239
rect 32398 42236 32404 42248
rect 32456 42276 32462 42288
rect 37461 42279 37519 42285
rect 37461 42276 37473 42279
rect 32456 42248 37473 42276
rect 32456 42236 32462 42248
rect 37461 42245 37473 42248
rect 37507 42276 37519 42279
rect 38102 42276 38108 42288
rect 37507 42248 38108 42276
rect 37507 42245 37519 42248
rect 37461 42239 37519 42245
rect 38102 42236 38108 42248
rect 38160 42276 38166 42288
rect 39206 42276 39212 42288
rect 38160 42248 39212 42276
rect 38160 42236 38166 42248
rect 39206 42236 39212 42248
rect 39264 42236 39270 42288
rect 44174 42236 44180 42288
rect 44232 42276 44238 42288
rect 44232 42248 44680 42276
rect 44232 42236 44238 42248
rect 33870 42217 33876 42220
rect 33864 42208 33876 42217
rect 24820 42180 28856 42208
rect 33831 42180 33876 42208
rect 24820 42168 24826 42180
rect 33864 42171 33876 42180
rect 33870 42168 33876 42171
rect 33928 42168 33934 42220
rect 35066 42168 35072 42220
rect 35124 42208 35130 42220
rect 36550 42211 36608 42217
rect 36550 42208 36562 42211
rect 35124 42180 36562 42208
rect 35124 42168 35130 42180
rect 36550 42177 36562 42180
rect 36596 42177 36608 42211
rect 36550 42171 36608 42177
rect 43990 42168 43996 42220
rect 44048 42208 44054 42220
rect 44269 42211 44327 42217
rect 44269 42208 44281 42211
rect 44048 42180 44281 42208
rect 44048 42168 44054 42180
rect 44269 42177 44281 42180
rect 44315 42177 44327 42211
rect 44269 42171 44327 42177
rect 44358 42168 44364 42220
rect 44416 42208 44422 42220
rect 44652 42217 44680 42248
rect 44545 42211 44603 42217
rect 44416 42180 44461 42208
rect 44416 42168 44422 42180
rect 44545 42177 44557 42211
rect 44591 42177 44603 42211
rect 44545 42171 44603 42177
rect 44637 42211 44695 42217
rect 44637 42177 44649 42211
rect 44683 42177 44695 42211
rect 44637 42171 44695 42177
rect 21499 42112 22140 42140
rect 21499 42109 21511 42112
rect 21453 42103 21511 42109
rect 23382 42100 23388 42152
rect 23440 42140 23446 42152
rect 23937 42143 23995 42149
rect 23937 42140 23949 42143
rect 23440 42112 23949 42140
rect 23440 42100 23446 42112
rect 23937 42109 23949 42112
rect 23983 42109 23995 42143
rect 23937 42103 23995 42109
rect 33318 42100 33324 42152
rect 33376 42140 33382 42152
rect 33597 42143 33655 42149
rect 33597 42140 33609 42143
rect 33376 42112 33609 42140
rect 33376 42100 33382 42112
rect 33597 42109 33609 42112
rect 33643 42109 33655 42143
rect 33597 42103 33655 42109
rect 36817 42143 36875 42149
rect 36817 42109 36829 42143
rect 36863 42140 36875 42143
rect 37274 42140 37280 42152
rect 36863 42112 37280 42140
rect 36863 42109 36875 42112
rect 36817 42103 36875 42109
rect 37274 42100 37280 42112
rect 37332 42140 37338 42152
rect 38562 42140 38568 42152
rect 37332 42112 38568 42140
rect 37332 42100 37338 42112
rect 38562 42100 38568 42112
rect 38620 42140 38626 42152
rect 38620 42112 38792 42140
rect 38620 42100 38626 42112
rect 28994 42032 29000 42084
rect 29052 42072 29058 42084
rect 38764 42081 38792 42112
rect 30101 42075 30159 42081
rect 30101 42072 30113 42075
rect 29052 42044 30113 42072
rect 29052 42032 29058 42044
rect 30101 42041 30113 42044
rect 30147 42041 30159 42075
rect 30101 42035 30159 42041
rect 38749 42075 38807 42081
rect 38749 42041 38761 42075
rect 38795 42041 38807 42075
rect 38749 42035 38807 42041
rect 39298 42032 39304 42084
rect 39356 42072 39362 42084
rect 44085 42075 44143 42081
rect 44085 42072 44097 42075
rect 39356 42044 44097 42072
rect 39356 42032 39362 42044
rect 44085 42041 44097 42044
rect 44131 42041 44143 42075
rect 44560 42072 44588 42171
rect 44634 42072 44640 42084
rect 44560 42044 44640 42072
rect 44085 42035 44143 42041
rect 44634 42032 44640 42044
rect 44692 42032 44698 42084
rect 5902 41964 5908 42016
rect 5960 42004 5966 42016
rect 6549 42007 6607 42013
rect 6549 42004 6561 42007
rect 5960 41976 6561 42004
rect 5960 41964 5966 41976
rect 6549 41973 6561 41976
rect 6595 41973 6607 42007
rect 12066 42004 12072 42016
rect 12027 41976 12072 42004
rect 6549 41967 6607 41973
rect 12066 41964 12072 41976
rect 12124 41964 12130 42016
rect 15286 42004 15292 42016
rect 15247 41976 15292 42004
rect 15286 41964 15292 41976
rect 15344 41964 15350 42016
rect 23014 41964 23020 42016
rect 23072 42004 23078 42016
rect 23385 42007 23443 42013
rect 23385 42004 23397 42007
rect 23072 41976 23397 42004
rect 23072 41964 23078 41976
rect 23385 41973 23397 41976
rect 23431 41973 23443 42007
rect 23385 41967 23443 41973
rect 25317 42007 25375 42013
rect 25317 41973 25329 42007
rect 25363 42004 25375 42007
rect 25590 42004 25596 42016
rect 25363 41976 25596 42004
rect 25363 41973 25375 41976
rect 25317 41967 25375 41973
rect 25590 41964 25596 41976
rect 25648 41964 25654 42016
rect 34790 41964 34796 42016
rect 34848 42004 34854 42016
rect 34977 42007 35035 42013
rect 34977 42004 34989 42007
rect 34848 41976 34989 42004
rect 34848 41964 34854 41976
rect 34977 41973 34989 41976
rect 35023 41973 35035 42007
rect 34977 41967 35035 41973
rect 35342 41964 35348 42016
rect 35400 42004 35406 42016
rect 35437 42007 35495 42013
rect 35437 42004 35449 42007
rect 35400 41976 35449 42004
rect 35400 41964 35406 41976
rect 35437 41973 35449 41976
rect 35483 41973 35495 42007
rect 40678 42004 40684 42016
rect 40639 41976 40684 42004
rect 35437 41967 35495 41973
rect 40678 41964 40684 41976
rect 40736 41964 40742 42016
rect 43438 42004 43444 42016
rect 43399 41976 43444 42004
rect 43438 41964 43444 41976
rect 43496 41964 43502 42016
rect 45094 42004 45100 42016
rect 45055 41976 45100 42004
rect 45094 41964 45100 41976
rect 45152 41964 45158 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 7009 41803 7067 41809
rect 7009 41769 7021 41803
rect 7055 41800 7067 41803
rect 7098 41800 7104 41812
rect 7055 41772 7104 41800
rect 7055 41769 7067 41772
rect 7009 41763 7067 41769
rect 7098 41760 7104 41772
rect 7156 41760 7162 41812
rect 7650 41800 7656 41812
rect 7611 41772 7656 41800
rect 7650 41760 7656 41772
rect 7708 41760 7714 41812
rect 13262 41800 13268 41812
rect 13223 41772 13268 41800
rect 13262 41760 13268 41772
rect 13320 41760 13326 41812
rect 27246 41800 27252 41812
rect 27207 41772 27252 41800
rect 27246 41760 27252 41772
rect 27304 41760 27310 41812
rect 35342 41800 35348 41812
rect 35303 41772 35348 41800
rect 35342 41760 35348 41772
rect 35400 41760 35406 41812
rect 35529 41803 35587 41809
rect 35529 41769 35541 41803
rect 35575 41800 35587 41803
rect 39025 41803 39083 41809
rect 39025 41800 39037 41803
rect 35575 41772 39037 41800
rect 35575 41769 35587 41772
rect 35529 41763 35587 41769
rect 39025 41769 39037 41772
rect 39071 41769 39083 41803
rect 39025 41763 39083 41769
rect 39485 41803 39543 41809
rect 39485 41769 39497 41803
rect 39531 41800 39543 41803
rect 41322 41800 41328 41812
rect 39531 41772 41328 41800
rect 39531 41769 39543 41772
rect 39485 41763 39543 41769
rect 41322 41760 41328 41772
rect 41380 41760 41386 41812
rect 44634 41800 44640 41812
rect 44595 41772 44640 41800
rect 44634 41760 44640 41772
rect 44692 41760 44698 41812
rect 34333 41735 34391 41741
rect 34333 41701 34345 41735
rect 34379 41701 34391 41735
rect 34333 41695 34391 41701
rect 7282 41624 7288 41676
rect 7340 41664 7346 41676
rect 7340 41636 7696 41664
rect 7340 41624 7346 41636
rect 5258 41556 5264 41608
rect 5316 41596 5322 41608
rect 5902 41605 5908 41608
rect 5629 41599 5687 41605
rect 5629 41596 5641 41599
rect 5316 41568 5641 41596
rect 5316 41556 5322 41568
rect 5629 41565 5641 41568
rect 5675 41565 5687 41599
rect 5896 41596 5908 41605
rect 5863 41568 5908 41596
rect 5629 41559 5687 41565
rect 5896 41559 5908 41568
rect 5902 41556 5908 41559
rect 5960 41556 5966 41608
rect 7190 41556 7196 41608
rect 7248 41596 7254 41608
rect 7668 41605 7696 41636
rect 9122 41624 9128 41676
rect 9180 41664 9186 41676
rect 9766 41664 9772 41676
rect 9180 41636 9772 41664
rect 9180 41624 9186 41636
rect 9766 41624 9772 41636
rect 9824 41664 9830 41676
rect 11149 41667 11207 41673
rect 11149 41664 11161 41667
rect 9824 41636 11161 41664
rect 9824 41624 9830 41636
rect 11149 41633 11161 41636
rect 11195 41633 11207 41667
rect 24578 41664 24584 41676
rect 24539 41636 24584 41664
rect 11149 41627 11207 41633
rect 24578 41624 24584 41636
rect 24636 41624 24642 41676
rect 28994 41664 29000 41676
rect 26206 41636 29000 41664
rect 7469 41599 7527 41605
rect 7469 41596 7481 41599
rect 7248 41568 7481 41596
rect 7248 41556 7254 41568
rect 7469 41565 7481 41568
rect 7515 41565 7527 41599
rect 7469 41559 7527 41565
rect 7653 41599 7711 41605
rect 7653 41565 7665 41599
rect 7699 41565 7711 41599
rect 7653 41559 7711 41565
rect 9309 41599 9367 41605
rect 9309 41565 9321 41599
rect 9355 41596 9367 41599
rect 9398 41596 9404 41608
rect 9355 41568 9404 41596
rect 9355 41565 9367 41568
rect 9309 41559 9367 41565
rect 7668 41460 7696 41559
rect 9398 41556 9404 41568
rect 9456 41556 9462 41608
rect 13170 41596 13176 41608
rect 13131 41568 13176 41596
rect 13170 41556 13176 41568
rect 13228 41556 13234 41608
rect 13262 41556 13268 41608
rect 13320 41596 13326 41608
rect 14918 41596 14924 41608
rect 13320 41568 13365 41596
rect 14879 41568 14924 41596
rect 13320 41556 13326 41568
rect 14918 41556 14924 41568
rect 14976 41556 14982 41608
rect 15188 41599 15246 41605
rect 15188 41565 15200 41599
rect 15234 41596 15246 41599
rect 16761 41599 16819 41605
rect 16761 41596 16773 41599
rect 15234 41568 16773 41596
rect 15234 41565 15246 41568
rect 15188 41559 15246 41565
rect 16761 41565 16773 41568
rect 16807 41565 16819 41599
rect 16761 41559 16819 41565
rect 20717 41599 20775 41605
rect 20717 41565 20729 41599
rect 20763 41596 20775 41599
rect 22094 41596 22100 41608
rect 20763 41568 22100 41596
rect 20763 41565 20775 41568
rect 20717 41559 20775 41565
rect 22094 41556 22100 41568
rect 22152 41556 22158 41608
rect 24029 41599 24087 41605
rect 24029 41565 24041 41599
rect 24075 41565 24087 41599
rect 24596 41596 24624 41624
rect 25222 41596 25228 41608
rect 24596 41568 25228 41596
rect 24029 41559 24087 41565
rect 11146 41488 11152 41540
rect 11204 41528 11210 41540
rect 11394 41531 11452 41537
rect 11394 41528 11406 41531
rect 11204 41500 11406 41528
rect 11204 41488 11210 41500
rect 11394 41497 11406 41500
rect 11440 41497 11452 41531
rect 12989 41531 13047 41537
rect 12989 41528 13001 41531
rect 11394 41491 11452 41497
rect 12544 41500 13001 41528
rect 12434 41460 12440 41472
rect 7668 41432 12440 41460
rect 12434 41420 12440 41432
rect 12492 41420 12498 41472
rect 12544 41469 12572 41500
rect 12989 41497 13001 41500
rect 13035 41497 13047 41531
rect 12989 41491 13047 41497
rect 20984 41531 21042 41537
rect 20984 41497 20996 41531
rect 21030 41528 21042 41531
rect 21082 41528 21088 41540
rect 21030 41500 21088 41528
rect 21030 41497 21042 41500
rect 20984 41491 21042 41497
rect 21082 41488 21088 41500
rect 21140 41488 21146 41540
rect 24044 41528 24072 41559
rect 25222 41556 25228 41568
rect 25280 41596 25286 41608
rect 26206 41596 26234 41636
rect 28994 41624 29000 41636
rect 29052 41664 29058 41676
rect 32953 41667 33011 41673
rect 32953 41664 32965 41667
rect 29052 41636 32965 41664
rect 29052 41624 29058 41636
rect 32953 41633 32965 41636
rect 32999 41633 33011 41667
rect 32953 41627 33011 41633
rect 27062 41596 27068 41608
rect 25280 41568 26234 41596
rect 27023 41568 27068 41596
rect 25280 41556 25286 41568
rect 27062 41556 27068 41568
rect 27120 41556 27126 41608
rect 27157 41599 27215 41605
rect 27157 41565 27169 41599
rect 27203 41596 27215 41599
rect 27430 41596 27436 41608
rect 27203 41568 27436 41596
rect 27203 41565 27215 41568
rect 27157 41559 27215 41565
rect 27430 41556 27436 41568
rect 27488 41556 27494 41608
rect 32968 41596 32996 41627
rect 34348 41596 34376 41695
rect 38562 41692 38568 41744
rect 38620 41732 38626 41744
rect 38620 41704 40448 41732
rect 38620 41692 38626 41704
rect 34790 41624 34796 41676
rect 34848 41664 34854 41676
rect 35161 41667 35219 41673
rect 35161 41664 35173 41667
rect 34848 41636 35173 41664
rect 34848 41624 34854 41636
rect 35161 41633 35173 41636
rect 35207 41633 35219 41667
rect 35161 41627 35219 41633
rect 38654 41624 38660 41676
rect 38712 41664 38718 41676
rect 40420 41673 40448 41704
rect 39117 41667 39175 41673
rect 39117 41664 39129 41667
rect 38712 41636 39129 41664
rect 38712 41624 38718 41636
rect 39117 41633 39129 41636
rect 39163 41633 39175 41667
rect 39117 41627 39175 41633
rect 40405 41667 40463 41673
rect 40405 41633 40417 41667
rect 40451 41633 40463 41667
rect 40405 41627 40463 41633
rect 35345 41599 35403 41605
rect 35345 41596 35357 41599
rect 32968 41568 33364 41596
rect 34348 41568 35357 41596
rect 33336 41540 33364 41568
rect 35345 41565 35357 41568
rect 35391 41565 35403 41599
rect 35345 41559 35403 41565
rect 37093 41599 37151 41605
rect 37093 41565 37105 41599
rect 37139 41596 37151 41599
rect 37182 41596 37188 41608
rect 37139 41568 37188 41596
rect 37139 41565 37151 41568
rect 37093 41559 37151 41565
rect 37182 41556 37188 41568
rect 37240 41556 37246 41608
rect 37366 41605 37372 41608
rect 37360 41596 37372 41605
rect 37327 41568 37372 41596
rect 37360 41559 37372 41568
rect 37366 41556 37372 41559
rect 37424 41556 37430 41608
rect 39298 41596 39304 41608
rect 39259 41568 39304 41596
rect 39298 41556 39304 41568
rect 39356 41556 39362 41608
rect 40678 41605 40684 41608
rect 40672 41596 40684 41605
rect 40639 41568 40684 41596
rect 40672 41559 40684 41568
rect 40678 41556 40684 41559
rect 40736 41556 40742 41608
rect 43257 41599 43315 41605
rect 43257 41565 43269 41599
rect 43303 41565 43315 41599
rect 43257 41559 43315 41565
rect 43524 41599 43582 41605
rect 43524 41565 43536 41599
rect 43570 41565 43582 41599
rect 43524 41559 43582 41565
rect 24826 41531 24884 41537
rect 24826 41528 24838 41531
rect 24044 41500 24838 41528
rect 24826 41497 24838 41500
rect 24872 41497 24884 41531
rect 27338 41528 27344 41540
rect 27299 41500 27344 41528
rect 24826 41491 24884 41497
rect 27338 41488 27344 41500
rect 27396 41488 27402 41540
rect 33220 41531 33278 41537
rect 33220 41497 33232 41531
rect 33266 41497 33278 41531
rect 33220 41491 33278 41497
rect 12529 41463 12587 41469
rect 12529 41429 12541 41463
rect 12575 41429 12587 41463
rect 13446 41460 13452 41472
rect 13407 41432 13452 41460
rect 12529 41423 12587 41429
rect 13446 41420 13452 41432
rect 13504 41420 13510 41472
rect 16301 41463 16359 41469
rect 16301 41429 16313 41463
rect 16347 41460 16359 41463
rect 16758 41460 16764 41472
rect 16347 41432 16764 41460
rect 16347 41429 16359 41432
rect 16301 41423 16359 41429
rect 16758 41420 16764 41432
rect 16816 41420 16822 41472
rect 22097 41463 22155 41469
rect 22097 41429 22109 41463
rect 22143 41460 22155 41463
rect 22738 41460 22744 41472
rect 22143 41432 22744 41460
rect 22143 41429 22155 41432
rect 22097 41423 22155 41429
rect 22738 41420 22744 41432
rect 22796 41420 22802 41472
rect 25774 41420 25780 41472
rect 25832 41460 25838 41472
rect 25961 41463 26019 41469
rect 25961 41460 25973 41463
rect 25832 41432 25973 41460
rect 25832 41420 25838 41432
rect 25961 41429 25973 41432
rect 26007 41429 26019 41463
rect 33244 41460 33272 41491
rect 33318 41488 33324 41540
rect 33376 41488 33382 41540
rect 35066 41528 35072 41540
rect 35027 41500 35072 41528
rect 35066 41488 35072 41500
rect 35124 41488 35130 41540
rect 39025 41531 39083 41537
rect 39025 41497 39037 41531
rect 39071 41528 39083 41531
rect 39114 41528 39120 41540
rect 39071 41500 39120 41528
rect 39071 41497 39083 41500
rect 39025 41491 39083 41497
rect 39114 41488 39120 41500
rect 39172 41488 39178 41540
rect 34974 41460 34980 41472
rect 33244 41432 34980 41460
rect 25961 41423 26019 41429
rect 34974 41420 34980 41432
rect 35032 41420 35038 41472
rect 38473 41463 38531 41469
rect 38473 41429 38485 41463
rect 38519 41460 38531 41463
rect 38746 41460 38752 41472
rect 38519 41432 38752 41460
rect 38519 41429 38531 41432
rect 38473 41423 38531 41429
rect 38746 41420 38752 41432
rect 38804 41420 38810 41472
rect 41785 41463 41843 41469
rect 41785 41429 41797 41463
rect 41831 41460 41843 41463
rect 42150 41460 42156 41472
rect 41831 41432 42156 41460
rect 41831 41429 41843 41432
rect 41785 41423 41843 41429
rect 42150 41420 42156 41432
rect 42208 41420 42214 41472
rect 43272 41460 43300 41559
rect 43438 41488 43444 41540
rect 43496 41528 43502 41540
rect 43548 41528 43576 41559
rect 43496 41500 43576 41528
rect 43496 41488 43502 41500
rect 45002 41460 45008 41472
rect 43272 41432 45008 41460
rect 45002 41420 45008 41432
rect 45060 41420 45066 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 12161 41259 12219 41265
rect 12161 41225 12173 41259
rect 12207 41256 12219 41259
rect 13262 41256 13268 41268
rect 12207 41228 13268 41256
rect 12207 41225 12219 41228
rect 12161 41219 12219 41225
rect 13262 41216 13268 41228
rect 13320 41216 13326 41268
rect 22094 41216 22100 41268
rect 22152 41256 22158 41268
rect 23382 41256 23388 41268
rect 22152 41228 23388 41256
rect 22152 41216 22158 41228
rect 23382 41216 23388 41228
rect 23440 41216 23446 41268
rect 25041 41259 25099 41265
rect 25041 41225 25053 41259
rect 25087 41256 25099 41259
rect 25087 41228 25544 41256
rect 25087 41225 25099 41228
rect 25041 41219 25099 41225
rect 22738 41188 22744 41200
rect 22699 41160 22744 41188
rect 22738 41148 22744 41160
rect 22796 41148 22802 41200
rect 9122 41120 9128 41132
rect 9083 41092 9128 41120
rect 9122 41080 9128 41092
rect 9180 41080 9186 41132
rect 9381 41123 9439 41129
rect 9381 41120 9393 41123
rect 9232 41092 9393 41120
rect 8570 41012 8576 41064
rect 8628 41052 8634 41064
rect 9232 41052 9260 41092
rect 9381 41089 9393 41092
rect 9427 41089 9439 41123
rect 11146 41120 11152 41132
rect 11107 41092 11152 41120
rect 9381 41083 9439 41089
rect 11146 41080 11152 41092
rect 11204 41080 11210 41132
rect 15194 41129 15200 41132
rect 13285 41123 13343 41129
rect 13285 41089 13297 41123
rect 13331 41120 13343 41123
rect 14001 41123 14059 41129
rect 14001 41120 14013 41123
rect 13331 41092 14013 41120
rect 13331 41089 13343 41092
rect 13285 41083 13343 41089
rect 14001 41089 14013 41092
rect 14047 41089 14059 41123
rect 14001 41083 14059 41089
rect 15188 41083 15200 41129
rect 15252 41120 15258 41132
rect 21082 41120 21088 41132
rect 15252 41092 15288 41120
rect 21043 41092 21088 41120
rect 15194 41080 15200 41083
rect 15252 41080 15258 41092
rect 21082 41080 21088 41092
rect 21140 41080 21146 41132
rect 23017 41123 23075 41129
rect 23017 41089 23029 41123
rect 23063 41089 23075 41123
rect 23400 41120 23428 41216
rect 25516 41197 25544 41228
rect 27338 41216 27344 41268
rect 27396 41256 27402 41268
rect 27525 41259 27583 41265
rect 27525 41256 27537 41259
rect 27396 41228 27537 41256
rect 27396 41216 27402 41228
rect 27525 41225 27537 41228
rect 27571 41256 27583 41259
rect 27982 41256 27988 41268
rect 27571 41228 27988 41256
rect 27571 41225 27583 41228
rect 27525 41219 27583 41225
rect 27982 41216 27988 41228
rect 28040 41216 28046 41268
rect 34609 41259 34667 41265
rect 34609 41225 34621 41259
rect 34655 41256 34667 41259
rect 35066 41256 35072 41268
rect 34655 41228 35072 41256
rect 34655 41225 34667 41228
rect 34609 41219 34667 41225
rect 35066 41216 35072 41228
rect 35124 41216 35130 41268
rect 43625 41259 43683 41265
rect 43625 41225 43637 41259
rect 43671 41256 43683 41259
rect 44174 41256 44180 41268
rect 43671 41228 44180 41256
rect 43671 41225 43683 41228
rect 43625 41219 43683 41225
rect 44174 41216 44180 41228
rect 44232 41216 44238 41268
rect 25501 41191 25559 41197
rect 25501 41157 25513 41191
rect 25547 41157 25559 41191
rect 25501 41151 25559 41157
rect 44760 41191 44818 41197
rect 44760 41157 44772 41191
rect 44806 41188 44818 41191
rect 45094 41188 45100 41200
rect 44806 41160 45100 41188
rect 44806 41157 44818 41160
rect 44760 41151 44818 41157
rect 45094 41148 45100 41160
rect 45152 41148 45158 41200
rect 23661 41123 23719 41129
rect 23661 41120 23673 41123
rect 23400 41092 23673 41120
rect 23017 41083 23075 41089
rect 23661 41089 23673 41092
rect 23707 41089 23719 41123
rect 23661 41083 23719 41089
rect 23928 41123 23986 41129
rect 23928 41089 23940 41123
rect 23974 41120 23986 41123
rect 24486 41120 24492 41132
rect 23974 41092 24492 41120
rect 23974 41089 23986 41092
rect 23928 41083 23986 41089
rect 8628 41024 9260 41052
rect 13541 41055 13599 41061
rect 8628 41012 8634 41024
rect 13541 41021 13553 41055
rect 13587 41052 13599 41055
rect 13814 41052 13820 41064
rect 13587 41024 13820 41052
rect 13587 41021 13599 41024
rect 13541 41015 13599 41021
rect 13814 41012 13820 41024
rect 13872 41052 13878 41064
rect 14918 41052 14924 41064
rect 13872 41024 14924 41052
rect 13872 41012 13878 41024
rect 14918 41012 14924 41024
rect 14976 41012 14982 41064
rect 22922 41052 22928 41064
rect 22883 41024 22928 41052
rect 22922 41012 22928 41024
rect 22980 41012 22986 41064
rect 23032 41052 23060 41083
rect 24486 41080 24492 41092
rect 24544 41080 24550 41132
rect 25774 41120 25780 41132
rect 25735 41092 25780 41120
rect 25774 41080 25780 41092
rect 25832 41080 25838 41132
rect 28258 41080 28264 41132
rect 28316 41120 28322 41132
rect 28638 41123 28696 41129
rect 28638 41120 28650 41123
rect 28316 41092 28650 41120
rect 28316 41080 28322 41092
rect 28638 41089 28650 41092
rect 28684 41089 28696 41123
rect 28638 41083 28696 41089
rect 28905 41123 28963 41129
rect 28905 41089 28917 41123
rect 28951 41120 28963 41123
rect 28994 41120 29000 41132
rect 28951 41092 29000 41120
rect 28951 41089 28963 41092
rect 28905 41083 28963 41089
rect 28994 41080 29000 41092
rect 29052 41080 29058 41132
rect 30285 41123 30343 41129
rect 30285 41089 30297 41123
rect 30331 41120 30343 41123
rect 30374 41120 30380 41132
rect 30331 41092 30380 41120
rect 30331 41089 30343 41092
rect 30285 41083 30343 41089
rect 30374 41080 30380 41092
rect 30432 41080 30438 41132
rect 33229 41123 33287 41129
rect 33229 41089 33241 41123
rect 33275 41120 33287 41123
rect 33318 41120 33324 41132
rect 33275 41092 33324 41120
rect 33275 41089 33287 41092
rect 33229 41083 33287 41089
rect 33318 41080 33324 41092
rect 33376 41080 33382 41132
rect 33502 41129 33508 41132
rect 33496 41083 33508 41129
rect 33560 41120 33566 41132
rect 33560 41092 33596 41120
rect 33502 41080 33508 41083
rect 33560 41080 33566 41092
rect 34974 41080 34980 41132
rect 35032 41120 35038 41132
rect 37734 41129 37740 41132
rect 35069 41123 35127 41129
rect 35069 41120 35081 41123
rect 35032 41092 35081 41120
rect 35032 41080 35038 41092
rect 35069 41089 35081 41092
rect 35115 41089 35127 41123
rect 35069 41083 35127 41089
rect 37728 41083 37740 41129
rect 37792 41120 37798 41132
rect 40856 41123 40914 41129
rect 37792 41092 37828 41120
rect 37734 41080 37740 41083
rect 37792 41080 37798 41092
rect 40856 41089 40868 41123
rect 40902 41120 40914 41123
rect 41322 41120 41328 41132
rect 40902 41092 41328 41120
rect 40902 41089 40914 41092
rect 40856 41083 40914 41089
rect 41322 41080 41328 41092
rect 41380 41080 41386 41132
rect 45002 41120 45008 41132
rect 44963 41092 45008 41120
rect 45002 41080 45008 41092
rect 45060 41080 45066 41132
rect 23566 41052 23572 41064
rect 23032 41024 23572 41052
rect 23566 41012 23572 41024
rect 23624 41012 23630 41064
rect 25590 41052 25596 41064
rect 25551 41024 25596 41052
rect 25590 41012 25596 41024
rect 25648 41012 25654 41064
rect 37274 41012 37280 41064
rect 37332 41052 37338 41064
rect 37461 41055 37519 41061
rect 37461 41052 37473 41055
rect 37332 41024 37473 41052
rect 37332 41012 37338 41024
rect 37461 41021 37473 41024
rect 37507 41021 37519 41055
rect 37461 41015 37519 41021
rect 40310 41012 40316 41064
rect 40368 41052 40374 41064
rect 40589 41055 40647 41061
rect 40589 41052 40601 41055
rect 40368 41024 40601 41052
rect 40368 41012 40374 41024
rect 40589 41021 40601 41024
rect 40635 41021 40647 41055
rect 40589 41015 40647 41021
rect 5534 40916 5540 40928
rect 5495 40888 5540 40916
rect 5534 40876 5540 40888
rect 5592 40876 5598 40928
rect 10505 40919 10563 40925
rect 10505 40885 10517 40919
rect 10551 40916 10563 40919
rect 11146 40916 11152 40928
rect 10551 40888 11152 40916
rect 10551 40885 10563 40888
rect 10505 40879 10563 40885
rect 11146 40876 11152 40888
rect 11204 40876 11210 40928
rect 16301 40919 16359 40925
rect 16301 40885 16313 40919
rect 16347 40916 16359 40919
rect 16850 40916 16856 40928
rect 16347 40888 16856 40916
rect 16347 40885 16359 40888
rect 16301 40879 16359 40885
rect 16850 40876 16856 40888
rect 16908 40876 16914 40928
rect 22189 40919 22247 40925
rect 22189 40885 22201 40919
rect 22235 40916 22247 40919
rect 22278 40916 22284 40928
rect 22235 40888 22284 40916
rect 22235 40885 22247 40888
rect 22189 40879 22247 40885
rect 22278 40876 22284 40888
rect 22336 40876 22342 40928
rect 23014 40916 23020 40928
rect 22975 40888 23020 40916
rect 23014 40876 23020 40888
rect 23072 40876 23078 40928
rect 23198 40916 23204 40928
rect 23159 40888 23204 40916
rect 23198 40876 23204 40888
rect 23256 40876 23262 40928
rect 25498 40916 25504 40928
rect 25459 40888 25504 40916
rect 25498 40876 25504 40888
rect 25556 40876 25562 40928
rect 25682 40876 25688 40928
rect 25740 40916 25746 40928
rect 25961 40919 26019 40925
rect 25961 40916 25973 40919
rect 25740 40888 25973 40916
rect 25740 40876 25746 40888
rect 25961 40885 25973 40888
rect 26007 40885 26019 40919
rect 30098 40916 30104 40928
rect 30059 40888 30104 40916
rect 25961 40879 26019 40885
rect 30098 40876 30104 40888
rect 30156 40876 30162 40928
rect 38841 40919 38899 40925
rect 38841 40885 38853 40919
rect 38887 40916 38899 40919
rect 39022 40916 39028 40928
rect 38887 40888 39028 40916
rect 38887 40885 38899 40888
rect 38841 40879 38899 40885
rect 39022 40876 39028 40888
rect 39080 40876 39086 40928
rect 40126 40916 40132 40928
rect 40087 40888 40132 40916
rect 40126 40876 40132 40888
rect 40184 40876 40190 40928
rect 41969 40919 42027 40925
rect 41969 40885 41981 40919
rect 42015 40916 42027 40919
rect 42426 40916 42432 40928
rect 42015 40888 42432 40916
rect 42015 40885 42027 40888
rect 41969 40879 42027 40885
rect 42426 40876 42432 40888
rect 42484 40876 42490 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 8570 40712 8576 40724
rect 8531 40684 8576 40712
rect 8570 40672 8576 40684
rect 8628 40672 8634 40724
rect 13170 40712 13176 40724
rect 13131 40684 13176 40712
rect 13170 40672 13176 40684
rect 13228 40672 13234 40724
rect 16758 40712 16764 40724
rect 16719 40684 16764 40712
rect 16758 40672 16764 40684
rect 16816 40672 16822 40724
rect 24486 40672 24492 40724
rect 24544 40712 24550 40724
rect 24581 40715 24639 40721
rect 24581 40712 24593 40715
rect 24544 40684 24593 40712
rect 24544 40672 24550 40684
rect 24581 40681 24593 40684
rect 24627 40681 24639 40715
rect 26326 40712 26332 40724
rect 26287 40684 26332 40712
rect 24581 40675 24639 40681
rect 26326 40672 26332 40684
rect 26384 40712 26390 40724
rect 27062 40712 27068 40724
rect 26384 40684 27068 40712
rect 26384 40672 26390 40684
rect 27062 40672 27068 40684
rect 27120 40712 27126 40724
rect 33502 40712 33508 40724
rect 27120 40684 27292 40712
rect 33463 40684 33508 40712
rect 27120 40672 27126 40684
rect 16301 40647 16359 40653
rect 16301 40613 16313 40647
rect 16347 40644 16359 40647
rect 16347 40616 16574 40644
rect 16347 40613 16359 40616
rect 16301 40607 16359 40613
rect 5258 40576 5264 40588
rect 5219 40548 5264 40576
rect 5258 40536 5264 40548
rect 5316 40536 5322 40588
rect 9122 40576 9128 40588
rect 9083 40548 9128 40576
rect 9122 40536 9128 40548
rect 9180 40536 9186 40588
rect 13814 40536 13820 40588
rect 13872 40576 13878 40588
rect 14918 40576 14924 40588
rect 13872 40548 14924 40576
rect 13872 40536 13878 40548
rect 14918 40536 14924 40548
rect 14976 40536 14982 40588
rect 5534 40517 5540 40520
rect 5528 40508 5540 40517
rect 5495 40480 5540 40508
rect 5528 40471 5540 40480
rect 5534 40468 5540 40471
rect 5592 40468 5598 40520
rect 9398 40517 9404 40520
rect 9392 40508 9404 40517
rect 9359 40480 9404 40508
rect 9392 40471 9404 40480
rect 9398 40468 9404 40471
rect 9456 40468 9462 40520
rect 11790 40508 11796 40520
rect 11751 40480 11796 40508
rect 11790 40468 11796 40480
rect 11848 40468 11854 40520
rect 12066 40517 12072 40520
rect 12060 40508 12072 40517
rect 12027 40480 12072 40508
rect 12060 40471 12072 40480
rect 12066 40468 12072 40471
rect 12124 40468 12130 40520
rect 14461 40511 14519 40517
rect 14461 40477 14473 40511
rect 14507 40508 14519 40511
rect 15177 40511 15235 40517
rect 15177 40508 15189 40511
rect 14507 40480 15189 40508
rect 14507 40477 14519 40480
rect 14461 40471 14519 40477
rect 15177 40477 15189 40480
rect 15223 40477 15235 40511
rect 16546 40508 16574 40616
rect 16850 40576 16856 40588
rect 16811 40548 16856 40576
rect 16850 40536 16856 40548
rect 16908 40536 16914 40588
rect 22094 40536 22100 40588
rect 22152 40576 22158 40588
rect 22281 40579 22339 40585
rect 22281 40576 22293 40579
rect 22152 40548 22293 40576
rect 22152 40536 22158 40548
rect 22281 40545 22293 40548
rect 22327 40545 22339 40579
rect 22281 40539 22339 40545
rect 25869 40579 25927 40585
rect 25869 40545 25881 40579
rect 25915 40576 25927 40579
rect 25915 40548 26556 40576
rect 27264 40562 27292 40684
rect 33502 40672 33508 40684
rect 33560 40672 33566 40724
rect 38746 40712 38752 40724
rect 38707 40684 38752 40712
rect 38746 40672 38752 40684
rect 38804 40672 38810 40724
rect 39114 40672 39120 40724
rect 39172 40712 39178 40724
rect 39209 40715 39267 40721
rect 39209 40712 39221 40715
rect 39172 40684 39221 40712
rect 39172 40672 39178 40684
rect 39209 40681 39221 40684
rect 39255 40681 39267 40715
rect 42150 40712 42156 40724
rect 42111 40684 42156 40712
rect 39209 40675 39267 40681
rect 42150 40672 42156 40684
rect 42208 40672 42214 40724
rect 42610 40712 42616 40724
rect 42571 40684 42616 40712
rect 42610 40672 42616 40684
rect 42668 40672 42674 40724
rect 38289 40647 38347 40653
rect 38289 40613 38301 40647
rect 38335 40644 38347 40647
rect 38335 40616 38884 40644
rect 38335 40613 38347 40616
rect 38289 40607 38347 40613
rect 38856 40585 38884 40616
rect 38841 40579 38899 40585
rect 25915 40545 25927 40548
rect 25869 40539 25927 40545
rect 17037 40511 17095 40517
rect 17037 40508 17049 40511
rect 16546 40480 17049 40508
rect 15177 40471 15235 40477
rect 17037 40477 17049 40480
rect 17083 40477 17095 40511
rect 17037 40471 17095 40477
rect 21729 40511 21787 40517
rect 21729 40477 21741 40511
rect 21775 40508 21787 40511
rect 22462 40508 22468 40520
rect 21775 40480 22468 40508
rect 21775 40477 21787 40480
rect 21729 40471 21787 40477
rect 22462 40468 22468 40480
rect 22520 40468 22526 40520
rect 23198 40468 23204 40520
rect 23256 40508 23262 40520
rect 25501 40511 25559 40517
rect 25501 40508 25513 40511
rect 23256 40480 25513 40508
rect 23256 40468 23262 40480
rect 25501 40477 25513 40480
rect 25547 40477 25559 40511
rect 25682 40508 25688 40520
rect 25643 40480 25688 40508
rect 25501 40471 25559 40477
rect 25682 40468 25688 40480
rect 25740 40468 25746 40520
rect 26528 40517 26556 40548
rect 38841 40545 38853 40579
rect 38887 40545 38899 40579
rect 38841 40539 38899 40545
rect 26329 40511 26387 40517
rect 26329 40477 26341 40511
rect 26375 40477 26387 40511
rect 26329 40471 26387 40477
rect 26513 40511 26571 40517
rect 26513 40477 26525 40511
rect 26559 40508 26571 40511
rect 27430 40508 27436 40520
rect 26559 40502 27292 40508
rect 27356 40502 27436 40508
rect 26559 40480 27436 40502
rect 26559 40477 26571 40480
rect 26513 40471 26571 40477
rect 27264 40474 27384 40480
rect 11808 40440 11836 40468
rect 13814 40440 13820 40452
rect 11808 40412 13820 40440
rect 13814 40400 13820 40412
rect 13872 40400 13878 40452
rect 16758 40440 16764 40452
rect 16719 40412 16764 40440
rect 16758 40400 16764 40412
rect 16816 40400 16822 40452
rect 24029 40443 24087 40449
rect 24029 40409 24041 40443
rect 24075 40440 24087 40443
rect 24210 40440 24216 40452
rect 24075 40412 24216 40440
rect 24075 40409 24087 40412
rect 24029 40403 24087 40409
rect 24210 40400 24216 40412
rect 24268 40440 24274 40452
rect 24762 40440 24768 40452
rect 24268 40412 24768 40440
rect 24268 40400 24274 40412
rect 24762 40400 24768 40412
rect 24820 40400 24826 40452
rect 26344 40440 26372 40471
rect 27430 40468 27436 40480
rect 27488 40468 27494 40520
rect 27893 40511 27951 40517
rect 27893 40477 27905 40511
rect 27939 40477 27951 40511
rect 27893 40471 27951 40477
rect 27522 40440 27528 40452
rect 26344 40412 27528 40440
rect 27522 40400 27528 40412
rect 27580 40440 27586 40452
rect 27908 40440 27936 40471
rect 27982 40468 27988 40520
rect 28040 40508 28046 40520
rect 28040 40480 28085 40508
rect 28040 40468 28046 40480
rect 29730 40468 29736 40520
rect 29788 40508 29794 40520
rect 30098 40517 30104 40520
rect 29825 40511 29883 40517
rect 29825 40508 29837 40511
rect 29788 40480 29837 40508
rect 29788 40468 29794 40480
rect 29825 40477 29837 40480
rect 29871 40477 29883 40511
rect 30092 40508 30104 40517
rect 30059 40480 30104 40508
rect 29825 40471 29883 40477
rect 30092 40471 30104 40480
rect 30098 40468 30104 40471
rect 30156 40468 30162 40520
rect 36449 40511 36507 40517
rect 36449 40477 36461 40511
rect 36495 40477 36507 40511
rect 36449 40471 36507 40477
rect 36909 40511 36967 40517
rect 36909 40477 36921 40511
rect 36955 40508 36967 40511
rect 39022 40508 39028 40520
rect 36955 40480 37320 40508
rect 38983 40480 39028 40508
rect 36955 40477 36967 40480
rect 36909 40471 36967 40477
rect 27580 40412 27936 40440
rect 36464 40440 36492 40471
rect 37292 40452 37320 40480
rect 39022 40468 39028 40480
rect 39080 40468 39086 40520
rect 40310 40508 40316 40520
rect 40271 40480 40316 40508
rect 40310 40468 40316 40480
rect 40368 40468 40374 40520
rect 41782 40468 41788 40520
rect 41840 40508 41846 40520
rect 42337 40511 42395 40517
rect 42337 40508 42349 40511
rect 41840 40480 42349 40508
rect 41840 40468 41846 40480
rect 42337 40477 42349 40480
rect 42383 40477 42395 40511
rect 42337 40471 42395 40477
rect 42426 40468 42432 40520
rect 42484 40508 42490 40520
rect 42484 40480 42529 40508
rect 42484 40468 42490 40480
rect 37154 40443 37212 40449
rect 37154 40440 37166 40443
rect 36464 40412 37166 40440
rect 27580 40400 27586 40412
rect 37154 40409 37166 40412
rect 37200 40409 37212 40443
rect 37154 40403 37212 40409
rect 37274 40400 37280 40452
rect 37332 40400 37338 40452
rect 38749 40443 38807 40449
rect 38749 40409 38761 40443
rect 38795 40440 38807 40443
rect 38838 40440 38844 40452
rect 38795 40412 38844 40440
rect 38795 40409 38807 40412
rect 38749 40403 38807 40409
rect 38838 40400 38844 40412
rect 38896 40400 38902 40452
rect 40586 40449 40592 40452
rect 40580 40403 40592 40449
rect 40644 40440 40650 40452
rect 42153 40443 42211 40449
rect 40644 40412 40680 40440
rect 40586 40400 40592 40403
rect 40644 40400 40650 40412
rect 42153 40409 42165 40443
rect 42199 40409 42211 40443
rect 42153 40403 42211 40409
rect 6641 40375 6699 40381
rect 6641 40341 6653 40375
rect 6687 40372 6699 40375
rect 6914 40372 6920 40384
rect 6687 40344 6920 40372
rect 6687 40341 6699 40344
rect 6641 40335 6699 40341
rect 6914 40332 6920 40344
rect 6972 40332 6978 40384
rect 10505 40375 10563 40381
rect 10505 40341 10517 40375
rect 10551 40372 10563 40375
rect 11238 40372 11244 40384
rect 10551 40344 11244 40372
rect 10551 40341 10563 40344
rect 10505 40335 10563 40341
rect 11238 40332 11244 40344
rect 11296 40332 11302 40384
rect 17218 40372 17224 40384
rect 17179 40344 17224 40372
rect 17218 40332 17224 40344
rect 17276 40332 17282 40384
rect 26694 40372 26700 40384
rect 26655 40344 26700 40372
rect 26694 40332 26700 40344
rect 26752 40332 26758 40384
rect 27776 40375 27834 40381
rect 27776 40341 27788 40375
rect 27822 40372 27834 40375
rect 28442 40372 28448 40384
rect 27822 40344 28448 40372
rect 27822 40341 27834 40344
rect 27776 40335 27834 40341
rect 28442 40332 28448 40344
rect 28500 40332 28506 40384
rect 31202 40372 31208 40384
rect 31163 40344 31208 40372
rect 31202 40332 31208 40344
rect 31260 40332 31266 40384
rect 41693 40375 41751 40381
rect 41693 40341 41705 40375
rect 41739 40372 41751 40375
rect 42168 40372 42196 40403
rect 41739 40344 42196 40372
rect 41739 40341 41751 40344
rect 41693 40335 41751 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 7190 40168 7196 40180
rect 7151 40140 7196 40168
rect 7190 40128 7196 40140
rect 7248 40128 7254 40180
rect 12434 40128 12440 40180
rect 12492 40168 12498 40180
rect 12713 40171 12771 40177
rect 12713 40168 12725 40171
rect 12492 40140 12725 40168
rect 12492 40128 12498 40140
rect 12713 40137 12725 40140
rect 12759 40137 12771 40171
rect 12713 40131 12771 40137
rect 12912 40140 16574 40168
rect 10505 40103 10563 40109
rect 10505 40069 10517 40103
rect 10551 40100 10563 40103
rect 10551 40072 11100 40100
rect 10551 40069 10563 40072
rect 10505 40063 10563 40069
rect 6825 40035 6883 40041
rect 6825 40001 6837 40035
rect 6871 40032 6883 40035
rect 7650 40032 7656 40044
rect 6871 40004 7656 40032
rect 6871 40001 6883 40004
rect 6825 39995 6883 40001
rect 7650 39992 7656 40004
rect 7708 39992 7714 40044
rect 8754 40032 8760 40044
rect 8715 40004 8760 40032
rect 8754 39992 8760 40004
rect 8812 39992 8818 40044
rect 6638 39924 6644 39976
rect 6696 39964 6702 39976
rect 6917 39967 6975 39973
rect 6917 39964 6929 39967
rect 6696 39936 6929 39964
rect 6696 39924 6702 39936
rect 6917 39933 6929 39936
rect 6963 39933 6975 39967
rect 6917 39927 6975 39933
rect 11072 39908 11100 40072
rect 12912 40041 12940 40140
rect 13814 40100 13820 40112
rect 13775 40072 13820 40100
rect 13814 40060 13820 40072
rect 13872 40060 13878 40112
rect 16546 40100 16574 40140
rect 22922 40128 22928 40180
rect 22980 40168 22986 40180
rect 23385 40171 23443 40177
rect 23385 40168 23397 40171
rect 22980 40140 23397 40168
rect 22980 40128 22986 40140
rect 23385 40137 23397 40140
rect 23431 40137 23443 40171
rect 23385 40131 23443 40137
rect 26605 40171 26663 40177
rect 26605 40137 26617 40171
rect 26651 40168 26663 40171
rect 28258 40168 28264 40180
rect 26651 40140 27844 40168
rect 28219 40140 28264 40168
rect 26651 40137 26663 40140
rect 26605 40131 26663 40137
rect 17218 40100 17224 40112
rect 16546 40072 17224 40100
rect 17218 40060 17224 40072
rect 17276 40060 17282 40112
rect 26694 40060 26700 40112
rect 26752 40100 26758 40112
rect 26752 40072 27384 40100
rect 26752 40060 26758 40072
rect 12897 40035 12955 40041
rect 12897 40001 12909 40035
rect 12943 40001 12955 40035
rect 13170 40032 13176 40044
rect 13131 40004 13176 40032
rect 12897 39995 12955 40001
rect 13170 39992 13176 40004
rect 13228 39992 13234 40044
rect 15381 40035 15439 40041
rect 15381 40001 15393 40035
rect 15427 40032 15439 40035
rect 15841 40035 15899 40041
rect 15841 40032 15853 40035
rect 15427 40004 15853 40032
rect 15427 40001 15439 40004
rect 15381 39995 15439 40001
rect 15841 40001 15853 40004
rect 15887 40001 15899 40035
rect 15841 39995 15899 40001
rect 22005 40035 22063 40041
rect 22005 40001 22017 40035
rect 22051 40032 22063 40035
rect 22094 40032 22100 40044
rect 22051 40004 22100 40032
rect 22051 40001 22063 40004
rect 22005 39995 22063 40001
rect 13081 39967 13139 39973
rect 13081 39933 13093 39967
rect 13127 39964 13139 39967
rect 13538 39964 13544 39976
rect 13127 39936 13544 39964
rect 13127 39933 13139 39936
rect 13081 39927 13139 39933
rect 13538 39924 13544 39936
rect 13596 39924 13602 39976
rect 11054 39896 11060 39908
rect 10967 39868 11060 39896
rect 11054 39856 11060 39868
rect 11112 39896 11118 39908
rect 15396 39896 15424 39995
rect 22094 39992 22100 40004
rect 22152 39992 22158 40044
rect 22278 40041 22284 40044
rect 22272 40032 22284 40041
rect 22239 40004 22284 40032
rect 22272 39995 22284 40004
rect 22278 39992 22284 39995
rect 22336 39992 22342 40044
rect 25222 40032 25228 40044
rect 25183 40004 25228 40032
rect 25222 39992 25228 40004
rect 25280 39992 25286 40044
rect 27356 40041 27384 40072
rect 25492 40035 25550 40041
rect 25492 40001 25504 40035
rect 25538 40032 25550 40035
rect 27157 40035 27215 40041
rect 27157 40032 27169 40035
rect 25538 40004 27169 40032
rect 25538 40001 25550 40004
rect 25492 39995 25550 40001
rect 27157 40001 27169 40004
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 27341 40035 27399 40041
rect 27341 40001 27353 40035
rect 27387 40001 27399 40035
rect 27614 40032 27620 40044
rect 27575 40004 27620 40032
rect 27341 39995 27399 40001
rect 27614 39992 27620 40004
rect 27672 39992 27678 40044
rect 27706 39992 27712 40044
rect 27764 40032 27770 40044
rect 27816 40041 27844 40140
rect 28258 40128 28264 40140
rect 28316 40128 28322 40180
rect 30374 40168 30380 40180
rect 30335 40140 30380 40168
rect 30374 40128 30380 40140
rect 30432 40128 30438 40180
rect 38838 40168 38844 40180
rect 38799 40140 38844 40168
rect 38838 40128 38844 40140
rect 38896 40128 38902 40180
rect 41782 40168 41788 40180
rect 41743 40140 41788 40168
rect 41782 40128 41788 40140
rect 41840 40128 41846 40180
rect 40126 40060 40132 40112
rect 40184 40100 40190 40112
rect 40650 40103 40708 40109
rect 40650 40100 40662 40103
rect 40184 40072 40662 40100
rect 40184 40060 40190 40072
rect 40650 40069 40662 40072
rect 40696 40069 40708 40103
rect 40650 40063 40708 40069
rect 27801 40035 27859 40041
rect 27801 40032 27813 40035
rect 27764 40004 27813 40032
rect 27764 39992 27770 40004
rect 27801 40001 27813 40004
rect 27847 40001 27859 40035
rect 28442 40032 28448 40044
rect 28403 40004 28448 40032
rect 27801 39995 27859 40001
rect 28442 39992 28448 40004
rect 28500 40032 28506 40044
rect 29917 40035 29975 40041
rect 28500 40004 28856 40032
rect 28500 39992 28506 40004
rect 27982 39924 27988 39976
rect 28040 39964 28046 39976
rect 28721 39967 28779 39973
rect 28721 39964 28733 39967
rect 28040 39936 28733 39964
rect 28040 39924 28046 39936
rect 28721 39933 28733 39936
rect 28767 39933 28779 39967
rect 28721 39927 28779 39933
rect 11112 39868 15424 39896
rect 11112 39856 11118 39868
rect 27522 39856 27528 39908
rect 27580 39896 27586 39908
rect 28629 39899 28687 39905
rect 28629 39896 28641 39899
rect 27580 39868 28641 39896
rect 27580 39856 27586 39868
rect 28629 39865 28641 39868
rect 28675 39865 28687 39899
rect 28828 39896 28856 40004
rect 29917 40001 29929 40035
rect 29963 40032 29975 40035
rect 30558 40032 30564 40044
rect 29963 40004 30564 40032
rect 29963 40001 29975 40004
rect 29917 39995 29975 40001
rect 30558 39992 30564 40004
rect 30616 40032 30622 40044
rect 31202 40032 31208 40044
rect 30616 40004 31208 40032
rect 30616 39992 30622 40004
rect 31202 39992 31208 40004
rect 31260 39992 31266 40044
rect 36909 40035 36967 40041
rect 36909 40001 36921 40035
rect 36955 40032 36967 40035
rect 37717 40035 37775 40041
rect 37717 40032 37729 40035
rect 36955 40004 37729 40032
rect 36955 40001 36967 40004
rect 36909 39995 36967 40001
rect 37717 40001 37729 40004
rect 37763 40001 37775 40035
rect 37717 39995 37775 40001
rect 37274 39924 37280 39976
rect 37332 39964 37338 39976
rect 37461 39967 37519 39973
rect 37461 39964 37473 39967
rect 37332 39936 37473 39964
rect 37332 39924 37338 39936
rect 37461 39933 37473 39936
rect 37507 39933 37519 39967
rect 37461 39927 37519 39933
rect 40310 39924 40316 39976
rect 40368 39964 40374 39976
rect 40405 39967 40463 39973
rect 40405 39964 40417 39967
rect 40368 39936 40417 39964
rect 40368 39924 40374 39936
rect 40405 39933 40417 39936
rect 40451 39933 40463 39967
rect 40405 39927 40463 39933
rect 30193 39899 30251 39905
rect 30193 39896 30205 39899
rect 28828 39868 30205 39896
rect 28629 39859 28687 39865
rect 30193 39865 30205 39868
rect 30239 39865 30251 39899
rect 30193 39859 30251 39865
rect 5534 39788 5540 39840
rect 5592 39828 5598 39840
rect 5629 39831 5687 39837
rect 5629 39828 5641 39831
rect 5592 39800 5641 39828
rect 5592 39788 5598 39800
rect 5629 39797 5641 39800
rect 5675 39797 5687 39831
rect 5629 39791 5687 39797
rect 6914 39788 6920 39840
rect 6972 39828 6978 39840
rect 8297 39831 8355 39837
rect 6972 39800 7017 39828
rect 6972 39788 6978 39800
rect 8297 39797 8309 39831
rect 8343 39828 8355 39831
rect 9214 39828 9220 39840
rect 8343 39800 9220 39828
rect 8343 39797 8355 39800
rect 8297 39791 8355 39797
rect 9214 39788 9220 39800
rect 9272 39788 9278 39840
rect 13173 39831 13231 39837
rect 13173 39797 13185 39831
rect 13219 39828 13231 39831
rect 13446 39828 13452 39840
rect 13219 39800 13452 39828
rect 13219 39797 13231 39800
rect 13173 39791 13231 39797
rect 13446 39788 13452 39800
rect 13504 39788 13510 39840
rect 24210 39828 24216 39840
rect 24171 39800 24216 39828
rect 24210 39788 24216 39800
rect 24268 39788 24274 39840
rect 40420 39828 40448 39927
rect 40678 39828 40684 39840
rect 40420 39800 40684 39828
rect 40678 39788 40684 39800
rect 40736 39788 40742 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 6638 39624 6644 39636
rect 6599 39596 6644 39624
rect 6638 39584 6644 39596
rect 6696 39584 6702 39636
rect 7282 39624 7288 39636
rect 7243 39596 7288 39624
rect 7282 39584 7288 39596
rect 7340 39584 7346 39636
rect 7650 39624 7656 39636
rect 7611 39596 7656 39624
rect 7650 39584 7656 39596
rect 7708 39584 7714 39636
rect 11146 39624 11152 39636
rect 11107 39596 11152 39624
rect 11146 39584 11152 39596
rect 11204 39584 11210 39636
rect 11333 39627 11391 39633
rect 11333 39593 11345 39627
rect 11379 39624 11391 39627
rect 13170 39624 13176 39636
rect 11379 39596 13176 39624
rect 11379 39593 11391 39596
rect 11333 39587 11391 39593
rect 13170 39584 13176 39596
rect 13228 39584 13234 39636
rect 14461 39627 14519 39633
rect 14461 39593 14473 39627
rect 14507 39624 14519 39627
rect 15194 39624 15200 39636
rect 14507 39596 15200 39624
rect 14507 39593 14519 39596
rect 14461 39587 14519 39593
rect 15194 39584 15200 39596
rect 15252 39584 15258 39636
rect 16393 39627 16451 39633
rect 16393 39593 16405 39627
rect 16439 39624 16451 39627
rect 16758 39624 16764 39636
rect 16439 39596 16764 39624
rect 16439 39593 16451 39596
rect 16393 39587 16451 39593
rect 16758 39584 16764 39596
rect 16816 39584 16822 39636
rect 23566 39624 23572 39636
rect 23527 39596 23572 39624
rect 23566 39584 23572 39596
rect 23624 39584 23630 39636
rect 37645 39627 37703 39633
rect 37645 39593 37657 39627
rect 37691 39624 37703 39627
rect 37734 39624 37740 39636
rect 37691 39596 37740 39624
rect 37691 39593 37703 39596
rect 37645 39587 37703 39593
rect 37734 39584 37740 39596
rect 37792 39584 37798 39636
rect 40586 39584 40592 39636
rect 40644 39624 40650 39636
rect 40681 39627 40739 39633
rect 40681 39624 40693 39627
rect 40644 39596 40693 39624
rect 40644 39584 40650 39596
rect 40681 39593 40693 39596
rect 40727 39593 40739 39627
rect 41322 39624 41328 39636
rect 41283 39596 41328 39624
rect 40681 39587 40739 39593
rect 41322 39584 41328 39596
rect 41380 39584 41386 39636
rect 5258 39488 5264 39500
rect 5219 39460 5264 39488
rect 5258 39448 5264 39460
rect 5316 39448 5322 39500
rect 7374 39488 7380 39500
rect 7335 39460 7380 39488
rect 7374 39448 7380 39460
rect 7432 39448 7438 39500
rect 14918 39448 14924 39500
rect 14976 39488 14982 39500
rect 15013 39491 15071 39497
rect 15013 39488 15025 39491
rect 14976 39460 15025 39488
rect 14976 39448 14982 39460
rect 15013 39457 15025 39460
rect 15059 39457 15071 39491
rect 15013 39451 15071 39457
rect 22094 39448 22100 39500
rect 22152 39488 22158 39500
rect 22189 39491 22247 39497
rect 22189 39488 22201 39491
rect 22152 39460 22201 39488
rect 22152 39448 22158 39460
rect 22189 39457 22201 39460
rect 22235 39457 22247 39491
rect 22189 39451 22247 39457
rect 5534 39429 5540 39432
rect 5528 39420 5540 39429
rect 5495 39392 5540 39420
rect 5528 39383 5540 39392
rect 5534 39380 5540 39383
rect 5592 39380 5598 39432
rect 7466 39420 7472 39432
rect 7427 39392 7472 39420
rect 7466 39380 7472 39392
rect 7524 39380 7530 39432
rect 8297 39423 8355 39429
rect 8297 39389 8309 39423
rect 8343 39420 8355 39423
rect 8386 39420 8392 39432
rect 8343 39392 8392 39420
rect 8343 39389 8355 39392
rect 8297 39383 8355 39389
rect 8386 39380 8392 39392
rect 8444 39380 8450 39432
rect 8754 39380 8760 39432
rect 8812 39420 8818 39432
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 8812 39392 9137 39420
rect 8812 39380 8818 39392
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9214 39380 9220 39432
rect 9272 39420 9278 39432
rect 9381 39423 9439 39429
rect 9381 39420 9393 39423
rect 9272 39392 9393 39420
rect 9272 39380 9278 39392
rect 9381 39389 9393 39392
rect 9427 39389 9439 39423
rect 10965 39423 11023 39429
rect 10965 39420 10977 39423
rect 9381 39383 9439 39389
rect 10520 39392 10977 39420
rect 7190 39352 7196 39364
rect 7151 39324 7196 39352
rect 7190 39312 7196 39324
rect 7248 39312 7254 39364
rect 10520 39293 10548 39392
rect 10965 39389 10977 39392
rect 11011 39389 11023 39423
rect 10965 39383 11023 39389
rect 11149 39423 11207 39429
rect 11149 39389 11161 39423
rect 11195 39420 11207 39423
rect 11238 39420 11244 39432
rect 11195 39392 11244 39420
rect 11195 39389 11207 39392
rect 11149 39383 11207 39389
rect 11238 39380 11244 39392
rect 11296 39380 11302 39432
rect 15286 39429 15292 39432
rect 15280 39420 15292 39429
rect 15247 39392 15292 39420
rect 15280 39383 15292 39392
rect 15286 39380 15292 39383
rect 15344 39380 15350 39432
rect 22462 39429 22468 39432
rect 22456 39383 22468 39429
rect 22520 39420 22526 39432
rect 22520 39392 22556 39420
rect 22462 39380 22468 39383
rect 22520 39380 22526 39392
rect 10505 39287 10563 39293
rect 10505 39253 10517 39287
rect 10551 39253 10563 39287
rect 10505 39247 10563 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 9585 39083 9643 39089
rect 9585 39080 9597 39083
rect 7300 39052 9597 39080
rect 7300 39021 7328 39052
rect 9585 39049 9597 39052
rect 9631 39080 9643 39083
rect 11054 39080 11060 39092
rect 9631 39052 11060 39080
rect 9631 39049 9643 39052
rect 9585 39043 9643 39049
rect 11054 39040 11060 39052
rect 11112 39040 11118 39092
rect 27157 39083 27215 39089
rect 27157 39049 27169 39083
rect 27203 39080 27215 39083
rect 27522 39080 27528 39092
rect 27203 39052 27528 39080
rect 27203 39049 27215 39052
rect 27157 39043 27215 39049
rect 27522 39040 27528 39052
rect 27580 39040 27586 39092
rect 7285 39015 7343 39021
rect 7285 38981 7297 39015
rect 7331 38981 7343 39015
rect 27341 39015 27399 39021
rect 27341 39012 27353 39015
rect 7285 38975 7343 38981
rect 27264 38984 27353 39012
rect 22094 38904 22100 38956
rect 22152 38944 22158 38956
rect 23201 38947 23259 38953
rect 23201 38944 23213 38947
rect 22152 38916 23213 38944
rect 22152 38904 22158 38916
rect 23201 38913 23213 38916
rect 23247 38944 23259 38947
rect 23290 38944 23296 38956
rect 23247 38916 23296 38944
rect 23247 38913 23259 38916
rect 23201 38907 23259 38913
rect 23290 38904 23296 38916
rect 23348 38904 23354 38956
rect 23474 38953 23480 38956
rect 23468 38907 23480 38953
rect 23532 38944 23538 38956
rect 23532 38916 23568 38944
rect 23474 38904 23480 38907
rect 23532 38904 23538 38916
rect 27264 38876 27292 38984
rect 27341 38981 27353 38984
rect 27387 38981 27399 39015
rect 27706 39012 27712 39024
rect 27667 38984 27712 39012
rect 27341 38975 27399 38981
rect 27706 38972 27712 38984
rect 27764 38972 27770 39024
rect 27430 38944 27436 38956
rect 27391 38916 27436 38944
rect 27430 38904 27436 38916
rect 27488 38904 27494 38956
rect 27525 38947 27583 38953
rect 27525 38913 27537 38947
rect 27571 38944 27583 38947
rect 28166 38944 28172 38956
rect 27571 38916 28172 38944
rect 27571 38913 27583 38916
rect 27525 38907 27583 38913
rect 28166 38904 28172 38916
rect 28224 38904 28230 38956
rect 30558 38944 30564 38956
rect 30519 38916 30564 38944
rect 30558 38904 30564 38916
rect 30616 38904 30622 38956
rect 30745 38947 30803 38953
rect 30745 38913 30757 38947
rect 30791 38944 30803 38947
rect 30834 38944 30840 38956
rect 30791 38916 30840 38944
rect 30791 38913 30803 38916
rect 30745 38907 30803 38913
rect 30834 38904 30840 38916
rect 30892 38904 30898 38956
rect 40770 38944 40776 38956
rect 40731 38916 40776 38944
rect 40770 38904 40776 38916
rect 40828 38904 40834 38956
rect 40957 38947 41015 38953
rect 40957 38913 40969 38947
rect 41003 38944 41015 38947
rect 41598 38944 41604 38956
rect 41003 38916 41604 38944
rect 41003 38913 41015 38916
rect 40957 38907 41015 38913
rect 41598 38904 41604 38916
rect 41656 38904 41662 38956
rect 28350 38876 28356 38888
rect 27264 38848 28356 38876
rect 28350 38836 28356 38848
rect 28408 38836 28414 38888
rect 5258 38768 5264 38820
rect 5316 38808 5322 38820
rect 6914 38808 6920 38820
rect 5316 38780 6920 38808
rect 5316 38768 5322 38780
rect 6914 38768 6920 38780
rect 6972 38768 6978 38820
rect 5534 38700 5540 38752
rect 5592 38740 5598 38752
rect 5721 38743 5779 38749
rect 5721 38740 5733 38743
rect 5592 38712 5733 38740
rect 5592 38700 5598 38712
rect 5721 38709 5733 38712
rect 5767 38709 5779 38743
rect 5721 38703 5779 38709
rect 6733 38743 6791 38749
rect 6733 38709 6745 38743
rect 6779 38740 6791 38743
rect 7006 38740 7012 38752
rect 6779 38712 7012 38740
rect 6779 38709 6791 38712
rect 6733 38703 6791 38709
rect 7006 38700 7012 38712
rect 7064 38700 7070 38752
rect 8754 38740 8760 38752
rect 8715 38712 8760 38740
rect 8754 38700 8760 38712
rect 8812 38700 8818 38752
rect 11698 38740 11704 38752
rect 11659 38712 11704 38740
rect 11698 38700 11704 38712
rect 11756 38700 11762 38752
rect 24578 38740 24584 38752
rect 24539 38712 24584 38740
rect 24578 38700 24584 38712
rect 24636 38700 24642 38752
rect 30653 38743 30711 38749
rect 30653 38709 30665 38743
rect 30699 38740 30711 38743
rect 30742 38740 30748 38752
rect 30699 38712 30748 38740
rect 30699 38709 30711 38712
rect 30653 38703 30711 38709
rect 30742 38700 30748 38712
rect 30800 38700 30806 38752
rect 36630 38700 36636 38752
rect 36688 38740 36694 38752
rect 36725 38743 36783 38749
rect 36725 38740 36737 38743
rect 36688 38712 36737 38740
rect 36688 38700 36694 38712
rect 36725 38709 36737 38712
rect 36771 38709 36783 38743
rect 36725 38703 36783 38709
rect 41141 38743 41199 38749
rect 41141 38709 41153 38743
rect 41187 38740 41199 38743
rect 41966 38740 41972 38752
rect 41187 38712 41972 38740
rect 41187 38709 41199 38712
rect 41141 38703 41199 38709
rect 41966 38700 41972 38712
rect 42024 38700 42030 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 7101 38539 7159 38545
rect 7101 38505 7113 38539
rect 7147 38536 7159 38539
rect 7466 38536 7472 38548
rect 7147 38508 7472 38536
rect 7147 38505 7159 38508
rect 7101 38499 7159 38505
rect 7466 38496 7472 38508
rect 7524 38496 7530 38548
rect 12621 38539 12679 38545
rect 12621 38505 12633 38539
rect 12667 38536 12679 38539
rect 13081 38539 13139 38545
rect 13081 38536 13093 38539
rect 12667 38508 13093 38536
rect 12667 38505 12679 38508
rect 12621 38499 12679 38505
rect 13081 38505 13093 38508
rect 13127 38505 13139 38539
rect 13538 38536 13544 38548
rect 13499 38508 13544 38536
rect 13081 38499 13139 38505
rect 13538 38496 13544 38508
rect 13596 38496 13602 38548
rect 23109 38539 23167 38545
rect 23109 38505 23121 38539
rect 23155 38536 23167 38539
rect 23474 38536 23480 38548
rect 23155 38508 23480 38536
rect 23155 38505 23167 38508
rect 23109 38499 23167 38505
rect 23474 38496 23480 38508
rect 23532 38496 23538 38548
rect 26881 38539 26939 38545
rect 26881 38505 26893 38539
rect 26927 38536 26939 38539
rect 27706 38536 27712 38548
rect 26927 38508 27712 38536
rect 26927 38505 26939 38508
rect 26881 38499 26939 38505
rect 27706 38496 27712 38508
rect 27764 38536 27770 38548
rect 28442 38536 28448 38548
rect 27764 38508 28448 38536
rect 27764 38496 27770 38508
rect 28442 38496 28448 38508
rect 28500 38496 28506 38548
rect 28813 38539 28871 38545
rect 28813 38505 28825 38539
rect 28859 38505 28871 38539
rect 28813 38499 28871 38505
rect 6641 38471 6699 38477
rect 6641 38437 6653 38471
rect 6687 38468 6699 38471
rect 7282 38468 7288 38480
rect 6687 38440 7288 38468
rect 6687 38437 6699 38440
rect 6641 38431 6699 38437
rect 7282 38428 7288 38440
rect 7340 38428 7346 38480
rect 26697 38471 26755 38477
rect 26697 38437 26709 38471
rect 26743 38437 26755 38471
rect 26697 38431 26755 38437
rect 27249 38471 27307 38477
rect 27249 38437 27261 38471
rect 27295 38468 27307 38471
rect 27614 38468 27620 38480
rect 27295 38440 27620 38468
rect 27295 38437 27307 38440
rect 27249 38431 27307 38437
rect 5258 38400 5264 38412
rect 5219 38372 5264 38400
rect 5258 38360 5264 38372
rect 5316 38360 5322 38412
rect 13170 38400 13176 38412
rect 13131 38372 13176 38400
rect 13170 38360 13176 38372
rect 13228 38360 13234 38412
rect 5534 38341 5540 38344
rect 5528 38332 5540 38341
rect 5495 38304 5540 38332
rect 5528 38295 5540 38304
rect 5534 38292 5540 38295
rect 5592 38292 5598 38344
rect 8225 38335 8283 38341
rect 8225 38301 8237 38335
rect 8271 38332 8283 38335
rect 8386 38332 8392 38344
rect 8271 38304 8392 38332
rect 8271 38301 8283 38304
rect 8225 38295 8283 38301
rect 8386 38292 8392 38304
rect 8444 38292 8450 38344
rect 8481 38335 8539 38341
rect 8481 38301 8493 38335
rect 8527 38332 8539 38335
rect 8754 38332 8760 38344
rect 8527 38304 8760 38332
rect 8527 38301 8539 38304
rect 8481 38295 8539 38301
rect 8754 38292 8760 38304
rect 8812 38332 8818 38344
rect 9766 38332 9772 38344
rect 8812 38304 9772 38332
rect 8812 38292 8818 38304
rect 9766 38292 9772 38304
rect 9824 38292 9830 38344
rect 10594 38332 10600 38344
rect 10555 38304 10600 38332
rect 10594 38292 10600 38304
rect 10652 38292 10658 38344
rect 11241 38335 11299 38341
rect 11241 38301 11253 38335
rect 11287 38332 11299 38335
rect 11790 38332 11796 38344
rect 11287 38304 11796 38332
rect 11287 38301 11299 38304
rect 11241 38295 11299 38301
rect 11790 38292 11796 38304
rect 11848 38332 11854 38344
rect 12526 38332 12532 38344
rect 11848 38304 12532 38332
rect 11848 38292 11854 38304
rect 12526 38292 12532 38304
rect 12584 38292 12590 38344
rect 13357 38335 13415 38341
rect 13357 38301 13369 38335
rect 13403 38332 13415 38335
rect 13906 38332 13912 38344
rect 13403 38304 13912 38332
rect 13403 38301 13415 38304
rect 13357 38295 13415 38301
rect 13906 38292 13912 38304
rect 13964 38292 13970 38344
rect 23566 38332 23572 38344
rect 23527 38304 23572 38332
rect 23566 38292 23572 38304
rect 23624 38292 23630 38344
rect 26053 38335 26111 38341
rect 26053 38301 26065 38335
rect 26099 38332 26111 38335
rect 26712 38332 26740 38431
rect 27614 38428 27620 38440
rect 27672 38468 27678 38480
rect 28629 38471 28687 38477
rect 28629 38468 28641 38471
rect 27672 38440 28641 38468
rect 27672 38428 27678 38440
rect 28629 38437 28641 38440
rect 28675 38437 28687 38471
rect 28629 38431 28687 38437
rect 28828 38400 28856 38499
rect 28902 38496 28908 38548
rect 28960 38536 28966 38548
rect 30009 38539 30067 38545
rect 30009 38536 30021 38539
rect 28960 38508 30021 38536
rect 28960 38496 28966 38508
rect 30009 38505 30021 38508
rect 30055 38536 30067 38539
rect 30929 38539 30987 38545
rect 30929 38536 30941 38539
rect 30055 38508 30941 38536
rect 30055 38505 30067 38508
rect 30009 38499 30067 38505
rect 30929 38505 30941 38508
rect 30975 38505 30987 38539
rect 39206 38536 39212 38548
rect 39167 38508 39212 38536
rect 30929 38499 30987 38505
rect 39206 38496 39212 38508
rect 39264 38536 39270 38548
rect 42613 38539 42671 38545
rect 42613 38536 42625 38539
rect 39264 38508 42625 38536
rect 39264 38496 39270 38508
rect 42613 38505 42625 38508
rect 42659 38536 42671 38539
rect 42794 38536 42800 38548
rect 42659 38508 42800 38536
rect 42659 38505 42671 38508
rect 42613 38499 42671 38505
rect 42794 38496 42800 38508
rect 42852 38496 42858 38548
rect 43441 38539 43499 38545
rect 43441 38505 43453 38539
rect 43487 38536 43499 38539
rect 44450 38536 44456 38548
rect 43487 38508 44456 38536
rect 43487 38505 43499 38508
rect 43441 38499 43499 38505
rect 44450 38496 44456 38508
rect 44508 38496 44514 38548
rect 30193 38471 30251 38477
rect 30193 38437 30205 38471
rect 30239 38468 30251 38471
rect 31754 38468 31760 38480
rect 30239 38440 31760 38468
rect 30239 38437 30251 38440
rect 30193 38431 30251 38437
rect 31754 38428 31760 38440
rect 31812 38428 31818 38480
rect 27908 38372 28856 38400
rect 26099 38304 26740 38332
rect 26099 38301 26111 38304
rect 26053 38295 26111 38301
rect 27430 38292 27436 38344
rect 27488 38332 27494 38344
rect 27908 38341 27936 38372
rect 27893 38335 27951 38341
rect 27893 38332 27905 38335
rect 27488 38304 27905 38332
rect 27488 38292 27494 38304
rect 27893 38301 27905 38304
rect 27939 38301 27951 38335
rect 27893 38295 27951 38301
rect 28169 38335 28227 38341
rect 28169 38301 28181 38335
rect 28215 38332 28227 38335
rect 28350 38332 28356 38344
rect 28215 38304 28356 38332
rect 28215 38301 28227 38304
rect 28169 38295 28227 38301
rect 28350 38292 28356 38304
rect 28408 38292 28414 38344
rect 31665 38335 31723 38341
rect 31665 38332 31677 38335
rect 31128 38304 31677 38332
rect 11508 38267 11566 38273
rect 11508 38233 11520 38267
rect 11554 38264 11566 38267
rect 11698 38264 11704 38276
rect 11554 38236 11704 38264
rect 11554 38233 11566 38236
rect 11508 38227 11566 38233
rect 11698 38224 11704 38236
rect 11756 38224 11762 38276
rect 13078 38264 13084 38276
rect 13039 38236 13084 38264
rect 13078 38224 13084 38236
rect 13136 38224 13142 38276
rect 28997 38267 29055 38273
rect 28997 38264 29009 38267
rect 28184 38236 29009 38264
rect 28184 38208 28212 38236
rect 28997 38233 29009 38236
rect 29043 38233 29055 38267
rect 28997 38227 29055 38233
rect 29638 38224 29644 38276
rect 29696 38264 29702 38276
rect 29825 38267 29883 38273
rect 29825 38264 29837 38267
rect 29696 38236 29837 38264
rect 29696 38224 29702 38236
rect 29825 38233 29837 38236
rect 29871 38233 29883 38267
rect 30742 38264 30748 38276
rect 30703 38236 30748 38264
rect 29825 38227 29883 38233
rect 30742 38224 30748 38236
rect 30800 38224 30806 38276
rect 26234 38196 26240 38208
rect 26195 38168 26240 38196
rect 26234 38156 26240 38168
rect 26292 38156 26298 38208
rect 26881 38199 26939 38205
rect 26881 38165 26893 38199
rect 26927 38196 26939 38199
rect 27709 38199 27767 38205
rect 27709 38196 27721 38199
rect 26927 38168 27721 38196
rect 26927 38165 26939 38168
rect 26881 38159 26939 38165
rect 27709 38165 27721 38168
rect 27755 38165 27767 38199
rect 27709 38159 27767 38165
rect 28077 38199 28135 38205
rect 28077 38165 28089 38199
rect 28123 38196 28135 38199
rect 28166 38196 28172 38208
rect 28123 38168 28172 38196
rect 28123 38165 28135 38168
rect 28077 38159 28135 38165
rect 28166 38156 28172 38168
rect 28224 38156 28230 38208
rect 28350 38156 28356 38208
rect 28408 38196 28414 38208
rect 28787 38199 28845 38205
rect 28787 38196 28799 38199
rect 28408 38168 28799 38196
rect 28408 38156 28414 38168
rect 28787 38165 28799 38168
rect 28833 38165 28845 38199
rect 28787 38159 28845 38165
rect 30006 38156 30012 38208
rect 30064 38205 30070 38208
rect 30064 38199 30083 38205
rect 30071 38165 30083 38199
rect 30064 38159 30083 38165
rect 30064 38156 30070 38159
rect 30926 38156 30932 38208
rect 30984 38205 30990 38208
rect 31128 38205 31156 38304
rect 31665 38301 31677 38304
rect 31711 38301 31723 38335
rect 31665 38295 31723 38301
rect 36081 38335 36139 38341
rect 36081 38301 36093 38335
rect 36127 38301 36139 38335
rect 36081 38295 36139 38301
rect 36541 38335 36599 38341
rect 36541 38301 36553 38335
rect 36587 38332 36599 38335
rect 37274 38332 37280 38344
rect 36587 38304 37280 38332
rect 36587 38301 36599 38304
rect 36541 38295 36599 38301
rect 36096 38264 36124 38295
rect 37274 38292 37280 38304
rect 37332 38292 37338 38344
rect 40037 38335 40095 38341
rect 40037 38301 40049 38335
rect 40083 38332 40095 38335
rect 40126 38332 40132 38344
rect 40083 38304 40132 38332
rect 40083 38301 40095 38304
rect 40037 38295 40095 38301
rect 40126 38292 40132 38304
rect 40184 38292 40190 38344
rect 40678 38332 40684 38344
rect 40639 38304 40684 38332
rect 40678 38292 40684 38304
rect 40736 38292 40742 38344
rect 42058 38292 42064 38344
rect 42116 38332 42122 38344
rect 43257 38335 43315 38341
rect 43257 38332 43269 38335
rect 42116 38304 43269 38332
rect 42116 38292 42122 38304
rect 43257 38301 43269 38304
rect 43303 38301 43315 38335
rect 43257 38295 43315 38301
rect 36786 38267 36844 38273
rect 36786 38264 36798 38267
rect 36096 38236 36798 38264
rect 36786 38233 36798 38236
rect 36832 38233 36844 38267
rect 36786 38227 36844 38233
rect 40948 38267 41006 38273
rect 40948 38233 40960 38267
rect 40994 38264 41006 38267
rect 42702 38264 42708 38276
rect 40994 38236 42708 38264
rect 40994 38233 41006 38236
rect 40948 38227 41006 38233
rect 42702 38224 42708 38236
rect 42760 38224 42766 38276
rect 30984 38199 31003 38205
rect 30991 38165 31003 38199
rect 30984 38159 31003 38165
rect 31113 38199 31171 38205
rect 31113 38165 31125 38199
rect 31159 38165 31171 38199
rect 31846 38196 31852 38208
rect 31807 38168 31852 38196
rect 31113 38159 31171 38165
rect 30984 38156 30990 38159
rect 31846 38156 31852 38168
rect 31904 38156 31910 38208
rect 37921 38199 37979 38205
rect 37921 38165 37933 38199
rect 37967 38196 37979 38199
rect 38286 38196 38292 38208
rect 37967 38168 38292 38196
rect 37967 38165 37979 38168
rect 37921 38159 37979 38165
rect 38286 38156 38292 38168
rect 38344 38156 38350 38208
rect 40221 38199 40279 38205
rect 40221 38165 40233 38199
rect 40267 38196 40279 38199
rect 40310 38196 40316 38208
rect 40267 38168 40316 38196
rect 40267 38165 40279 38168
rect 40221 38159 40279 38165
rect 40310 38156 40316 38168
rect 40368 38156 40374 38208
rect 41598 38156 41604 38208
rect 41656 38196 41662 38208
rect 42061 38199 42119 38205
rect 42061 38196 42073 38199
rect 41656 38168 42073 38196
rect 41656 38156 41662 38168
rect 42061 38165 42073 38168
rect 42107 38165 42119 38199
rect 42061 38159 42119 38165
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 6914 37952 6920 38004
rect 6972 37952 6978 38004
rect 7374 37952 7380 38004
rect 7432 37992 7438 38004
rect 8113 37995 8171 38001
rect 8113 37992 8125 37995
rect 7432 37964 8125 37992
rect 7432 37952 7438 37964
rect 8113 37961 8125 37964
rect 8159 37961 8171 37995
rect 8113 37955 8171 37961
rect 11149 37995 11207 38001
rect 11149 37961 11161 37995
rect 11195 37992 11207 37995
rect 13078 37992 13084 38004
rect 11195 37964 13084 37992
rect 11195 37961 11207 37964
rect 11149 37955 11207 37961
rect 13078 37952 13084 37964
rect 13136 37952 13142 38004
rect 13906 37992 13912 38004
rect 13867 37964 13912 37992
rect 13906 37952 13912 37964
rect 13964 37952 13970 38004
rect 27325 37995 27383 38001
rect 27325 37961 27337 37995
rect 27371 37992 27383 37995
rect 27985 37995 28043 38001
rect 27985 37992 27997 37995
rect 27371 37964 27997 37992
rect 27371 37961 27383 37964
rect 27325 37955 27383 37961
rect 27985 37961 27997 37964
rect 28031 37961 28043 37995
rect 30285 37995 30343 38001
rect 30285 37992 30297 37995
rect 27985 37955 28043 37961
rect 29472 37964 30297 37992
rect 6932 37924 6960 37952
rect 8754 37924 8760 37936
rect 6886 37896 8760 37924
rect 6733 37859 6791 37865
rect 6733 37825 6745 37859
rect 6779 37856 6791 37859
rect 6886 37856 6914 37896
rect 8754 37884 8760 37896
rect 8812 37884 8818 37936
rect 10036 37927 10094 37933
rect 10036 37893 10048 37927
rect 10082 37924 10094 37927
rect 10594 37924 10600 37936
rect 10082 37896 10600 37924
rect 10082 37893 10094 37896
rect 10036 37887 10094 37893
rect 10594 37884 10600 37896
rect 10652 37884 10658 37936
rect 23566 37933 23572 37936
rect 12774 37927 12832 37933
rect 12774 37924 12786 37927
rect 12084 37896 12786 37924
rect 7006 37865 7012 37868
rect 6779 37828 6914 37856
rect 6779 37825 6791 37828
rect 6733 37819 6791 37825
rect 7000 37819 7012 37865
rect 7064 37856 7070 37868
rect 12084 37865 12112 37896
rect 12774 37893 12786 37896
rect 12820 37893 12832 37927
rect 23560 37924 23572 37933
rect 23527 37896 23572 37924
rect 12774 37887 12832 37893
rect 23560 37887 23572 37896
rect 23566 37884 23572 37887
rect 23624 37884 23630 37936
rect 27522 37924 27528 37936
rect 27483 37896 27528 37924
rect 27522 37884 27528 37896
rect 27580 37884 27586 37936
rect 29365 37927 29423 37933
rect 29365 37893 29377 37927
rect 29411 37924 29423 37927
rect 29472 37924 29500 37964
rect 30285 37961 30297 37964
rect 30331 37992 30343 37995
rect 30558 37992 30564 38004
rect 30331 37964 30564 37992
rect 30331 37961 30343 37964
rect 30285 37955 30343 37961
rect 30558 37952 30564 37964
rect 30616 37952 30622 38004
rect 30926 37952 30932 38004
rect 30984 37992 30990 38004
rect 31113 37995 31171 38001
rect 31113 37992 31125 37995
rect 30984 37964 31125 37992
rect 30984 37952 30990 37964
rect 31113 37961 31125 37964
rect 31159 37961 31171 37995
rect 42058 37992 42064 38004
rect 42019 37964 42064 37992
rect 31113 37955 31171 37961
rect 42058 37952 42064 37964
rect 42116 37952 42122 38004
rect 29411 37896 29500 37924
rect 29549 37927 29607 37933
rect 29411 37893 29423 37896
rect 29365 37887 29423 37893
rect 29549 37893 29561 37927
rect 29595 37924 29607 37927
rect 30834 37924 30840 37936
rect 29595 37896 30144 37924
rect 29595 37893 29607 37896
rect 29549 37887 29607 37893
rect 12069 37859 12127 37865
rect 7064 37828 7100 37856
rect 7006 37816 7012 37819
rect 7064 37816 7070 37828
rect 12069 37825 12081 37859
rect 12115 37825 12127 37859
rect 12526 37856 12532 37868
rect 12487 37828 12532 37856
rect 12069 37819 12127 37825
rect 12526 37816 12532 37828
rect 12584 37816 12590 37868
rect 23290 37856 23296 37868
rect 23251 37828 23296 37856
rect 23290 37816 23296 37828
rect 23348 37816 23354 37868
rect 28166 37856 28172 37868
rect 28127 37828 28172 37856
rect 28166 37816 28172 37828
rect 28224 37816 28230 37868
rect 28350 37856 28356 37868
rect 28311 37828 28356 37856
rect 28350 37816 28356 37828
rect 28408 37816 28414 37868
rect 29641 37862 29699 37865
rect 29641 37859 29776 37862
rect 29641 37825 29653 37859
rect 29687 37856 29776 37859
rect 30116 37856 30144 37896
rect 30392 37896 30840 37924
rect 30392 37868 30420 37896
rect 30834 37884 30840 37896
rect 30892 37924 30898 37936
rect 31297 37927 31355 37933
rect 31297 37924 31309 37927
rect 30892 37896 31309 37924
rect 30892 37884 30898 37896
rect 31297 37893 31309 37896
rect 31343 37924 31355 37927
rect 31343 37896 31754 37924
rect 31343 37893 31355 37896
rect 31297 37887 31355 37893
rect 30374 37856 30380 37868
rect 29687 37834 30052 37856
rect 29687 37825 29699 37834
rect 29748 37828 30052 37834
rect 30116 37828 30380 37856
rect 29641 37819 29699 37825
rect 9766 37788 9772 37800
rect 9727 37760 9772 37788
rect 9766 37748 9772 37760
rect 9824 37748 9830 37800
rect 30024 37788 30052 37828
rect 30374 37816 30380 37828
rect 30432 37816 30438 37868
rect 30469 37859 30527 37865
rect 30469 37825 30481 37859
rect 30515 37856 30527 37859
rect 31110 37856 31116 37868
rect 30515 37828 31116 37856
rect 30515 37825 30527 37828
rect 30469 37819 30527 37825
rect 31110 37816 31116 37828
rect 31168 37816 31174 37868
rect 31478 37856 31484 37868
rect 31439 37828 31484 37856
rect 31478 37816 31484 37828
rect 31536 37816 31542 37868
rect 30024 37760 30328 37788
rect 30300 37732 30328 37760
rect 28350 37680 28356 37732
rect 28408 37720 28414 37732
rect 30101 37723 30159 37729
rect 30101 37720 30113 37723
rect 28408 37692 30113 37720
rect 28408 37680 28414 37692
rect 30101 37689 30113 37692
rect 30147 37689 30159 37723
rect 30101 37683 30159 37689
rect 30282 37680 30288 37732
rect 30340 37720 30346 37732
rect 30653 37723 30711 37729
rect 30653 37720 30665 37723
rect 30340 37692 30665 37720
rect 30340 37680 30346 37692
rect 30653 37689 30665 37692
rect 30699 37689 30711 37723
rect 30653 37683 30711 37689
rect 5810 37652 5816 37664
rect 5771 37624 5816 37652
rect 5810 37612 5816 37624
rect 5868 37612 5874 37664
rect 24670 37652 24676 37664
rect 24631 37624 24676 37652
rect 24670 37612 24676 37624
rect 24728 37612 24734 37664
rect 27062 37612 27068 37664
rect 27120 37652 27126 37664
rect 27157 37655 27215 37661
rect 27157 37652 27169 37655
rect 27120 37624 27169 37652
rect 27120 37612 27126 37624
rect 27157 37621 27169 37624
rect 27203 37621 27215 37655
rect 27157 37615 27215 37621
rect 27341 37655 27399 37661
rect 27341 37621 27353 37655
rect 27387 37652 27399 37655
rect 27706 37652 27712 37664
rect 27387 37624 27712 37652
rect 27387 37621 27399 37624
rect 27341 37615 27399 37621
rect 27706 37612 27712 37624
rect 27764 37652 27770 37664
rect 28810 37652 28816 37664
rect 27764 37624 28816 37652
rect 27764 37612 27770 37624
rect 28810 37612 28816 37624
rect 28868 37612 28874 37664
rect 29638 37652 29644 37664
rect 29599 37624 29644 37652
rect 29638 37612 29644 37624
rect 29696 37612 29702 37664
rect 31726 37652 31754 37896
rect 31846 37884 31852 37936
rect 31904 37924 31910 37936
rect 32554 37927 32612 37933
rect 32554 37924 32566 37927
rect 31904 37896 32566 37924
rect 31904 37884 31910 37896
rect 32554 37893 32566 37896
rect 32600 37893 32612 37927
rect 32554 37887 32612 37893
rect 39206 37884 39212 37936
rect 39264 37924 39270 37936
rect 39390 37924 39396 37936
rect 39264 37896 39396 37924
rect 39264 37884 39270 37896
rect 39390 37884 39396 37896
rect 39448 37884 39454 37936
rect 42794 37924 42800 37936
rect 42755 37896 42800 37924
rect 42794 37884 42800 37896
rect 42852 37884 42858 37936
rect 44542 37924 44548 37936
rect 44503 37896 44548 37924
rect 44542 37884 44548 37896
rect 44600 37884 44606 37936
rect 36630 37816 36636 37868
rect 36688 37865 36694 37868
rect 36688 37856 36700 37865
rect 36909 37859 36967 37865
rect 36688 37828 36733 37856
rect 36688 37819 36700 37828
rect 36909 37825 36921 37859
rect 36955 37856 36967 37859
rect 37274 37856 37280 37868
rect 36955 37828 37280 37856
rect 36955 37825 36967 37828
rect 36909 37819 36967 37825
rect 36688 37816 36694 37819
rect 37274 37816 37280 37828
rect 37332 37816 37338 37868
rect 37734 37865 37740 37868
rect 37728 37819 37740 37865
rect 37792 37856 37798 37868
rect 37792 37828 37828 37856
rect 37734 37816 37740 37819
rect 37792 37816 37798 37828
rect 32306 37788 32312 37800
rect 32267 37760 32312 37788
rect 32306 37748 32312 37760
rect 32364 37748 32370 37800
rect 37458 37788 37464 37800
rect 37419 37760 37464 37788
rect 37458 37748 37464 37760
rect 37516 37748 37522 37800
rect 41598 37788 41604 37800
rect 41559 37760 41604 37788
rect 41598 37748 41604 37760
rect 41656 37748 41662 37800
rect 41874 37720 41880 37732
rect 41835 37692 41880 37720
rect 41874 37680 41880 37692
rect 41932 37680 41938 37732
rect 31846 37652 31852 37664
rect 31726 37624 31852 37652
rect 31846 37612 31852 37624
rect 31904 37652 31910 37664
rect 33689 37655 33747 37661
rect 33689 37652 33701 37655
rect 31904 37624 33701 37652
rect 31904 37612 31910 37624
rect 33689 37621 33701 37624
rect 33735 37621 33747 37655
rect 33689 37615 33747 37621
rect 35529 37655 35587 37661
rect 35529 37621 35541 37655
rect 35575 37652 35587 37655
rect 38194 37652 38200 37664
rect 35575 37624 38200 37652
rect 35575 37621 35587 37624
rect 35529 37615 35587 37621
rect 38194 37612 38200 37624
rect 38252 37612 38258 37664
rect 38838 37652 38844 37664
rect 38799 37624 38844 37652
rect 38838 37612 38844 37624
rect 38896 37612 38902 37664
rect 40034 37612 40040 37664
rect 40092 37652 40098 37664
rect 40678 37652 40684 37664
rect 40092 37624 40684 37652
rect 40092 37612 40098 37624
rect 40678 37612 40684 37624
rect 40736 37612 40742 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 12989 37451 13047 37457
rect 12989 37417 13001 37451
rect 13035 37448 13047 37451
rect 13170 37448 13176 37460
rect 13035 37420 13176 37448
rect 13035 37417 13047 37420
rect 12989 37411 13047 37417
rect 13170 37408 13176 37420
rect 13228 37408 13234 37460
rect 24578 37448 24584 37460
rect 24539 37420 24584 37448
rect 24578 37408 24584 37420
rect 24636 37408 24642 37460
rect 27430 37448 27436 37460
rect 27391 37420 27436 37448
rect 27430 37408 27436 37420
rect 27488 37408 27494 37460
rect 28350 37408 28356 37460
rect 28408 37448 28414 37460
rect 28408 37420 28764 37448
rect 28408 37408 28414 37420
rect 28629 37383 28687 37389
rect 28629 37349 28641 37383
rect 28675 37349 28687 37383
rect 28736 37380 28764 37420
rect 28810 37408 28816 37460
rect 28868 37448 28874 37460
rect 28868 37420 28913 37448
rect 28868 37408 28874 37420
rect 30650 37408 30656 37460
rect 30708 37408 30714 37460
rect 31110 37448 31116 37460
rect 31071 37420 31116 37448
rect 31110 37408 31116 37420
rect 31168 37448 31174 37460
rect 38194 37448 38200 37460
rect 31168 37420 32076 37448
rect 38155 37420 38200 37448
rect 31168 37408 31174 37420
rect 29181 37383 29239 37389
rect 29181 37380 29193 37383
rect 28736 37352 29193 37380
rect 28629 37343 28687 37349
rect 29181 37349 29193 37352
rect 29227 37349 29239 37383
rect 30668 37380 30696 37408
rect 31478 37380 31484 37392
rect 30668 37352 31484 37380
rect 29181 37343 29239 37349
rect 5258 37272 5264 37324
rect 5316 37312 5322 37324
rect 5537 37315 5595 37321
rect 5537 37312 5549 37315
rect 5316 37284 5549 37312
rect 5316 37272 5322 37284
rect 5537 37281 5549 37284
rect 5583 37281 5595 37315
rect 24670 37312 24676 37324
rect 24631 37284 24676 37312
rect 5537 37275 5595 37281
rect 24670 37272 24676 37284
rect 24728 37272 24734 37324
rect 5810 37253 5816 37256
rect 5804 37244 5816 37253
rect 5771 37216 5816 37244
rect 5804 37207 5816 37216
rect 5810 37204 5816 37207
rect 5868 37204 5874 37256
rect 9766 37204 9772 37256
rect 9824 37244 9830 37256
rect 11609 37247 11667 37253
rect 11609 37244 11621 37247
rect 9824 37216 11621 37244
rect 9824 37204 9830 37216
rect 11609 37213 11621 37216
rect 11655 37213 11667 37247
rect 11609 37207 11667 37213
rect 22649 37247 22707 37253
rect 22649 37213 22661 37247
rect 22695 37244 22707 37247
rect 23290 37244 23296 37256
rect 22695 37216 23296 37244
rect 22695 37213 22707 37216
rect 22649 37207 22707 37213
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 24854 37244 24860 37256
rect 24815 37216 24860 37244
rect 24854 37204 24860 37216
rect 24912 37204 24918 37256
rect 26053 37247 26111 37253
rect 26053 37213 26065 37247
rect 26099 37213 26111 37247
rect 26053 37207 26111 37213
rect 26320 37247 26378 37253
rect 26320 37213 26332 37247
rect 26366 37213 26378 37247
rect 26320 37207 26378 37213
rect 27985 37247 28043 37253
rect 27985 37213 27997 37247
rect 28031 37244 28043 37247
rect 28644 37244 28672 37343
rect 31478 37340 31484 37352
rect 31536 37380 31542 37392
rect 31536 37352 31800 37380
rect 31536 37340 31542 37352
rect 29564 37284 29868 37312
rect 29564 37244 29592 37284
rect 29730 37244 29736 37256
rect 28031 37216 28672 37244
rect 28736 37216 29592 37244
rect 29643 37216 29736 37244
rect 28031 37213 28043 37216
rect 27985 37207 28043 37213
rect 11882 37185 11888 37188
rect 11876 37139 11888 37185
rect 11940 37176 11946 37188
rect 22922 37185 22928 37188
rect 11940 37148 11976 37176
rect 11882 37136 11888 37139
rect 11940 37136 11946 37148
rect 22916 37139 22928 37185
rect 22980 37176 22986 37188
rect 24581 37179 24639 37185
rect 22980 37148 23016 37176
rect 22922 37136 22928 37139
rect 22980 37136 22986 37148
rect 24581 37145 24593 37179
rect 24627 37145 24639 37179
rect 24581 37139 24639 37145
rect 6917 37111 6975 37117
rect 6917 37077 6929 37111
rect 6963 37108 6975 37111
rect 7190 37108 7196 37120
rect 6963 37080 7196 37108
rect 6963 37077 6975 37080
rect 6917 37071 6975 37077
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 24029 37111 24087 37117
rect 24029 37077 24041 37111
rect 24075 37108 24087 37111
rect 24596 37108 24624 37139
rect 24075 37080 24624 37108
rect 25041 37111 25099 37117
rect 24075 37077 24087 37080
rect 24029 37071 24087 37077
rect 25041 37077 25053 37111
rect 25087 37108 25099 37111
rect 25590 37108 25596 37120
rect 25087 37080 25596 37108
rect 25087 37077 25099 37080
rect 25041 37071 25099 37077
rect 25590 37068 25596 37080
rect 25648 37068 25654 37120
rect 26068 37108 26096 37207
rect 26234 37136 26240 37188
rect 26292 37176 26298 37188
rect 26344 37176 26372 37207
rect 27798 37176 27804 37188
rect 26292 37148 26372 37176
rect 27172 37148 27804 37176
rect 26292 37136 26298 37148
rect 27172 37120 27200 37148
rect 27798 37136 27804 37148
rect 27856 37176 27862 37188
rect 28626 37176 28632 37188
rect 27856 37148 28632 37176
rect 27856 37136 27862 37148
rect 28626 37136 28632 37148
rect 28684 37136 28690 37188
rect 27154 37108 27160 37120
rect 26068 37080 27160 37108
rect 27154 37068 27160 37080
rect 27212 37068 27218 37120
rect 28169 37111 28227 37117
rect 28169 37077 28181 37111
rect 28215 37108 28227 37111
rect 28736 37108 28764 37216
rect 28902 37136 28908 37188
rect 28960 37176 28966 37188
rect 29656 37176 29684 37216
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 29840 37244 29868 37284
rect 29989 37247 30047 37253
rect 29989 37244 30001 37247
rect 29840 37216 30001 37244
rect 29989 37213 30001 37216
rect 30035 37213 30047 37247
rect 29989 37207 30047 37213
rect 30282 37204 30288 37256
rect 30340 37244 30346 37256
rect 31772 37253 31800 37352
rect 31846 37272 31852 37324
rect 31904 37312 31910 37324
rect 31904 37284 31949 37312
rect 31904 37272 31910 37284
rect 32048 37253 32076 37420
rect 38194 37408 38200 37420
rect 38252 37408 38258 37460
rect 39393 37451 39451 37457
rect 39393 37417 39405 37451
rect 39439 37448 39451 37451
rect 40218 37448 40224 37460
rect 39439 37420 40224 37448
rect 39439 37417 39451 37420
rect 39393 37411 39451 37417
rect 40218 37408 40224 37420
rect 40276 37448 40282 37460
rect 42061 37451 42119 37457
rect 42061 37448 42073 37451
rect 40276 37420 42073 37448
rect 40276 37408 40282 37420
rect 42061 37417 42073 37420
rect 42107 37417 42119 37451
rect 42702 37448 42708 37460
rect 42663 37420 42708 37448
rect 42061 37411 42119 37417
rect 42702 37408 42708 37420
rect 42760 37408 42766 37460
rect 38286 37312 38292 37324
rect 38247 37284 38292 37312
rect 38286 37272 38292 37284
rect 38344 37272 38350 37324
rect 40034 37312 40040 37324
rect 38396 37284 40040 37312
rect 31757 37247 31815 37253
rect 30340 37216 31708 37244
rect 30340 37204 30346 37216
rect 28960 37148 29684 37176
rect 31680 37176 31708 37216
rect 31757 37213 31769 37247
rect 31803 37213 31815 37247
rect 31757 37207 31815 37213
rect 31941 37247 31999 37253
rect 31941 37213 31953 37247
rect 31987 37213 31999 37247
rect 31941 37207 31999 37213
rect 32033 37247 32091 37253
rect 32033 37213 32045 37247
rect 32079 37213 32091 37247
rect 32033 37207 32091 37213
rect 31956 37176 31984 37207
rect 36170 37204 36176 37256
rect 36228 37244 36234 37256
rect 36357 37247 36415 37253
rect 36357 37244 36369 37247
rect 36228 37216 36369 37244
rect 36228 37204 36234 37216
rect 36357 37213 36369 37216
rect 36403 37244 36415 37247
rect 37458 37244 37464 37256
rect 36403 37216 37464 37244
rect 36403 37213 36415 37216
rect 36357 37207 36415 37213
rect 37458 37204 37464 37216
rect 37516 37244 37522 37256
rect 38396 37244 38424 37284
rect 40034 37272 40040 37284
rect 40092 37272 40098 37324
rect 37516 37216 38424 37244
rect 38473 37247 38531 37253
rect 37516 37204 37522 37216
rect 38473 37213 38485 37247
rect 38519 37244 38531 37247
rect 38838 37244 38844 37256
rect 38519 37216 38844 37244
rect 38519 37213 38531 37216
rect 38473 37207 38531 37213
rect 38838 37204 38844 37216
rect 38896 37204 38902 37256
rect 39298 37244 39304 37256
rect 39259 37216 39304 37244
rect 39298 37204 39304 37216
rect 39356 37204 39362 37256
rect 40310 37253 40316 37256
rect 39485 37247 39543 37253
rect 39485 37213 39497 37247
rect 39531 37213 39543 37247
rect 40304 37244 40316 37253
rect 40271 37216 40316 37244
rect 39485 37207 39543 37213
rect 40304 37207 40316 37216
rect 36630 37185 36636 37188
rect 31680 37148 31984 37176
rect 28960 37136 28966 37148
rect 36624 37139 36636 37185
rect 36688 37176 36694 37188
rect 38197 37179 38255 37185
rect 36688 37148 36724 37176
rect 36630 37136 36636 37139
rect 36688 37136 36694 37148
rect 38197 37145 38209 37179
rect 38243 37145 38255 37179
rect 39500 37176 39528 37207
rect 40310 37204 40316 37207
rect 40368 37204 40374 37256
rect 42889 37247 42947 37253
rect 42889 37244 42901 37247
rect 42260 37216 42901 37244
rect 41598 37176 41604 37188
rect 39500 37148 41604 37176
rect 38197 37139 38255 37145
rect 28215 37080 28764 37108
rect 28813 37111 28871 37117
rect 28215 37077 28227 37080
rect 28169 37071 28227 37077
rect 28813 37077 28825 37111
rect 28859 37108 28871 37111
rect 31573 37111 31631 37117
rect 31573 37108 31585 37111
rect 28859 37080 31585 37108
rect 28859 37077 28871 37080
rect 28813 37071 28871 37077
rect 31573 37077 31585 37080
rect 31619 37077 31631 37111
rect 31573 37071 31631 37077
rect 37737 37111 37795 37117
rect 37737 37077 37749 37111
rect 37783 37108 37795 37111
rect 38212 37108 38240 37139
rect 41598 37136 41604 37148
rect 41656 37136 41662 37188
rect 41874 37176 41880 37188
rect 41835 37148 41880 37176
rect 41874 37136 41880 37148
rect 41932 37136 41938 37188
rect 41966 37136 41972 37188
rect 42024 37176 42030 37188
rect 42077 37179 42135 37185
rect 42077 37176 42089 37179
rect 42024 37148 42089 37176
rect 42024 37136 42030 37148
rect 42077 37145 42089 37148
rect 42123 37145 42135 37179
rect 42077 37139 42135 37145
rect 38654 37108 38660 37120
rect 37783 37080 38240 37108
rect 38615 37080 38660 37108
rect 37783 37077 37795 37080
rect 37737 37071 37795 37077
rect 38654 37068 38660 37080
rect 38712 37068 38718 37120
rect 41414 37108 41420 37120
rect 41375 37080 41420 37108
rect 41414 37068 41420 37080
rect 41472 37068 41478 37120
rect 42260 37117 42288 37216
rect 42889 37213 42901 37216
rect 42935 37213 42947 37247
rect 42889 37207 42947 37213
rect 42245 37111 42303 37117
rect 42245 37077 42257 37111
rect 42291 37077 42303 37111
rect 42245 37071 42303 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 24854 36904 24860 36916
rect 24815 36876 24860 36904
rect 24854 36864 24860 36876
rect 24912 36864 24918 36916
rect 26605 36907 26663 36913
rect 26605 36873 26617 36907
rect 26651 36904 26663 36907
rect 27522 36904 27528 36916
rect 26651 36876 27528 36904
rect 26651 36873 26663 36876
rect 26605 36867 26663 36873
rect 27522 36864 27528 36876
rect 27580 36864 27586 36916
rect 28537 36907 28595 36913
rect 28537 36873 28549 36907
rect 28583 36873 28595 36907
rect 28537 36867 28595 36873
rect 28166 36836 28172 36848
rect 26620 36808 28172 36836
rect 11882 36768 11888 36780
rect 11843 36740 11888 36768
rect 11882 36728 11888 36740
rect 11940 36728 11946 36780
rect 22833 36771 22891 36777
rect 22833 36737 22845 36771
rect 22879 36768 22891 36771
rect 22922 36768 22928 36780
rect 22879 36740 22928 36768
rect 22879 36737 22891 36740
rect 22833 36731 22891 36737
rect 22922 36728 22928 36740
rect 22980 36728 22986 36780
rect 23750 36777 23756 36780
rect 23744 36731 23756 36777
rect 23808 36768 23814 36780
rect 26620 36777 26648 36808
rect 28166 36796 28172 36808
rect 28224 36836 28230 36848
rect 28552 36836 28580 36867
rect 29730 36864 29736 36916
rect 29788 36904 29794 36916
rect 31110 36904 31116 36916
rect 29788 36876 31116 36904
rect 29788 36864 29794 36876
rect 31110 36864 31116 36876
rect 31168 36904 31174 36916
rect 31297 36907 31355 36913
rect 31297 36904 31309 36907
rect 31168 36876 31309 36904
rect 31168 36864 31174 36876
rect 31297 36873 31309 36876
rect 31343 36904 31355 36907
rect 32306 36904 32312 36916
rect 31343 36876 32312 36904
rect 31343 36873 31355 36876
rect 31297 36867 31355 36873
rect 32306 36864 32312 36876
rect 32364 36864 32370 36916
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 40126 36904 40132 36916
rect 32456 36876 32501 36904
rect 40087 36876 40132 36904
rect 32456 36864 32462 36876
rect 40126 36864 40132 36876
rect 40184 36864 40190 36916
rect 40310 36864 40316 36916
rect 40368 36904 40374 36916
rect 41874 36904 41880 36916
rect 40368 36876 41880 36904
rect 40368 36864 40374 36876
rect 41874 36864 41880 36876
rect 41932 36864 41938 36916
rect 28224 36808 28580 36836
rect 30009 36839 30067 36845
rect 28224 36796 28230 36808
rect 30009 36805 30021 36839
rect 30055 36836 30067 36839
rect 32416 36836 32444 36864
rect 30055 36808 32444 36836
rect 30055 36805 30067 36808
rect 30009 36799 30067 36805
rect 26421 36771 26479 36777
rect 23808 36740 23844 36768
rect 23750 36728 23756 36731
rect 23808 36728 23814 36740
rect 26421 36737 26433 36771
rect 26467 36737 26479 36771
rect 26421 36731 26479 36737
rect 26605 36771 26663 36777
rect 26605 36737 26617 36771
rect 26651 36737 26663 36771
rect 27154 36768 27160 36780
rect 27115 36740 27160 36768
rect 26605 36731 26663 36737
rect 23474 36700 23480 36712
rect 23435 36672 23480 36700
rect 23474 36660 23480 36672
rect 23532 36660 23538 36712
rect 26436 36564 26464 36731
rect 27154 36728 27160 36740
rect 27212 36728 27218 36780
rect 27246 36728 27252 36780
rect 27304 36768 27310 36780
rect 27413 36771 27471 36777
rect 27413 36768 27425 36771
rect 27304 36740 27425 36768
rect 27304 36728 27310 36740
rect 27413 36737 27425 36740
rect 27459 36737 27471 36771
rect 36630 36768 36636 36780
rect 36591 36740 36636 36768
rect 27413 36731 27471 36737
rect 36630 36728 36636 36740
rect 36688 36728 36694 36780
rect 37645 36771 37703 36777
rect 37645 36737 37657 36771
rect 37691 36768 37703 36771
rect 37734 36768 37740 36780
rect 37691 36740 37740 36768
rect 37691 36737 37703 36740
rect 37645 36731 37703 36737
rect 37734 36728 37740 36740
rect 37792 36728 37798 36780
rect 39482 36768 39488 36780
rect 39395 36740 39488 36768
rect 39482 36728 39488 36740
rect 39540 36768 39546 36780
rect 41141 36771 41199 36777
rect 41141 36768 41153 36771
rect 39540 36740 41153 36768
rect 39540 36728 39546 36740
rect 41141 36737 41153 36740
rect 41187 36737 41199 36771
rect 41141 36731 41199 36737
rect 41325 36771 41383 36777
rect 41325 36737 41337 36771
rect 41371 36768 41383 36771
rect 41414 36768 41420 36780
rect 41371 36740 41420 36768
rect 41371 36737 41383 36740
rect 41325 36731 41383 36737
rect 39669 36703 39727 36709
rect 39669 36669 39681 36703
rect 39715 36700 39727 36703
rect 41340 36700 41368 36731
rect 41414 36728 41420 36740
rect 41472 36728 41478 36780
rect 39715 36672 41368 36700
rect 39715 36669 39727 36672
rect 39669 36663 39727 36669
rect 39298 36632 39304 36644
rect 39211 36604 39304 36632
rect 39298 36592 39304 36604
rect 39356 36632 39362 36644
rect 40681 36635 40739 36641
rect 40681 36632 40693 36635
rect 39356 36604 40693 36632
rect 39356 36592 39362 36604
rect 40681 36601 40693 36604
rect 40727 36632 40739 36635
rect 40770 36632 40776 36644
rect 40727 36604 40776 36632
rect 40727 36601 40739 36604
rect 40681 36595 40739 36601
rect 40770 36592 40776 36604
rect 40828 36592 40834 36644
rect 28350 36564 28356 36576
rect 26436 36536 28356 36564
rect 28350 36524 28356 36536
rect 28408 36524 28414 36576
rect 33226 36524 33232 36576
rect 33284 36564 33290 36576
rect 33321 36567 33379 36573
rect 33321 36564 33333 36567
rect 33284 36536 33333 36564
rect 33284 36524 33290 36536
rect 33321 36533 33333 36536
rect 33367 36533 33379 36567
rect 33321 36527 33379 36533
rect 40313 36567 40371 36573
rect 40313 36533 40325 36567
rect 40359 36564 40371 36567
rect 41509 36567 41567 36573
rect 41509 36564 41521 36567
rect 40359 36536 41521 36564
rect 40359 36533 40371 36536
rect 40313 36527 40371 36533
rect 41509 36533 41521 36536
rect 41555 36533 41567 36567
rect 41509 36527 41567 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 23750 36360 23756 36372
rect 23711 36332 23756 36360
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 27246 36360 27252 36372
rect 27207 36332 27252 36360
rect 27246 36320 27252 36332
rect 27304 36320 27310 36372
rect 29733 36363 29791 36369
rect 29733 36329 29745 36363
rect 29779 36360 29791 36363
rect 30190 36360 30196 36372
rect 29779 36332 30196 36360
rect 29779 36329 29791 36332
rect 29733 36323 29791 36329
rect 30190 36320 30196 36332
rect 30248 36320 30254 36372
rect 40310 36360 40316 36372
rect 40271 36332 40316 36360
rect 40310 36320 40316 36332
rect 40368 36320 40374 36372
rect 31110 36224 31116 36236
rect 31071 36196 31116 36224
rect 31110 36184 31116 36196
rect 31168 36184 31174 36236
rect 32306 36184 32312 36236
rect 32364 36224 32370 36236
rect 32950 36224 32956 36236
rect 32364 36196 32956 36224
rect 32364 36184 32370 36196
rect 32950 36184 32956 36196
rect 33008 36184 33014 36236
rect 36170 36224 36176 36236
rect 36131 36196 36176 36224
rect 36170 36184 36176 36196
rect 36228 36184 36234 36236
rect 27062 36156 27068 36168
rect 27023 36128 27068 36156
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 31754 36156 31760 36168
rect 31715 36128 31760 36156
rect 31754 36116 31760 36128
rect 31812 36116 31818 36168
rect 33226 36165 33232 36168
rect 33220 36156 33232 36165
rect 33187 36128 33232 36156
rect 33220 36119 33232 36128
rect 33226 36116 33232 36119
rect 33284 36116 33290 36168
rect 40681 36159 40739 36165
rect 40681 36125 40693 36159
rect 40727 36156 40739 36159
rect 41138 36156 41144 36168
rect 40727 36128 41144 36156
rect 40727 36125 40739 36128
rect 40681 36119 40739 36125
rect 41138 36116 41144 36128
rect 41196 36116 41202 36168
rect 30868 36091 30926 36097
rect 30868 36057 30880 36091
rect 30914 36088 30926 36091
rect 36440 36091 36498 36097
rect 30914 36060 31616 36088
rect 30914 36057 30926 36060
rect 30868 36051 30926 36057
rect 31588 36029 31616 36060
rect 36440 36057 36452 36091
rect 36486 36088 36498 36091
rect 38102 36088 38108 36100
rect 36486 36060 38108 36088
rect 36486 36057 36498 36060
rect 36440 36051 36498 36057
rect 38102 36048 38108 36060
rect 38160 36048 38166 36100
rect 40218 36048 40224 36100
rect 40276 36088 40282 36100
rect 40313 36091 40371 36097
rect 40313 36088 40325 36091
rect 40276 36060 40325 36088
rect 40276 36048 40282 36060
rect 40313 36057 40325 36060
rect 40359 36057 40371 36091
rect 40313 36051 40371 36057
rect 31573 36023 31631 36029
rect 31573 35989 31585 36023
rect 31619 35989 31631 36023
rect 31573 35983 31631 35989
rect 34333 36023 34391 36029
rect 34333 35989 34345 36023
rect 34379 36020 34391 36023
rect 34790 36020 34796 36032
rect 34379 35992 34796 36020
rect 34379 35989 34391 35992
rect 34333 35983 34391 35989
rect 34790 35980 34796 35992
rect 34848 35980 34854 36032
rect 37553 36023 37611 36029
rect 37553 35989 37565 36023
rect 37599 36020 37611 36023
rect 37642 36020 37648 36032
rect 37599 35992 37648 36020
rect 37599 35989 37611 35992
rect 37553 35983 37611 35989
rect 37642 35980 37648 35992
rect 37700 35980 37706 36032
rect 40126 36020 40132 36032
rect 40087 35992 40132 36020
rect 40126 35980 40132 35992
rect 40184 35980 40190 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 25961 35819 26019 35825
rect 25961 35785 25973 35819
rect 26007 35816 26019 35819
rect 26326 35816 26332 35828
rect 26007 35788 26332 35816
rect 26007 35785 26019 35788
rect 25961 35779 26019 35785
rect 26326 35776 26332 35788
rect 26384 35776 26390 35828
rect 30006 35816 30012 35828
rect 29967 35788 30012 35816
rect 30006 35776 30012 35788
rect 30064 35776 30070 35828
rect 30374 35816 30380 35828
rect 30335 35788 30380 35816
rect 30374 35776 30380 35788
rect 30432 35776 30438 35828
rect 41138 35816 41144 35828
rect 41099 35788 41144 35816
rect 41138 35776 41144 35788
rect 41196 35776 41202 35828
rect 33290 35751 33348 35757
rect 33290 35748 33302 35751
rect 32600 35720 33302 35748
rect 23566 35640 23572 35692
rect 23624 35680 23630 35692
rect 25593 35683 25651 35689
rect 25593 35680 25605 35683
rect 23624 35652 25605 35680
rect 23624 35640 23630 35652
rect 25593 35649 25605 35652
rect 25639 35649 25651 35683
rect 25593 35643 25651 35649
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35680 25835 35683
rect 27062 35680 27068 35692
rect 25823 35652 27068 35680
rect 25823 35649 25835 35652
rect 25777 35643 25835 35649
rect 27062 35640 27068 35652
rect 27120 35640 27126 35692
rect 30190 35680 30196 35692
rect 30151 35652 30196 35680
rect 30190 35640 30196 35652
rect 30248 35640 30254 35692
rect 30469 35683 30527 35689
rect 30469 35649 30481 35683
rect 30515 35680 30527 35683
rect 30558 35680 30564 35692
rect 30515 35652 30564 35680
rect 30515 35649 30527 35652
rect 30469 35643 30527 35649
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 32600 35689 32628 35720
rect 33290 35717 33302 35720
rect 33336 35717 33348 35751
rect 33290 35711 33348 35717
rect 40028 35751 40086 35757
rect 40028 35717 40040 35751
rect 40074 35748 40086 35751
rect 40218 35748 40224 35760
rect 40074 35720 40224 35748
rect 40074 35717 40086 35720
rect 40028 35711 40086 35717
rect 40218 35708 40224 35720
rect 40276 35708 40282 35760
rect 32585 35683 32643 35689
rect 32585 35649 32597 35683
rect 32631 35649 32643 35683
rect 32585 35643 32643 35649
rect 32950 35640 32956 35692
rect 33008 35680 33014 35692
rect 33045 35683 33103 35689
rect 33045 35680 33057 35683
rect 33008 35652 33057 35680
rect 33008 35640 33014 35652
rect 33045 35649 33057 35652
rect 33091 35649 33103 35683
rect 33045 35643 33103 35649
rect 39761 35615 39819 35621
rect 39761 35581 39773 35615
rect 39807 35581 39819 35615
rect 39761 35575 39819 35581
rect 22002 35476 22008 35488
rect 21963 35448 22008 35476
rect 22002 35436 22008 35448
rect 22060 35436 22066 35488
rect 25590 35476 25596 35488
rect 25551 35448 25596 35476
rect 25590 35436 25596 35448
rect 25648 35436 25654 35488
rect 34422 35476 34428 35488
rect 34383 35448 34428 35476
rect 34422 35436 34428 35448
rect 34480 35436 34486 35488
rect 34514 35436 34520 35488
rect 34572 35476 34578 35488
rect 34885 35479 34943 35485
rect 34885 35476 34897 35479
rect 34572 35448 34897 35476
rect 34572 35436 34578 35448
rect 34885 35445 34897 35448
rect 34931 35445 34943 35479
rect 36538 35476 36544 35488
rect 36499 35448 36544 35476
rect 34885 35439 34943 35445
rect 36538 35436 36544 35448
rect 36596 35436 36602 35488
rect 39776 35476 39804 35575
rect 40034 35476 40040 35488
rect 39776 35448 40040 35476
rect 40034 35436 40040 35448
rect 40092 35476 40098 35488
rect 40494 35476 40500 35488
rect 40092 35448 40500 35476
rect 40092 35436 40098 35448
rect 40494 35436 40500 35448
rect 40552 35436 40558 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 20070 35232 20076 35284
rect 20128 35272 20134 35284
rect 23109 35275 23167 35281
rect 23109 35272 23121 35275
rect 20128 35244 23121 35272
rect 20128 35232 20134 35244
rect 23109 35241 23121 35244
rect 23155 35241 23167 35275
rect 23566 35272 23572 35284
rect 23527 35244 23572 35272
rect 23109 35235 23167 35241
rect 23566 35232 23572 35244
rect 23624 35232 23630 35284
rect 34790 35232 34796 35284
rect 34848 35272 34854 35284
rect 34885 35275 34943 35281
rect 34885 35272 34897 35275
rect 34848 35244 34897 35272
rect 34848 35232 34854 35244
rect 34885 35241 34897 35244
rect 34931 35241 34943 35275
rect 38102 35272 38108 35284
rect 38063 35244 38108 35272
rect 34885 35235 34943 35241
rect 38102 35232 38108 35244
rect 38160 35232 38166 35284
rect 40218 35272 40224 35284
rect 40179 35244 40224 35272
rect 40218 35232 40224 35244
rect 40276 35232 40282 35284
rect 34333 35207 34391 35213
rect 34333 35173 34345 35207
rect 34379 35204 34391 35207
rect 34379 35176 35020 35204
rect 34379 35173 34391 35176
rect 34333 35167 34391 35173
rect 23474 35096 23480 35148
rect 23532 35136 23538 35148
rect 24578 35136 24584 35148
rect 23532 35108 24584 35136
rect 23532 35096 23538 35108
rect 24578 35096 24584 35108
rect 24636 35136 24642 35148
rect 25041 35139 25099 35145
rect 25041 35136 25053 35139
rect 24636 35108 25053 35136
rect 24636 35096 24642 35108
rect 25041 35105 25053 35108
rect 25087 35105 25099 35139
rect 32950 35136 32956 35148
rect 32911 35108 32956 35136
rect 25041 35099 25099 35105
rect 32950 35096 32956 35108
rect 33008 35096 33014 35148
rect 34514 35136 34520 35148
rect 34072 35108 34520 35136
rect 20809 35071 20867 35077
rect 20809 35037 20821 35071
rect 20855 35037 20867 35071
rect 20809 35031 20867 35037
rect 21269 35071 21327 35077
rect 21269 35037 21281 35071
rect 21315 35068 21327 35071
rect 21358 35068 21364 35080
rect 21315 35040 21364 35068
rect 21315 35037 21327 35040
rect 21269 35031 21327 35037
rect 20824 35000 20852 35031
rect 21358 35028 21364 35040
rect 21416 35028 21422 35080
rect 23290 35068 23296 35080
rect 23251 35040 23296 35068
rect 23290 35028 23296 35040
rect 23348 35028 23354 35080
rect 23382 35028 23388 35080
rect 23440 35068 23446 35080
rect 25308 35071 25366 35077
rect 23440 35040 23485 35068
rect 23440 35028 23446 35040
rect 25308 35037 25320 35071
rect 25354 35068 25366 35071
rect 26881 35071 26939 35077
rect 26881 35068 26893 35071
rect 25354 35040 26893 35068
rect 25354 35037 25366 35040
rect 25308 35031 25366 35037
rect 26881 35037 26893 35040
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 33220 35071 33278 35077
rect 33220 35037 33232 35071
rect 33266 35068 33278 35071
rect 34072 35068 34100 35108
rect 34514 35096 34520 35108
rect 34572 35096 34578 35148
rect 34992 35145 35020 35176
rect 34977 35139 35035 35145
rect 34977 35105 34989 35139
rect 35023 35105 35035 35139
rect 34977 35099 35035 35105
rect 33266 35040 34100 35068
rect 33266 35037 33278 35040
rect 33220 35031 33278 35037
rect 34422 35028 34428 35080
rect 34480 35068 34486 35080
rect 34885 35071 34943 35077
rect 34885 35068 34897 35071
rect 34480 35040 34897 35068
rect 34480 35028 34486 35040
rect 34885 35037 34897 35040
rect 34931 35037 34943 35071
rect 35158 35068 35164 35080
rect 35119 35040 35164 35068
rect 34885 35031 34943 35037
rect 35158 35028 35164 35040
rect 35216 35028 35222 35080
rect 36262 35068 36268 35080
rect 36223 35040 36268 35068
rect 36262 35028 36268 35040
rect 36320 35028 36326 35080
rect 36538 35077 36544 35080
rect 36532 35068 36544 35077
rect 36499 35040 36544 35068
rect 36532 35031 36544 35040
rect 36538 35028 36544 35031
rect 36596 35028 36602 35080
rect 40126 35028 40132 35080
rect 40184 35068 40190 35080
rect 40405 35071 40463 35077
rect 40405 35068 40417 35071
rect 40184 35040 40417 35068
rect 40184 35028 40190 35040
rect 40405 35037 40417 35040
rect 40451 35037 40463 35071
rect 40405 35031 40463 35037
rect 21514 35003 21572 35009
rect 21514 35000 21526 35003
rect 20824 34972 21526 35000
rect 21514 34969 21526 34972
rect 21560 34969 21572 35003
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 21514 34963 21572 34969
rect 22664 34972 23121 35000
rect 22664 34941 22692 34972
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 22649 34935 22707 34941
rect 22649 34901 22661 34935
rect 22695 34901 22707 34935
rect 22649 34895 22707 34901
rect 26421 34935 26479 34941
rect 26421 34901 26433 34935
rect 26467 34932 26479 34935
rect 26602 34932 26608 34944
rect 26467 34904 26608 34932
rect 26467 34901 26479 34904
rect 26421 34895 26479 34901
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 35345 34935 35403 34941
rect 35345 34901 35357 34935
rect 35391 34932 35403 34935
rect 37458 34932 37464 34944
rect 35391 34904 37464 34932
rect 35391 34901 35403 34904
rect 35345 34895 35403 34901
rect 37458 34892 37464 34904
rect 37516 34892 37522 34944
rect 37645 34935 37703 34941
rect 37645 34901 37657 34935
rect 37691 34932 37703 34935
rect 37734 34932 37740 34944
rect 37691 34904 37740 34932
rect 37691 34901 37703 34904
rect 37645 34895 37703 34901
rect 37734 34892 37740 34904
rect 37792 34892 37798 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 20070 34728 20076 34740
rect 20031 34700 20076 34728
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 23290 34688 23296 34740
rect 23348 34728 23354 34740
rect 23385 34731 23443 34737
rect 23385 34728 23397 34731
rect 23348 34700 23397 34728
rect 23348 34688 23354 34700
rect 23385 34697 23397 34700
rect 23431 34697 23443 34731
rect 23385 34691 23443 34697
rect 25961 34731 26019 34737
rect 25961 34697 25973 34731
rect 26007 34728 26019 34731
rect 26694 34728 26700 34740
rect 26007 34700 26700 34728
rect 26007 34697 26019 34700
rect 25961 34691 26019 34697
rect 26694 34688 26700 34700
rect 26752 34688 26758 34740
rect 34977 34731 35035 34737
rect 34977 34697 34989 34731
rect 35023 34728 35035 34731
rect 35158 34728 35164 34740
rect 35023 34700 35164 34728
rect 35023 34697 35035 34700
rect 34977 34691 35035 34697
rect 35158 34688 35164 34700
rect 35216 34688 35222 34740
rect 21208 34663 21266 34669
rect 21208 34629 21220 34663
rect 21254 34660 21266 34663
rect 22002 34660 22008 34672
rect 21254 34632 22008 34660
rect 21254 34629 21266 34632
rect 21208 34623 21266 34629
rect 22002 34620 22008 34632
rect 22060 34620 22066 34672
rect 37458 34660 37464 34672
rect 37419 34632 37464 34660
rect 37458 34620 37464 34632
rect 37516 34620 37522 34672
rect 22278 34601 22284 34604
rect 22272 34555 22284 34601
rect 22336 34592 22342 34604
rect 24578 34592 24584 34604
rect 22336 34564 22372 34592
rect 24539 34564 24584 34592
rect 22278 34552 22284 34555
rect 22336 34552 22342 34564
rect 24578 34552 24584 34564
rect 24636 34552 24642 34604
rect 24854 34601 24860 34604
rect 24848 34555 24860 34601
rect 24912 34592 24918 34604
rect 33870 34601 33876 34604
rect 24912 34564 24948 34592
rect 24854 34552 24860 34555
rect 24912 34552 24918 34564
rect 33864 34555 33876 34601
rect 33928 34592 33934 34604
rect 37734 34592 37740 34604
rect 33928 34564 33964 34592
rect 37695 34564 37740 34592
rect 33870 34552 33876 34555
rect 33928 34552 33934 34564
rect 37734 34552 37740 34564
rect 37792 34552 37798 34604
rect 39669 34595 39727 34601
rect 39669 34561 39681 34595
rect 39715 34561 39727 34595
rect 39669 34555 39727 34561
rect 21453 34527 21511 34533
rect 21453 34493 21465 34527
rect 21499 34524 21511 34527
rect 21542 34524 21548 34536
rect 21499 34496 21548 34524
rect 21499 34493 21511 34496
rect 21453 34487 21511 34493
rect 21542 34484 21548 34496
rect 21600 34524 21606 34536
rect 22005 34527 22063 34533
rect 22005 34524 22017 34527
rect 21600 34496 22017 34524
rect 21600 34484 21606 34496
rect 22005 34493 22017 34496
rect 22051 34493 22063 34527
rect 33597 34527 33655 34533
rect 33597 34524 33609 34527
rect 22005 34487 22063 34493
rect 33060 34496 33609 34524
rect 22020 34388 22048 34487
rect 23474 34456 23480 34468
rect 23308 34428 23480 34456
rect 23308 34388 23336 34428
rect 23474 34416 23480 34428
rect 23532 34416 23538 34468
rect 32306 34416 32312 34468
rect 32364 34456 32370 34468
rect 33060 34456 33088 34496
rect 33597 34493 33609 34496
rect 33643 34493 33655 34527
rect 37550 34524 37556 34536
rect 37511 34496 37556 34524
rect 33597 34487 33655 34493
rect 37550 34484 37556 34496
rect 37608 34484 37614 34536
rect 39298 34484 39304 34536
rect 39356 34524 39362 34536
rect 39684 34524 39712 34555
rect 39758 34552 39764 34604
rect 39816 34592 39822 34604
rect 39942 34592 39948 34604
rect 39816 34564 39861 34592
rect 39903 34564 39948 34592
rect 39816 34552 39822 34564
rect 39942 34552 39948 34564
rect 40000 34552 40006 34604
rect 39850 34524 39856 34536
rect 39356 34496 39856 34524
rect 39356 34484 39362 34496
rect 39850 34484 39856 34496
rect 39908 34524 39914 34536
rect 41046 34524 41052 34536
rect 39908 34496 41052 34524
rect 39908 34484 39914 34496
rect 41046 34484 41052 34496
rect 41104 34484 41110 34536
rect 32364 34428 33088 34456
rect 32364 34416 32370 34428
rect 28166 34388 28172 34400
rect 22020 34360 23336 34388
rect 28127 34360 28172 34388
rect 28166 34348 28172 34360
rect 28224 34348 28230 34400
rect 28810 34388 28816 34400
rect 28771 34360 28816 34388
rect 28810 34348 28816 34360
rect 28868 34348 28874 34400
rect 31202 34348 31208 34400
rect 31260 34388 31266 34400
rect 31297 34391 31355 34397
rect 31297 34388 31309 34391
rect 31260 34360 31309 34388
rect 31260 34348 31266 34360
rect 31297 34357 31309 34360
rect 31343 34357 31355 34391
rect 36446 34388 36452 34400
rect 36407 34360 36452 34388
rect 31297 34351 31355 34357
rect 36446 34348 36452 34360
rect 36504 34348 36510 34400
rect 37642 34388 37648 34400
rect 37603 34360 37648 34388
rect 37642 34348 37648 34360
rect 37700 34348 37706 34400
rect 37921 34391 37979 34397
rect 37921 34357 37933 34391
rect 37967 34388 37979 34391
rect 38010 34388 38016 34400
rect 37967 34360 38016 34388
rect 37967 34357 37979 34360
rect 37921 34351 37979 34357
rect 38010 34348 38016 34360
rect 38068 34348 38074 34400
rect 40129 34391 40187 34397
rect 40129 34357 40141 34391
rect 40175 34388 40187 34391
rect 40218 34388 40224 34400
rect 40175 34360 40224 34388
rect 40175 34357 40187 34360
rect 40129 34351 40187 34357
rect 40218 34348 40224 34360
rect 40276 34348 40282 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 21085 34187 21143 34193
rect 21085 34153 21097 34187
rect 21131 34184 21143 34187
rect 22278 34184 22284 34196
rect 21131 34156 22284 34184
rect 21131 34153 21143 34156
rect 21085 34147 21143 34153
rect 22278 34144 22284 34156
rect 22336 34144 22342 34196
rect 22925 34187 22983 34193
rect 22925 34153 22937 34187
rect 22971 34184 22983 34187
rect 23382 34184 23388 34196
rect 22971 34156 23388 34184
rect 22971 34153 22983 34156
rect 22925 34147 22983 34153
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 26602 34184 26608 34196
rect 26563 34156 26608 34184
rect 26602 34144 26608 34156
rect 26660 34144 26666 34196
rect 27062 34184 27068 34196
rect 27023 34156 27068 34184
rect 27062 34144 27068 34156
rect 27120 34144 27126 34196
rect 33042 34184 33048 34196
rect 33003 34156 33048 34184
rect 33042 34144 33048 34156
rect 33100 34144 33106 34196
rect 33870 34144 33876 34196
rect 33928 34184 33934 34196
rect 33965 34187 34023 34193
rect 33965 34184 33977 34187
rect 33928 34156 33977 34184
rect 33928 34144 33934 34156
rect 33965 34153 33977 34156
rect 34011 34153 34023 34187
rect 37550 34184 37556 34196
rect 37511 34156 37556 34184
rect 33965 34147 34023 34153
rect 37550 34144 37556 34156
rect 37608 34144 37614 34196
rect 39298 34184 39304 34196
rect 39259 34156 39304 34184
rect 39298 34144 39304 34156
rect 39356 34144 39362 34196
rect 39482 34184 39488 34196
rect 39443 34156 39488 34184
rect 39482 34144 39488 34156
rect 39540 34144 39546 34196
rect 40218 34184 40224 34196
rect 40179 34156 40224 34184
rect 40218 34144 40224 34156
rect 40276 34144 40282 34196
rect 26145 34119 26203 34125
rect 26145 34085 26157 34119
rect 26191 34085 26203 34119
rect 26145 34079 26203 34085
rect 32309 34119 32367 34125
rect 32309 34085 32321 34119
rect 32355 34116 32367 34119
rect 39500 34116 39528 34144
rect 40589 34119 40647 34125
rect 40589 34116 40601 34119
rect 32355 34088 32904 34116
rect 39500 34088 40601 34116
rect 32355 34085 32367 34088
rect 32309 34079 32367 34085
rect 21542 34048 21548 34060
rect 21503 34020 21548 34048
rect 21542 34008 21548 34020
rect 21600 34008 21606 34060
rect 24578 34008 24584 34060
rect 24636 34048 24642 34060
rect 24765 34051 24823 34057
rect 24765 34048 24777 34051
rect 24636 34020 24777 34048
rect 24636 34008 24642 34020
rect 24765 34017 24777 34020
rect 24811 34017 24823 34051
rect 24765 34011 24823 34017
rect 24029 33983 24087 33989
rect 24029 33949 24041 33983
rect 24075 33980 24087 33983
rect 24854 33980 24860 33992
rect 24075 33952 24860 33980
rect 24075 33949 24087 33952
rect 24029 33943 24087 33949
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 26160 33980 26188 34079
rect 26694 34048 26700 34060
rect 26655 34020 26700 34048
rect 26694 34008 26700 34020
rect 26752 34008 26758 34060
rect 27798 34048 27804 34060
rect 27759 34020 27804 34048
rect 27798 34008 27804 34020
rect 27856 34008 27862 34060
rect 32876 34057 32904 34088
rect 40589 34085 40601 34088
rect 40635 34085 40647 34119
rect 40589 34079 40647 34085
rect 32861 34051 32919 34057
rect 32861 34017 32873 34051
rect 32907 34017 32919 34051
rect 39758 34048 39764 34060
rect 32861 34011 32919 34017
rect 39132 34020 39764 34048
rect 26881 33983 26939 33989
rect 26881 33980 26893 33983
rect 26160 33952 26893 33980
rect 26881 33949 26893 33952
rect 26927 33949 26939 33983
rect 26881 33943 26939 33949
rect 28068 33983 28126 33989
rect 28068 33949 28080 33983
rect 28114 33980 28126 33983
rect 28810 33980 28816 33992
rect 28114 33952 28816 33980
rect 28114 33949 28126 33952
rect 28068 33943 28126 33949
rect 28810 33940 28816 33952
rect 28868 33940 28874 33992
rect 30466 33980 30472 33992
rect 30427 33952 30472 33980
rect 30466 33940 30472 33952
rect 30524 33940 30530 33992
rect 30929 33983 30987 33989
rect 30929 33949 30941 33983
rect 30975 33980 30987 33983
rect 31018 33980 31024 33992
rect 30975 33952 31024 33980
rect 30975 33949 30987 33952
rect 30929 33943 30987 33949
rect 31018 33940 31024 33952
rect 31076 33940 31082 33992
rect 31202 33989 31208 33992
rect 31196 33980 31208 33989
rect 31163 33952 31208 33980
rect 31196 33943 31208 33952
rect 31202 33940 31208 33943
rect 31260 33940 31266 33992
rect 32490 33940 32496 33992
rect 32548 33980 32554 33992
rect 33045 33983 33103 33989
rect 33045 33980 33057 33983
rect 32548 33952 33057 33980
rect 32548 33940 32554 33952
rect 33045 33949 33057 33952
rect 33091 33949 33103 33983
rect 33045 33943 33103 33949
rect 36173 33983 36231 33989
rect 36173 33949 36185 33983
rect 36219 33980 36231 33983
rect 36262 33980 36268 33992
rect 36219 33952 36268 33980
rect 36219 33949 36231 33952
rect 36173 33943 36231 33949
rect 36262 33940 36268 33952
rect 36320 33980 36326 33992
rect 38010 33980 38016 33992
rect 36320 33952 37412 33980
rect 37971 33952 38016 33980
rect 36320 33940 36326 33952
rect 21812 33915 21870 33921
rect 21812 33881 21824 33915
rect 21858 33912 21870 33915
rect 22002 33912 22008 33924
rect 21858 33884 22008 33912
rect 21858 33881 21870 33884
rect 21812 33875 21870 33881
rect 22002 33872 22008 33884
rect 22060 33872 22066 33924
rect 25032 33915 25090 33921
rect 25032 33881 25044 33915
rect 25078 33912 25090 33915
rect 26142 33912 26148 33924
rect 25078 33884 26148 33912
rect 25078 33881 25090 33884
rect 25032 33875 25090 33881
rect 26142 33872 26148 33884
rect 26200 33872 26206 33924
rect 26234 33872 26240 33924
rect 26292 33912 26298 33924
rect 26605 33915 26663 33921
rect 26605 33912 26617 33915
rect 26292 33884 26617 33912
rect 26292 33872 26298 33884
rect 26605 33881 26617 33884
rect 26651 33881 26663 33915
rect 26605 33875 26663 33881
rect 31754 33872 31760 33924
rect 31812 33912 31818 33924
rect 36446 33921 36452 33924
rect 32769 33915 32827 33921
rect 32769 33912 32781 33915
rect 31812 33884 32781 33912
rect 31812 33872 31818 33884
rect 32769 33881 32781 33884
rect 32815 33881 32827 33915
rect 36440 33912 36452 33921
rect 36407 33884 36452 33912
rect 32769 33875 32827 33881
rect 36440 33875 36452 33884
rect 36446 33872 36452 33875
rect 36504 33872 36510 33924
rect 37384 33912 37412 33952
rect 38010 33940 38016 33952
rect 38068 33940 38074 33992
rect 38194 33980 38200 33992
rect 38155 33952 38200 33980
rect 38194 33940 38200 33952
rect 38252 33940 38258 33992
rect 38378 33912 38384 33924
rect 37384 33884 38384 33912
rect 38378 33872 38384 33884
rect 38436 33872 38442 33924
rect 39132 33921 39160 34020
rect 39758 34008 39764 34020
rect 39816 34048 39822 34060
rect 39816 34020 41276 34048
rect 39816 34008 39822 34020
rect 41248 33992 41276 34020
rect 40310 33980 40316 33992
rect 40236 33952 40316 33980
rect 39117 33915 39175 33921
rect 39117 33881 39129 33915
rect 39163 33881 39175 33915
rect 40126 33912 40132 33924
rect 39117 33875 39175 33881
rect 39224 33884 40132 33912
rect 29181 33847 29239 33853
rect 29181 33813 29193 33847
rect 29227 33844 29239 33847
rect 29730 33844 29736 33856
rect 29227 33816 29736 33844
rect 29227 33813 29239 33816
rect 29181 33807 29239 33813
rect 29730 33804 29736 33816
rect 29788 33804 29794 33856
rect 33226 33844 33232 33856
rect 33187 33816 33232 33844
rect 33226 33804 33232 33816
rect 33284 33804 33290 33856
rect 38105 33847 38163 33853
rect 38105 33813 38117 33847
rect 38151 33844 38163 33847
rect 39224 33844 39252 33884
rect 40126 33872 40132 33884
rect 40184 33912 40190 33924
rect 40236 33921 40264 33952
rect 40310 33940 40316 33952
rect 40368 33940 40374 33992
rect 41046 33980 41052 33992
rect 41007 33952 41052 33980
rect 41046 33940 41052 33952
rect 41104 33940 41110 33992
rect 41230 33980 41236 33992
rect 41191 33952 41236 33980
rect 41230 33940 41236 33952
rect 41288 33940 41294 33992
rect 43438 33980 43444 33992
rect 43399 33952 43444 33980
rect 43438 33940 43444 33952
rect 43496 33940 43502 33992
rect 40221 33915 40279 33921
rect 40221 33912 40233 33915
rect 40184 33884 40233 33912
rect 40184 33872 40190 33884
rect 40221 33881 40233 33884
rect 40267 33881 40279 33915
rect 40221 33875 40279 33881
rect 38151 33816 39252 33844
rect 38151 33813 38163 33816
rect 38105 33807 38163 33813
rect 39298 33804 39304 33856
rect 39356 33853 39362 33856
rect 39356 33847 39375 33853
rect 39363 33813 39375 33847
rect 40034 33844 40040 33856
rect 39995 33816 40040 33844
rect 39356 33807 39375 33813
rect 39356 33804 39362 33807
rect 40034 33804 40040 33816
rect 40092 33804 40098 33856
rect 40310 33804 40316 33856
rect 40368 33844 40374 33856
rect 41141 33847 41199 33853
rect 41141 33844 41153 33847
rect 40368 33816 41153 33844
rect 40368 33804 40374 33816
rect 41141 33813 41153 33816
rect 41187 33813 41199 33847
rect 43254 33844 43260 33856
rect 43215 33816 43260 33844
rect 41141 33807 41199 33813
rect 43254 33804 43260 33816
rect 43312 33804 43318 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 24578 33600 24584 33652
rect 24636 33640 24642 33652
rect 25225 33643 25283 33649
rect 25225 33640 25237 33643
rect 24636 33612 25237 33640
rect 24636 33600 24642 33612
rect 25225 33609 25237 33612
rect 25271 33609 25283 33643
rect 25225 33603 25283 33609
rect 30466 33600 30472 33652
rect 30524 33640 30530 33652
rect 31754 33640 31760 33652
rect 30524 33612 31156 33640
rect 31715 33612 31760 33640
rect 30524 33600 30530 33612
rect 28166 33581 28172 33584
rect 28160 33572 28172 33581
rect 28127 33544 28172 33572
rect 28160 33535 28172 33544
rect 28166 33532 28172 33535
rect 28224 33532 28230 33584
rect 31018 33572 31024 33584
rect 30392 33544 31024 33572
rect 22002 33504 22008 33516
rect 21963 33476 22008 33504
rect 22002 33464 22008 33476
rect 22060 33464 22066 33516
rect 23937 33507 23995 33513
rect 23937 33473 23949 33507
rect 23983 33504 23995 33507
rect 24210 33504 24216 33516
rect 23983 33476 24216 33504
rect 23983 33473 23995 33476
rect 23937 33467 23995 33473
rect 24210 33464 24216 33476
rect 24268 33504 24274 33516
rect 26418 33504 26424 33516
rect 24268 33476 26424 33504
rect 24268 33464 24274 33476
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 30392 33513 30420 33544
rect 31018 33532 31024 33544
rect 31076 33532 31082 33584
rect 31128 33572 31156 33612
rect 31754 33600 31760 33612
rect 31812 33600 31818 33652
rect 33042 33600 33048 33652
rect 33100 33640 33106 33652
rect 33689 33643 33747 33649
rect 33689 33640 33701 33643
rect 33100 33612 33701 33640
rect 33100 33600 33106 33612
rect 33689 33609 33701 33612
rect 33735 33609 33747 33643
rect 33689 33603 33747 33609
rect 39298 33600 39304 33652
rect 39356 33640 39362 33652
rect 39942 33640 39948 33652
rect 39356 33612 39948 33640
rect 39356 33600 39362 33612
rect 39942 33600 39948 33612
rect 40000 33640 40006 33652
rect 40037 33643 40095 33649
rect 40037 33640 40049 33643
rect 40000 33612 40049 33640
rect 40000 33600 40006 33612
rect 40037 33609 40049 33612
rect 40083 33609 40095 33643
rect 40037 33603 40095 33609
rect 41230 33600 41236 33652
rect 41288 33640 41294 33652
rect 41877 33643 41935 33649
rect 41877 33640 41889 33643
rect 41288 33612 41889 33640
rect 41288 33600 41294 33612
rect 41877 33609 41889 33612
rect 41923 33609 41935 33643
rect 41877 33603 41935 33609
rect 43254 33581 43260 33584
rect 32554 33575 32612 33581
rect 32554 33572 32566 33575
rect 31128 33544 32566 33572
rect 32554 33541 32566 33544
rect 32600 33541 32612 33575
rect 43248 33572 43260 33581
rect 43215 33544 43260 33572
rect 32554 33535 32612 33541
rect 43248 33535 43260 33544
rect 43254 33532 43260 33535
rect 43312 33532 43318 33584
rect 30377 33507 30435 33513
rect 30377 33473 30389 33507
rect 30423 33473 30435 33507
rect 30377 33467 30435 33473
rect 30644 33507 30702 33513
rect 30644 33473 30656 33507
rect 30690 33504 30702 33507
rect 30926 33504 30932 33516
rect 30690 33476 30932 33504
rect 30690 33473 30702 33476
rect 30644 33467 30702 33473
rect 30926 33464 30932 33476
rect 30984 33464 30990 33516
rect 38924 33507 38982 33513
rect 38924 33473 38936 33507
rect 38970 33504 38982 33507
rect 39206 33504 39212 33516
rect 38970 33476 39212 33504
rect 38970 33473 38982 33476
rect 38924 33467 38982 33473
rect 39206 33464 39212 33476
rect 39264 33464 39270 33516
rect 40494 33504 40500 33516
rect 40455 33476 40500 33504
rect 40494 33464 40500 33476
rect 40552 33464 40558 33516
rect 40770 33513 40776 33516
rect 40764 33467 40776 33513
rect 40828 33504 40834 33516
rect 40828 33476 40864 33504
rect 40770 33464 40776 33467
rect 40828 33464 40834 33476
rect 26142 33436 26148 33448
rect 26103 33408 26148 33436
rect 26142 33396 26148 33408
rect 26200 33396 26206 33448
rect 27798 33396 27804 33448
rect 27856 33436 27862 33448
rect 27893 33439 27951 33445
rect 27893 33436 27905 33439
rect 27856 33408 27905 33436
rect 27856 33396 27862 33408
rect 27893 33405 27905 33408
rect 27939 33405 27951 33439
rect 32306 33436 32312 33448
rect 32267 33408 32312 33436
rect 27893 33399 27951 33405
rect 32306 33396 32312 33408
rect 32364 33396 32370 33448
rect 38378 33396 38384 33448
rect 38436 33436 38442 33448
rect 38657 33439 38715 33445
rect 38657 33436 38669 33439
rect 38436 33408 38669 33436
rect 38436 33396 38442 33408
rect 38657 33405 38669 33408
rect 38703 33405 38715 33439
rect 38657 33399 38715 33405
rect 42794 33396 42800 33448
rect 42852 33436 42858 33448
rect 42981 33439 43039 33445
rect 42981 33436 42993 33439
rect 42852 33408 42993 33436
rect 42852 33396 42858 33408
rect 42981 33405 42993 33408
rect 43027 33405 43039 33439
rect 42981 33399 43039 33405
rect 27433 33303 27491 33309
rect 27433 33269 27445 33303
rect 27479 33300 27491 33303
rect 27890 33300 27896 33312
rect 27479 33272 27896 33300
rect 27479 33269 27491 33272
rect 27433 33263 27491 33269
rect 27890 33260 27896 33272
rect 27948 33260 27954 33312
rect 29270 33300 29276 33312
rect 29231 33272 29276 33300
rect 29270 33260 29276 33272
rect 29328 33260 29334 33312
rect 29917 33303 29975 33309
rect 29917 33269 29929 33303
rect 29963 33300 29975 33303
rect 31386 33300 31392 33312
rect 29963 33272 31392 33300
rect 29963 33269 29975 33272
rect 29917 33263 29975 33269
rect 31386 33260 31392 33272
rect 31444 33260 31450 33312
rect 44358 33300 44364 33312
rect 44319 33272 44364 33300
rect 44358 33260 44364 33272
rect 44416 33260 44422 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 25961 33099 26019 33105
rect 25961 33065 25973 33099
rect 26007 33096 26019 33099
rect 26234 33096 26240 33108
rect 26007 33068 26240 33096
rect 26007 33065 26019 33068
rect 25961 33059 26019 33065
rect 26234 33056 26240 33068
rect 26292 33056 26298 33108
rect 26418 33096 26424 33108
rect 26379 33068 26424 33096
rect 26418 33056 26424 33068
rect 26476 33056 26482 33108
rect 29730 33096 29736 33108
rect 29691 33068 29736 33096
rect 29730 33056 29736 33068
rect 29788 33056 29794 33108
rect 32490 33096 32496 33108
rect 32451 33068 32496 33096
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 33045 33099 33103 33105
rect 33045 33065 33057 33099
rect 33091 33096 33103 33099
rect 33226 33096 33232 33108
rect 33091 33068 33232 33096
rect 33091 33065 33103 33068
rect 33045 33059 33103 33065
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 33413 33099 33471 33105
rect 33413 33065 33425 33099
rect 33459 33096 33471 33099
rect 38194 33096 38200 33108
rect 33459 33068 38200 33096
rect 33459 33065 33471 33068
rect 33413 33059 33471 33065
rect 38194 33056 38200 33068
rect 38252 33056 38258 33108
rect 39206 33096 39212 33108
rect 39167 33068 39212 33096
rect 39206 33056 39212 33068
rect 39264 33056 39270 33108
rect 40221 33099 40279 33105
rect 40221 33065 40233 33099
rect 40267 33096 40279 33099
rect 40310 33096 40316 33108
rect 40267 33068 40316 33096
rect 40267 33065 40279 33068
rect 40221 33059 40279 33065
rect 40310 33056 40316 33068
rect 40368 33056 40374 33108
rect 40770 33056 40776 33108
rect 40828 33096 40834 33108
rect 40865 33099 40923 33105
rect 40865 33096 40877 33099
rect 40828 33068 40877 33096
rect 40828 33056 40834 33068
rect 40865 33065 40877 33068
rect 40911 33065 40923 33099
rect 40865 33059 40923 33065
rect 42429 33099 42487 33105
rect 42429 33065 42441 33099
rect 42475 33096 42487 33099
rect 42475 33068 43392 33096
rect 42475 33065 42487 33068
rect 42429 33059 42487 33065
rect 43364 33040 43392 33068
rect 43438 33056 43444 33108
rect 43496 33096 43502 33108
rect 43533 33099 43591 33105
rect 43533 33096 43545 33099
rect 43496 33068 43545 33096
rect 43496 33056 43502 33068
rect 43533 33065 43545 33068
rect 43579 33065 43591 33099
rect 43533 33059 43591 33065
rect 45373 33099 45431 33105
rect 45373 33065 45385 33099
rect 45419 33065 45431 33099
rect 45373 33059 45431 33065
rect 29181 33031 29239 33037
rect 29181 32997 29193 33031
rect 29227 33028 29239 33031
rect 40405 33031 40463 33037
rect 29227 33000 29868 33028
rect 29227 32997 29239 33000
rect 29181 32991 29239 32997
rect 23290 32920 23296 32972
rect 23348 32960 23354 32972
rect 24578 32960 24584 32972
rect 23348 32932 24584 32960
rect 23348 32920 23354 32932
rect 24578 32920 24584 32932
rect 24636 32920 24642 32972
rect 29840 32969 29868 33000
rect 40405 32997 40417 33031
rect 40451 32997 40463 33031
rect 43346 33028 43352 33040
rect 43307 33000 43352 33028
rect 40405 32991 40463 32997
rect 29825 32963 29883 32969
rect 29825 32929 29837 32963
rect 29871 32929 29883 32963
rect 40034 32960 40040 32972
rect 29825 32923 29883 32929
rect 39408 32932 40040 32960
rect 27798 32892 27804 32904
rect 27759 32864 27804 32892
rect 27798 32852 27804 32864
rect 27856 32852 27862 32904
rect 27890 32852 27896 32904
rect 27948 32892 27954 32904
rect 28057 32895 28115 32901
rect 28057 32892 28069 32895
rect 27948 32864 28069 32892
rect 27948 32852 27954 32864
rect 28057 32861 28069 32864
rect 28103 32861 28115 32895
rect 28057 32855 28115 32861
rect 29270 32852 29276 32904
rect 29328 32892 29334 32904
rect 30009 32895 30067 32901
rect 30009 32892 30021 32895
rect 29328 32864 30021 32892
rect 29328 32852 29334 32864
rect 30009 32861 30021 32864
rect 30055 32861 30067 32895
rect 31110 32892 31116 32904
rect 31071 32864 31116 32892
rect 30009 32855 30067 32861
rect 31110 32852 31116 32864
rect 31168 32892 31174 32904
rect 32306 32892 32312 32904
rect 31168 32864 32312 32892
rect 31168 32852 31174 32864
rect 32306 32852 32312 32864
rect 32364 32852 32370 32904
rect 33134 32892 33140 32904
rect 33095 32864 33140 32892
rect 33134 32852 33140 32864
rect 33192 32852 33198 32904
rect 33226 32852 33232 32904
rect 33284 32892 33290 32904
rect 35069 32895 35127 32901
rect 33284 32864 33329 32892
rect 33284 32852 33290 32864
rect 35069 32861 35081 32895
rect 35115 32892 35127 32895
rect 35434 32892 35440 32904
rect 35115 32864 35440 32892
rect 35115 32861 35127 32864
rect 35069 32855 35127 32861
rect 35434 32852 35440 32864
rect 35492 32852 35498 32904
rect 39408 32901 39436 32932
rect 40034 32920 40040 32932
rect 40092 32920 40098 32972
rect 39393 32895 39451 32901
rect 39393 32861 39405 32895
rect 39439 32861 39451 32895
rect 40420 32892 40448 32991
rect 43346 32988 43352 33000
rect 43404 33028 43410 33040
rect 45388 33028 45416 33059
rect 43404 33000 45416 33028
rect 43404 32988 43410 33000
rect 41049 32895 41107 32901
rect 41049 32892 41061 32895
rect 40420 32864 41061 32892
rect 39393 32855 39451 32861
rect 41049 32861 41061 32864
rect 41095 32861 41107 32895
rect 41049 32855 41107 32861
rect 24854 32833 24860 32836
rect 24848 32787 24860 32833
rect 24912 32824 24918 32836
rect 24912 32796 24948 32824
rect 24854 32784 24860 32787
rect 24912 32784 24918 32796
rect 28902 32784 28908 32836
rect 28960 32824 28966 32836
rect 31386 32833 31392 32836
rect 29733 32827 29791 32833
rect 29733 32824 29745 32827
rect 28960 32796 29745 32824
rect 28960 32784 28966 32796
rect 29733 32793 29745 32796
rect 29779 32793 29791 32827
rect 31380 32824 31392 32833
rect 31347 32796 31392 32824
rect 29733 32787 29791 32793
rect 31380 32787 31392 32796
rect 31386 32784 31392 32787
rect 31444 32784 31450 32836
rect 32953 32827 33011 32833
rect 32953 32824 32965 32827
rect 31726 32796 32965 32824
rect 30193 32759 30251 32765
rect 30193 32725 30205 32759
rect 30239 32756 30251 32759
rect 31726 32756 31754 32796
rect 32953 32793 32965 32796
rect 32999 32793 33011 32827
rect 32953 32787 33011 32793
rect 40037 32827 40095 32833
rect 40037 32793 40049 32827
rect 40083 32824 40095 32827
rect 40126 32824 40132 32836
rect 40083 32796 40132 32824
rect 40083 32793 40095 32796
rect 40037 32787 40095 32793
rect 40126 32784 40132 32796
rect 40184 32784 40190 32836
rect 42058 32784 42064 32836
rect 42116 32824 42122 32836
rect 42613 32827 42671 32833
rect 42613 32824 42625 32827
rect 42116 32796 42625 32824
rect 42116 32784 42122 32796
rect 42613 32793 42625 32796
rect 42659 32793 42671 32827
rect 42613 32787 42671 32793
rect 43073 32827 43131 32833
rect 43073 32793 43085 32827
rect 43119 32824 43131 32827
rect 43622 32824 43628 32836
rect 43119 32796 43628 32824
rect 43119 32793 43131 32796
rect 43073 32787 43131 32793
rect 43622 32784 43628 32796
rect 43680 32824 43686 32836
rect 44358 32824 44364 32836
rect 43680 32796 44364 32824
rect 43680 32784 43686 32796
rect 44358 32784 44364 32796
rect 44416 32784 44422 32836
rect 44542 32784 44548 32836
rect 44600 32824 44606 32836
rect 45189 32827 45247 32833
rect 45189 32824 45201 32827
rect 44600 32796 45201 32824
rect 44600 32784 44606 32796
rect 45189 32793 45201 32796
rect 45235 32793 45247 32827
rect 45189 32787 45247 32793
rect 30239 32728 31754 32756
rect 30239 32725 30251 32728
rect 30193 32719 30251 32725
rect 40218 32716 40224 32768
rect 40276 32765 40282 32768
rect 40276 32759 40295 32765
rect 40283 32725 40295 32759
rect 40276 32719 40295 32725
rect 40276 32716 40282 32719
rect 41138 32716 41144 32768
rect 41196 32756 41202 32768
rect 42245 32759 42303 32765
rect 42245 32756 42257 32759
rect 41196 32728 42257 32756
rect 41196 32716 41202 32728
rect 42245 32725 42257 32728
rect 42291 32725 42303 32759
rect 42245 32719 42303 32725
rect 42413 32759 42471 32765
rect 42413 32725 42425 32759
rect 42459 32756 42471 32759
rect 42518 32756 42524 32768
rect 42459 32728 42524 32756
rect 42459 32725 42471 32728
rect 42413 32719 42471 32725
rect 42518 32716 42524 32728
rect 42576 32716 42582 32768
rect 45370 32716 45376 32768
rect 45428 32765 45434 32768
rect 45428 32759 45447 32765
rect 45435 32725 45447 32759
rect 45428 32719 45447 32725
rect 45557 32759 45615 32765
rect 45557 32725 45569 32759
rect 45603 32756 45615 32759
rect 46014 32756 46020 32768
rect 45603 32728 46020 32756
rect 45603 32725 45615 32728
rect 45557 32719 45615 32725
rect 45428 32716 45434 32719
rect 46014 32716 46020 32728
rect 46072 32716 46078 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 33226 32512 33232 32564
rect 33284 32552 33290 32564
rect 35621 32555 35679 32561
rect 35621 32552 35633 32555
rect 33284 32524 35633 32552
rect 33284 32512 33290 32524
rect 35621 32521 35633 32524
rect 35667 32521 35679 32555
rect 35621 32515 35679 32521
rect 40218 32512 40224 32564
rect 40276 32552 40282 32564
rect 40313 32555 40371 32561
rect 40313 32552 40325 32555
rect 40276 32524 40325 32552
rect 40276 32512 40282 32524
rect 40313 32521 40325 32524
rect 40359 32521 40371 32555
rect 42058 32552 42064 32564
rect 42019 32524 42064 32552
rect 40313 32515 40371 32521
rect 42058 32512 42064 32524
rect 42116 32512 42122 32564
rect 42518 32512 42524 32564
rect 42576 32552 42582 32564
rect 42613 32555 42671 32561
rect 42613 32552 42625 32555
rect 42576 32524 42625 32552
rect 42576 32512 42582 32524
rect 42613 32521 42625 32524
rect 42659 32521 42671 32555
rect 42613 32515 42671 32521
rect 42702 32512 42708 32564
rect 42760 32552 42766 32564
rect 42981 32555 43039 32561
rect 42981 32552 42993 32555
rect 42760 32524 42993 32552
rect 42760 32512 42766 32524
rect 42981 32521 42993 32524
rect 43027 32552 43039 32555
rect 43714 32552 43720 32564
rect 43027 32524 43720 32552
rect 43027 32521 43039 32524
rect 42981 32515 43039 32521
rect 43714 32512 43720 32524
rect 43772 32552 43778 32564
rect 43809 32555 43867 32561
rect 43809 32552 43821 32555
rect 43772 32524 43821 32552
rect 43772 32512 43778 32524
rect 43809 32521 43821 32524
rect 43855 32552 43867 32555
rect 45097 32555 45155 32561
rect 45097 32552 45109 32555
rect 43855 32524 45109 32552
rect 43855 32521 43867 32524
rect 43809 32515 43867 32521
rect 45097 32521 45109 32524
rect 45143 32521 45155 32555
rect 45097 32515 45155 32521
rect 36906 32484 36912 32496
rect 36819 32456 36912 32484
rect 36906 32444 36912 32456
rect 36964 32484 36970 32496
rect 37461 32487 37519 32493
rect 37461 32484 37473 32487
rect 36964 32456 37473 32484
rect 36964 32444 36970 32456
rect 37461 32453 37473 32456
rect 37507 32484 37519 32487
rect 39390 32484 39396 32496
rect 37507 32456 39396 32484
rect 37507 32453 37519 32456
rect 37461 32447 37519 32453
rect 39390 32444 39396 32456
rect 39448 32484 39454 32496
rect 44450 32484 44456 32496
rect 39448 32456 44456 32484
rect 39448 32444 39454 32456
rect 44450 32444 44456 32456
rect 44508 32444 44514 32496
rect 24765 32419 24823 32425
rect 24765 32385 24777 32419
rect 24811 32416 24823 32419
rect 24854 32416 24860 32428
rect 24811 32388 24860 32416
rect 24811 32385 24823 32388
rect 24765 32379 24823 32385
rect 24854 32376 24860 32388
rect 24912 32376 24918 32428
rect 30926 32376 30932 32428
rect 30984 32416 30990 32428
rect 31113 32419 31171 32425
rect 31113 32416 31125 32419
rect 30984 32388 31125 32416
rect 30984 32376 30990 32388
rect 31113 32385 31125 32388
rect 31159 32385 31171 32419
rect 35802 32416 35808 32428
rect 35763 32388 35808 32416
rect 31113 32379 31171 32385
rect 35802 32376 35808 32388
rect 35860 32376 35866 32428
rect 36081 32419 36139 32425
rect 36081 32385 36093 32419
rect 36127 32416 36139 32419
rect 36446 32416 36452 32428
rect 36127 32388 36452 32416
rect 36127 32385 36139 32388
rect 36081 32379 36139 32385
rect 36446 32376 36452 32388
rect 36504 32376 36510 32428
rect 39850 32376 39856 32428
rect 39908 32416 39914 32428
rect 39945 32419 40003 32425
rect 39945 32416 39957 32419
rect 39908 32388 39957 32416
rect 39908 32376 39914 32388
rect 39945 32385 39957 32388
rect 39991 32385 40003 32419
rect 39945 32379 40003 32385
rect 40129 32419 40187 32425
rect 40129 32385 40141 32419
rect 40175 32385 40187 32419
rect 41138 32416 41144 32428
rect 41099 32388 41144 32416
rect 40129 32379 40187 32385
rect 35986 32348 35992 32360
rect 35947 32320 35992 32348
rect 35986 32308 35992 32320
rect 36044 32308 36050 32360
rect 40144 32348 40172 32379
rect 41138 32376 41144 32388
rect 41196 32376 41202 32428
rect 41785 32419 41843 32425
rect 41785 32385 41797 32419
rect 41831 32385 41843 32419
rect 41785 32379 41843 32385
rect 41969 32419 42027 32425
rect 41969 32385 41981 32419
rect 42015 32385 42027 32419
rect 41969 32379 42027 32385
rect 42061 32419 42119 32425
rect 42061 32385 42073 32419
rect 42107 32416 42119 32419
rect 42794 32416 42800 32428
rect 42107 32388 42800 32416
rect 42107 32385 42119 32388
rect 42061 32379 42119 32385
rect 41230 32348 41236 32360
rect 40144 32320 41236 32348
rect 41230 32308 41236 32320
rect 41288 32308 41294 32360
rect 41800 32280 41828 32379
rect 41984 32348 42012 32379
rect 42794 32376 42800 32388
rect 42852 32376 42858 32428
rect 43073 32419 43131 32425
rect 43073 32385 43085 32419
rect 43119 32416 43131 32419
rect 43622 32416 43628 32428
rect 43119 32388 43628 32416
rect 43119 32385 43131 32388
rect 43073 32379 43131 32385
rect 43622 32376 43628 32388
rect 43680 32416 43686 32428
rect 43717 32419 43775 32425
rect 43717 32416 43729 32419
rect 43680 32388 43729 32416
rect 43680 32376 43686 32388
rect 43717 32385 43729 32388
rect 43763 32385 43775 32419
rect 43717 32379 43775 32385
rect 43901 32419 43959 32425
rect 43901 32385 43913 32419
rect 43947 32385 43959 32419
rect 46198 32416 46204 32428
rect 46256 32425 46262 32428
rect 46168 32388 46204 32416
rect 43901 32379 43959 32385
rect 42702 32348 42708 32360
rect 41984 32320 42708 32348
rect 42702 32308 42708 32320
rect 42760 32308 42766 32360
rect 42812 32348 42840 32376
rect 43916 32348 43944 32379
rect 46198 32376 46204 32388
rect 46256 32379 46268 32425
rect 46256 32376 46262 32379
rect 46474 32348 46480 32360
rect 42812 32320 43944 32348
rect 46435 32320 46480 32348
rect 46474 32308 46480 32320
rect 46532 32308 46538 32360
rect 43622 32280 43628 32292
rect 41800 32252 43628 32280
rect 43622 32240 43628 32252
rect 43680 32240 43686 32292
rect 44082 32280 44088 32292
rect 44043 32252 44088 32280
rect 44082 32240 44088 32252
rect 44140 32240 44146 32292
rect 27614 32172 27620 32224
rect 27672 32212 27678 32224
rect 27801 32215 27859 32221
rect 27801 32212 27813 32215
rect 27672 32184 27813 32212
rect 27672 32172 27678 32184
rect 27801 32181 27813 32184
rect 27847 32181 27859 32215
rect 27801 32175 27859 32181
rect 34977 32215 35035 32221
rect 34977 32181 34989 32215
rect 35023 32212 35035 32215
rect 35342 32212 35348 32224
rect 35023 32184 35348 32212
rect 35023 32181 35035 32184
rect 34977 32175 35035 32181
rect 35342 32172 35348 32184
rect 35400 32172 35406 32224
rect 36078 32212 36084 32224
rect 36039 32184 36084 32212
rect 36078 32172 36084 32184
rect 36136 32172 36142 32224
rect 38378 32172 38384 32224
rect 38436 32212 38442 32224
rect 38749 32215 38807 32221
rect 38749 32212 38761 32215
rect 38436 32184 38761 32212
rect 38436 32172 38442 32184
rect 38749 32181 38761 32184
rect 38795 32181 38807 32215
rect 38749 32175 38807 32181
rect 41325 32215 41383 32221
rect 41325 32181 41337 32215
rect 41371 32212 41383 32215
rect 41782 32212 41788 32224
rect 41371 32184 41788 32212
rect 41371 32181 41383 32184
rect 41325 32175 41383 32181
rect 41782 32172 41788 32184
rect 41840 32172 41846 32224
rect 43530 32212 43536 32224
rect 43491 32184 43536 32212
rect 43530 32172 43536 32184
rect 43588 32172 43594 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 27798 32008 27804 32020
rect 27540 31980 27804 32008
rect 24578 31832 24584 31884
rect 24636 31872 24642 31884
rect 27540 31881 27568 31980
rect 27798 31968 27804 31980
rect 27856 31968 27862 32020
rect 28902 32008 28908 32020
rect 28863 31980 28908 32008
rect 28902 31968 28908 31980
rect 28960 31968 28966 32020
rect 36078 31968 36084 32020
rect 36136 32008 36142 32020
rect 36265 32011 36323 32017
rect 36265 32008 36277 32011
rect 36136 31980 36277 32008
rect 36136 31968 36142 31980
rect 36265 31977 36277 31980
rect 36311 31977 36323 32011
rect 36265 31971 36323 31977
rect 42794 31968 42800 32020
rect 42852 32008 42858 32020
rect 42981 32011 43039 32017
rect 42981 32008 42993 32011
rect 42852 31980 42993 32008
rect 42852 31968 42858 31980
rect 42981 31977 42993 31980
rect 43027 31977 43039 32011
rect 44542 32008 44548 32020
rect 44503 31980 44548 32008
rect 42981 31971 43039 31977
rect 42996 31940 43024 31971
rect 44542 31968 44548 31980
rect 44600 31968 44606 32020
rect 45370 31968 45376 32020
rect 45428 32008 45434 32020
rect 45557 32011 45615 32017
rect 45557 32008 45569 32011
rect 45428 31980 45569 32008
rect 45428 31968 45434 31980
rect 45557 31977 45569 31980
rect 45603 31977 45615 32011
rect 46198 32008 46204 32020
rect 46159 31980 46204 32008
rect 45557 31971 45615 31977
rect 46198 31968 46204 31980
rect 46256 31968 46262 32020
rect 42996 31912 43852 31940
rect 27525 31875 27583 31881
rect 27525 31872 27537 31875
rect 24636 31844 27537 31872
rect 24636 31832 24642 31844
rect 27525 31841 27537 31844
rect 27571 31841 27583 31875
rect 27525 31835 27583 31841
rect 42886 31832 42892 31884
rect 42944 31872 42950 31884
rect 43441 31875 43499 31881
rect 43441 31872 43453 31875
rect 42944 31844 43453 31872
rect 42944 31832 42950 31844
rect 43441 31841 43453 31844
rect 43487 31841 43499 31875
rect 43714 31872 43720 31884
rect 43675 31844 43720 31872
rect 43441 31835 43499 31841
rect 43714 31832 43720 31844
rect 43772 31832 43778 31884
rect 43824 31881 43852 31912
rect 43809 31875 43867 31881
rect 43809 31841 43821 31875
rect 43855 31841 43867 31875
rect 43809 31835 43867 31841
rect 43901 31875 43959 31881
rect 43901 31841 43913 31875
rect 43947 31872 43959 31875
rect 44082 31872 44088 31884
rect 43947 31844 44088 31872
rect 43947 31841 43959 31844
rect 43901 31835 43959 31841
rect 44082 31832 44088 31844
rect 44140 31832 44146 31884
rect 44376 31844 44680 31872
rect 27614 31764 27620 31816
rect 27672 31804 27678 31816
rect 27781 31807 27839 31813
rect 27781 31804 27793 31807
rect 27672 31776 27793 31804
rect 27672 31764 27678 31776
rect 27781 31773 27793 31776
rect 27827 31773 27839 31807
rect 27781 31767 27839 31773
rect 34333 31807 34391 31813
rect 34333 31773 34345 31807
rect 34379 31804 34391 31807
rect 34698 31804 34704 31816
rect 34379 31776 34704 31804
rect 34379 31773 34391 31776
rect 34333 31767 34391 31773
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34790 31764 34796 31816
rect 34848 31804 34854 31816
rect 34885 31807 34943 31813
rect 34885 31804 34897 31807
rect 34848 31776 34897 31804
rect 34848 31764 34854 31776
rect 34885 31773 34897 31776
rect 34931 31773 34943 31807
rect 34885 31767 34943 31773
rect 35152 31807 35210 31813
rect 35152 31773 35164 31807
rect 35198 31804 35210 31807
rect 35434 31804 35440 31816
rect 35198 31776 35440 31804
rect 35198 31773 35210 31776
rect 35152 31767 35210 31773
rect 35434 31764 35440 31776
rect 35492 31764 35498 31816
rect 36722 31804 36728 31816
rect 36683 31776 36728 31804
rect 36722 31764 36728 31776
rect 36780 31764 36786 31816
rect 41601 31807 41659 31813
rect 41601 31773 41613 31807
rect 41647 31804 41659 31807
rect 41868 31807 41926 31813
rect 41647 31776 41736 31804
rect 41647 31773 41659 31776
rect 41601 31767 41659 31773
rect 41708 31668 41736 31776
rect 41868 31773 41880 31807
rect 41914 31773 41926 31807
rect 43622 31804 43628 31816
rect 43535 31776 43628 31804
rect 41868 31767 41926 31773
rect 41782 31696 41788 31748
rect 41840 31736 41846 31748
rect 41892 31736 41920 31767
rect 43622 31764 43628 31776
rect 43680 31764 43686 31816
rect 43732 31804 43760 31832
rect 44376 31804 44404 31844
rect 44652 31813 44680 31844
rect 43732 31776 44404 31804
rect 44453 31807 44511 31813
rect 44453 31773 44465 31807
rect 44499 31804 44511 31807
rect 44637 31807 44695 31813
rect 44499 31776 44588 31804
rect 44499 31773 44511 31776
rect 44453 31767 44511 31773
rect 41840 31708 41920 31736
rect 43640 31736 43668 31764
rect 44560 31736 44588 31776
rect 44637 31773 44649 31807
rect 44683 31804 44695 31807
rect 45373 31807 45431 31813
rect 45373 31804 45385 31807
rect 44683 31776 45385 31804
rect 44683 31773 44695 31776
rect 44637 31767 44695 31773
rect 45373 31773 45385 31776
rect 45419 31773 45431 31807
rect 46014 31804 46020 31816
rect 45975 31776 46020 31804
rect 45373 31767 45431 31773
rect 46014 31764 46020 31776
rect 46072 31764 46078 31816
rect 45189 31739 45247 31745
rect 45189 31736 45201 31739
rect 43640 31708 45201 31736
rect 41840 31696 41846 31708
rect 45189 31705 45201 31708
rect 45235 31705 45247 31739
rect 45189 31699 45247 31705
rect 42610 31668 42616 31680
rect 41708 31640 42616 31668
rect 42610 31628 42616 31640
rect 42668 31628 42674 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 36446 31464 36452 31476
rect 36407 31436 36452 31464
rect 36446 31424 36452 31436
rect 36504 31424 36510 31476
rect 32401 31399 32459 31405
rect 32401 31365 32413 31399
rect 32447 31396 32459 31399
rect 32490 31396 32496 31408
rect 32447 31368 32496 31396
rect 32447 31365 32459 31368
rect 32401 31359 32459 31365
rect 32490 31356 32496 31368
rect 32548 31396 32554 31408
rect 32861 31399 32919 31405
rect 32861 31396 32873 31399
rect 32548 31368 32873 31396
rect 32548 31356 32554 31368
rect 32861 31365 32873 31368
rect 32907 31396 32919 31399
rect 36906 31396 36912 31408
rect 32907 31368 36912 31396
rect 32907 31365 32919 31368
rect 32861 31359 32919 31365
rect 36906 31356 36912 31368
rect 36964 31356 36970 31408
rect 43530 31356 43536 31408
rect 43588 31396 43594 31408
rect 43717 31399 43775 31405
rect 43717 31396 43729 31399
rect 43588 31368 43729 31396
rect 43588 31356 43594 31368
rect 43717 31365 43729 31368
rect 43763 31365 43775 31399
rect 43717 31359 43775 31365
rect 44269 31399 44327 31405
rect 44269 31365 44281 31399
rect 44315 31396 44327 31399
rect 44450 31396 44456 31408
rect 44315 31368 44456 31396
rect 44315 31365 44327 31368
rect 44269 31359 44327 31365
rect 44450 31356 44456 31368
rect 44508 31356 44514 31408
rect 23201 31331 23259 31337
rect 23201 31297 23213 31331
rect 23247 31328 23259 31331
rect 23290 31328 23296 31340
rect 23247 31300 23296 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 23468 31331 23526 31337
rect 23468 31297 23480 31331
rect 23514 31328 23526 31331
rect 25130 31328 25136 31340
rect 23514 31300 25136 31328
rect 23514 31297 23526 31300
rect 23468 31291 23526 31297
rect 25130 31288 25136 31300
rect 25188 31288 25194 31340
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 35325 31331 35383 31337
rect 35325 31328 35337 31331
rect 34756 31300 35337 31328
rect 34756 31288 34762 31300
rect 35325 31297 35337 31300
rect 35371 31297 35383 31331
rect 41874 31328 41880 31340
rect 41835 31300 41880 31328
rect 35325 31291 35383 31297
rect 41874 31288 41880 31300
rect 41932 31288 41938 31340
rect 34609 31263 34667 31269
rect 34609 31229 34621 31263
rect 34655 31260 34667 31263
rect 34790 31260 34796 31272
rect 34655 31232 34796 31260
rect 34655 31229 34667 31232
rect 34609 31223 34667 31229
rect 34790 31220 34796 31232
rect 34848 31260 34854 31272
rect 35069 31263 35127 31269
rect 35069 31260 35081 31263
rect 34848 31232 35081 31260
rect 34848 31220 34854 31232
rect 35069 31229 35081 31232
rect 35115 31229 35127 31263
rect 35069 31223 35127 31229
rect 42610 31152 42616 31204
rect 42668 31192 42674 31204
rect 45557 31195 45615 31201
rect 45557 31192 45569 31195
rect 42668 31164 45569 31192
rect 42668 31152 42674 31164
rect 45557 31161 45569 31164
rect 45603 31192 45615 31195
rect 46474 31192 46480 31204
rect 45603 31164 46480 31192
rect 45603 31161 45615 31164
rect 45557 31155 45615 31161
rect 46474 31152 46480 31164
rect 46532 31152 46538 31204
rect 24578 31124 24584 31136
rect 24539 31096 24584 31124
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 30834 31124 30840 31136
rect 30795 31096 30840 31124
rect 30834 31084 30840 31096
rect 30892 31084 30898 31136
rect 31478 31124 31484 31136
rect 31439 31096 31484 31124
rect 31478 31084 31484 31096
rect 31536 31084 31542 31136
rect 42061 31127 42119 31133
rect 42061 31093 42073 31127
rect 42107 31124 42119 31127
rect 42702 31124 42708 31136
rect 42107 31096 42708 31124
rect 42107 31093 42119 31096
rect 42061 31087 42119 31093
rect 42702 31084 42708 31096
rect 42760 31084 42766 31136
rect 43622 31124 43628 31136
rect 43583 31096 43628 31124
rect 43622 31084 43628 31096
rect 43680 31084 43686 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 31941 30923 31999 30929
rect 31941 30889 31953 30923
rect 31987 30920 31999 30923
rect 32401 30923 32459 30929
rect 32401 30920 32413 30923
rect 31987 30892 32413 30920
rect 31987 30889 31999 30892
rect 31941 30883 31999 30889
rect 32401 30889 32413 30892
rect 32447 30889 32459 30923
rect 32401 30883 32459 30889
rect 32861 30923 32919 30929
rect 32861 30889 32873 30923
rect 32907 30920 32919 30923
rect 33134 30920 33140 30932
rect 32907 30892 33140 30920
rect 32907 30889 32919 30892
rect 32861 30883 32919 30889
rect 33134 30880 33140 30892
rect 33192 30880 33198 30932
rect 35986 30880 35992 30932
rect 36044 30920 36050 30932
rect 36265 30923 36323 30929
rect 36265 30920 36277 30923
rect 36044 30892 36277 30920
rect 36044 30880 36050 30892
rect 36265 30889 36277 30892
rect 36311 30889 36323 30923
rect 36265 30883 36323 30889
rect 43993 30923 44051 30929
rect 43993 30889 44005 30923
rect 44039 30920 44051 30923
rect 44082 30920 44088 30932
rect 44039 30892 44088 30920
rect 44039 30889 44051 30892
rect 43993 30883 44051 30889
rect 44082 30880 44088 30892
rect 44140 30880 44146 30932
rect 44450 30920 44456 30932
rect 44411 30892 44456 30920
rect 44450 30880 44456 30892
rect 44508 30880 44514 30932
rect 31754 30744 31760 30796
rect 31812 30784 31818 30796
rect 32493 30787 32551 30793
rect 32493 30784 32505 30787
rect 31812 30756 32505 30784
rect 31812 30744 31818 30756
rect 32493 30753 32505 30756
rect 32539 30753 32551 30787
rect 32493 30747 32551 30753
rect 23566 30716 23572 30728
rect 23527 30688 23572 30716
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30561 30719 30619 30725
rect 30561 30716 30573 30719
rect 30432 30688 30573 30716
rect 30432 30676 30438 30688
rect 30561 30685 30573 30688
rect 30607 30716 30619 30719
rect 31110 30716 31116 30728
rect 30607 30688 31116 30716
rect 30607 30685 30619 30688
rect 30561 30679 30619 30685
rect 31110 30676 31116 30688
rect 31168 30716 31174 30728
rect 31386 30716 31392 30728
rect 31168 30688 31392 30716
rect 31168 30676 31174 30688
rect 31386 30676 31392 30688
rect 31444 30676 31450 30728
rect 32674 30716 32680 30728
rect 32635 30688 32680 30716
rect 32674 30676 32680 30688
rect 32732 30676 32738 30728
rect 34790 30676 34796 30728
rect 34848 30716 34854 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34848 30688 34897 30716
rect 34848 30676 34854 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 42610 30716 42616 30728
rect 42571 30688 42616 30716
rect 34885 30679 34943 30685
rect 42610 30676 42616 30688
rect 42668 30676 42674 30728
rect 42702 30676 42708 30728
rect 42760 30716 42766 30728
rect 42869 30719 42927 30725
rect 42869 30716 42881 30719
rect 42760 30688 42881 30716
rect 42760 30676 42766 30688
rect 42869 30685 42881 30688
rect 42915 30685 42927 30719
rect 42869 30679 42927 30685
rect 30834 30657 30840 30660
rect 30828 30648 30840 30657
rect 30795 30620 30840 30648
rect 30828 30611 30840 30620
rect 30834 30608 30840 30611
rect 30892 30608 30898 30660
rect 32398 30648 32404 30660
rect 32359 30620 32404 30648
rect 32398 30608 32404 30620
rect 32456 30608 32462 30660
rect 35152 30651 35210 30657
rect 35152 30617 35164 30651
rect 35198 30648 35210 30651
rect 35342 30648 35348 30660
rect 35198 30620 35348 30648
rect 35198 30617 35210 30620
rect 35152 30611 35210 30617
rect 35342 30608 35348 30620
rect 35400 30608 35406 30660
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 31386 30336 31392 30388
rect 31444 30376 31450 30388
rect 34790 30376 34796 30388
rect 31444 30348 34796 30376
rect 31444 30336 31450 30348
rect 34790 30336 34796 30348
rect 34848 30336 34854 30388
rect 41874 30336 41880 30388
rect 41932 30376 41938 30388
rect 42705 30379 42763 30385
rect 42705 30376 42717 30379
rect 41932 30348 42717 30376
rect 41932 30336 41938 30348
rect 42705 30345 42717 30348
rect 42751 30345 42763 30379
rect 42705 30339 42763 30345
rect 23566 30317 23572 30320
rect 23560 30308 23572 30317
rect 23527 30280 23572 30308
rect 23560 30271 23572 30280
rect 23566 30268 23572 30271
rect 23624 30268 23630 30320
rect 30644 30311 30702 30317
rect 30644 30277 30656 30311
rect 30690 30308 30702 30311
rect 31478 30308 31484 30320
rect 30690 30280 31484 30308
rect 30690 30277 30702 30280
rect 30644 30271 30702 30277
rect 31478 30268 31484 30280
rect 31536 30268 31542 30320
rect 35928 30311 35986 30317
rect 35928 30277 35940 30311
rect 35974 30308 35986 30311
rect 36722 30308 36728 30320
rect 35974 30280 36728 30308
rect 35974 30277 35986 30280
rect 35928 30271 35986 30277
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 42886 30308 42892 30320
rect 42847 30280 42892 30308
rect 42886 30268 42892 30280
rect 42944 30268 42950 30320
rect 25130 30240 25136 30252
rect 25091 30212 25136 30240
rect 25130 30200 25136 30212
rect 25188 30200 25194 30252
rect 30374 30240 30380 30252
rect 30335 30212 30380 30240
rect 30374 30200 30380 30212
rect 30432 30200 30438 30252
rect 43070 30200 43076 30252
rect 43128 30240 43134 30252
rect 43257 30243 43315 30249
rect 43257 30240 43269 30243
rect 43128 30212 43269 30240
rect 43128 30200 43134 30212
rect 43257 30209 43269 30212
rect 43303 30240 43315 30243
rect 43622 30240 43628 30252
rect 43303 30212 43628 30240
rect 43303 30209 43315 30212
rect 43257 30203 43315 30209
rect 43622 30200 43628 30212
rect 43680 30200 43686 30252
rect 23290 30172 23296 30184
rect 23251 30144 23296 30172
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 36173 30175 36231 30181
rect 36173 30141 36185 30175
rect 36219 30172 36231 30175
rect 38378 30172 38384 30184
rect 36219 30144 38384 30172
rect 36219 30141 36231 30144
rect 36173 30135 36231 30141
rect 38378 30132 38384 30144
rect 38436 30132 38442 30184
rect 31754 30104 31760 30116
rect 31715 30076 31760 30104
rect 31754 30064 31760 30076
rect 31812 30064 31818 30116
rect 22830 30036 22836 30048
rect 22791 30008 22836 30036
rect 22830 29996 22836 30008
rect 22888 29996 22894 30048
rect 24670 30036 24676 30048
rect 24631 30008 24676 30036
rect 24670 29996 24676 30008
rect 24728 29996 24734 30048
rect 31938 29996 31944 30048
rect 31996 30036 32002 30048
rect 32309 30039 32367 30045
rect 32309 30036 32321 30039
rect 31996 30008 32321 30036
rect 31996 29996 32002 30008
rect 32309 30005 32321 30008
rect 32355 30005 32367 30039
rect 32309 29999 32367 30005
rect 34793 30039 34851 30045
rect 34793 30005 34805 30039
rect 34839 30036 34851 30039
rect 35802 30036 35808 30048
rect 34839 30008 35808 30036
rect 34839 30005 34851 30008
rect 34793 29999 34851 30005
rect 35802 29996 35808 30008
rect 35860 29996 35866 30048
rect 42889 30039 42947 30045
rect 42889 30005 42901 30039
rect 42935 30036 42947 30039
rect 43346 30036 43352 30048
rect 42935 30008 43352 30036
rect 42935 30005 42947 30008
rect 42889 29999 42947 30005
rect 43346 29996 43352 30008
rect 43404 29996 43410 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 24670 29832 24676 29844
rect 24631 29804 24676 29832
rect 24670 29792 24676 29804
rect 24728 29792 24734 29844
rect 32674 29792 32680 29844
rect 32732 29832 32738 29844
rect 32769 29835 32827 29841
rect 32769 29832 32781 29835
rect 32732 29804 32781 29832
rect 32732 29792 32738 29804
rect 32769 29801 32781 29804
rect 32815 29801 32827 29835
rect 32769 29795 32827 29801
rect 24578 29656 24584 29708
rect 24636 29696 24642 29708
rect 24673 29699 24731 29705
rect 24673 29696 24685 29699
rect 24636 29668 24685 29696
rect 24636 29656 24642 29668
rect 24673 29665 24685 29668
rect 24719 29665 24731 29699
rect 31386 29696 31392 29708
rect 31347 29668 31392 29696
rect 24673 29659 24731 29665
rect 31386 29656 31392 29668
rect 31444 29656 31450 29708
rect 22097 29631 22155 29637
rect 22097 29597 22109 29631
rect 22143 29597 22155 29631
rect 22097 29591 22155 29597
rect 22557 29631 22615 29637
rect 22557 29597 22569 29631
rect 22603 29628 22615 29631
rect 23290 29628 23296 29640
rect 22603 29600 23296 29628
rect 22603 29597 22615 29600
rect 22557 29591 22615 29597
rect 22112 29560 22140 29591
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 24854 29628 24860 29640
rect 24815 29600 24860 29628
rect 24854 29588 24860 29600
rect 24912 29588 24918 29640
rect 30282 29588 30288 29640
rect 30340 29628 30346 29640
rect 30377 29631 30435 29637
rect 30377 29628 30389 29631
rect 30340 29600 30389 29628
rect 30340 29588 30346 29600
rect 30377 29597 30389 29600
rect 30423 29597 30435 29631
rect 30377 29591 30435 29597
rect 31656 29631 31714 29637
rect 31656 29597 31668 29631
rect 31702 29628 31714 29631
rect 31938 29628 31944 29640
rect 31702 29600 31944 29628
rect 31702 29597 31714 29600
rect 31656 29591 31714 29597
rect 31938 29588 31944 29600
rect 31996 29588 32002 29640
rect 43898 29588 43904 29640
rect 43956 29628 43962 29640
rect 44361 29631 44419 29637
rect 44361 29628 44373 29631
rect 43956 29600 44373 29628
rect 43956 29588 43962 29600
rect 44361 29597 44373 29600
rect 44407 29597 44419 29631
rect 44361 29591 44419 29597
rect 46474 29588 46480 29640
rect 46532 29628 46538 29640
rect 46569 29631 46627 29637
rect 46569 29628 46581 29631
rect 46532 29600 46581 29628
rect 46532 29588 46538 29600
rect 46569 29597 46581 29600
rect 46615 29597 46627 29631
rect 46569 29591 46627 29597
rect 22802 29563 22860 29569
rect 22802 29560 22814 29563
rect 22112 29532 22814 29560
rect 22802 29529 22814 29532
rect 22848 29529 22860 29563
rect 24581 29563 24639 29569
rect 24581 29560 24593 29563
rect 22802 29523 22860 29529
rect 23952 29532 24593 29560
rect 23952 29501 23980 29532
rect 24581 29529 24593 29532
rect 24627 29529 24639 29563
rect 46302 29563 46360 29569
rect 46302 29560 46314 29563
rect 24581 29523 24639 29529
rect 44560 29532 46314 29560
rect 23937 29495 23995 29501
rect 23937 29461 23949 29495
rect 23983 29461 23995 29495
rect 23937 29455 23995 29461
rect 25041 29495 25099 29501
rect 25041 29461 25053 29495
rect 25087 29492 25099 29495
rect 25130 29492 25136 29504
rect 25087 29464 25136 29492
rect 25087 29461 25099 29464
rect 25041 29455 25099 29461
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 44560 29501 44588 29532
rect 46302 29529 46314 29532
rect 46348 29529 46360 29563
rect 46302 29523 46360 29529
rect 44545 29495 44603 29501
rect 44545 29461 44557 29495
rect 44591 29461 44603 29495
rect 44545 29455 44603 29461
rect 44634 29452 44640 29504
rect 44692 29492 44698 29504
rect 45189 29495 45247 29501
rect 45189 29492 45201 29495
rect 44692 29464 45201 29492
rect 44692 29452 44698 29464
rect 45189 29461 45201 29464
rect 45235 29461 45247 29495
rect 45189 29455 45247 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 24673 29291 24731 29297
rect 24673 29257 24685 29291
rect 24719 29288 24731 29291
rect 24854 29288 24860 29300
rect 24719 29260 24860 29288
rect 24719 29257 24731 29260
rect 24673 29251 24731 29257
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 31389 29291 31447 29297
rect 31389 29257 31401 29291
rect 31435 29288 31447 29291
rect 32398 29288 32404 29300
rect 31435 29260 32404 29288
rect 31435 29257 31447 29260
rect 31389 29251 31447 29257
rect 32398 29248 32404 29260
rect 32456 29248 32462 29300
rect 43898 29288 43904 29300
rect 43859 29260 43904 29288
rect 43898 29248 43904 29260
rect 43956 29248 43962 29300
rect 22830 29180 22836 29232
rect 22888 29220 22894 29232
rect 23538 29223 23596 29229
rect 23538 29220 23550 29223
rect 22888 29192 23550 29220
rect 22888 29180 22894 29192
rect 23538 29189 23550 29192
rect 23584 29189 23596 29223
rect 30374 29220 30380 29232
rect 23538 29183 23596 29189
rect 30024 29192 30380 29220
rect 23290 29152 23296 29164
rect 23251 29124 23296 29152
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 30024 29161 30052 29192
rect 30374 29180 30380 29192
rect 30432 29180 30438 29232
rect 42981 29223 43039 29229
rect 42981 29189 42993 29223
rect 43027 29220 43039 29223
rect 43533 29223 43591 29229
rect 43533 29220 43545 29223
rect 43027 29192 43545 29220
rect 43027 29189 43039 29192
rect 42981 29183 43039 29189
rect 43533 29189 43545 29192
rect 43579 29189 43591 29223
rect 43533 29183 43591 29189
rect 43749 29223 43807 29229
rect 43749 29189 43761 29223
rect 43795 29220 43807 29223
rect 44361 29223 44419 29229
rect 44361 29220 44373 29223
rect 43795 29192 44373 29220
rect 43795 29189 43807 29192
rect 43749 29183 43807 29189
rect 44361 29189 44373 29192
rect 44407 29189 44419 29223
rect 45278 29220 45284 29232
rect 44361 29183 44419 29189
rect 44468 29192 44864 29220
rect 45239 29192 45284 29220
rect 30282 29161 30288 29164
rect 30009 29155 30067 29161
rect 30009 29121 30021 29155
rect 30055 29121 30067 29155
rect 30276 29152 30288 29161
rect 30243 29124 30288 29152
rect 30009 29115 30067 29121
rect 30276 29115 30288 29124
rect 30282 29112 30288 29115
rect 30340 29112 30346 29164
rect 42889 29155 42947 29161
rect 42889 29121 42901 29155
rect 42935 29121 42947 29155
rect 43070 29152 43076 29164
rect 43031 29124 43076 29152
rect 42889 29115 42947 29121
rect 42904 29084 42932 29115
rect 43070 29112 43076 29124
rect 43128 29152 43134 29164
rect 44468 29152 44496 29192
rect 43128 29124 44496 29152
rect 43128 29112 43134 29124
rect 44542 29112 44548 29164
rect 44600 29152 44606 29164
rect 44726 29152 44732 29164
rect 44600 29124 44645 29152
rect 44687 29124 44732 29152
rect 44600 29112 44606 29124
rect 44726 29112 44732 29124
rect 44784 29112 44790 29164
rect 44836 29161 44864 29192
rect 45278 29180 45284 29192
rect 45336 29180 45342 29232
rect 45370 29180 45376 29232
rect 45428 29220 45434 29232
rect 45481 29223 45539 29229
rect 45481 29220 45493 29223
rect 45428 29192 45493 29220
rect 45428 29180 45434 29192
rect 45481 29189 45493 29192
rect 45527 29189 45539 29223
rect 45481 29183 45539 29189
rect 44821 29155 44879 29161
rect 44821 29121 44833 29155
rect 44867 29121 44879 29155
rect 46109 29155 46167 29161
rect 46109 29152 46121 29155
rect 44821 29115 44879 29121
rect 45664 29124 46121 29152
rect 43254 29084 43260 29096
rect 42904 29056 43260 29084
rect 43254 29044 43260 29056
rect 43312 29044 43318 29096
rect 35434 28976 35440 29028
rect 35492 29016 35498 29028
rect 35529 29019 35587 29025
rect 35529 29016 35541 29019
rect 35492 28988 35541 29016
rect 35492 28976 35498 28988
rect 35529 28985 35541 28988
rect 35575 28985 35587 29019
rect 38654 29016 38660 29028
rect 38615 28988 38660 29016
rect 35529 28979 35587 28985
rect 38654 28976 38660 28988
rect 38712 28976 38718 29028
rect 45664 29025 45692 29124
rect 46109 29121 46121 29124
rect 46155 29121 46167 29155
rect 46109 29115 46167 29121
rect 45649 29019 45707 29025
rect 45649 28985 45661 29019
rect 45695 28985 45707 29019
rect 45649 28979 45707 28985
rect 17310 28948 17316 28960
rect 17271 28920 17316 28948
rect 17310 28908 17316 28920
rect 17368 28908 17374 28960
rect 18322 28948 18328 28960
rect 18283 28920 18328 28948
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 36170 28948 36176 28960
rect 36131 28920 36176 28948
rect 36170 28908 36176 28920
rect 36228 28908 36234 28960
rect 42886 28908 42892 28960
rect 42944 28948 42950 28960
rect 43346 28948 43352 28960
rect 42944 28920 43352 28948
rect 42944 28908 42950 28920
rect 43346 28908 43352 28920
rect 43404 28948 43410 28960
rect 43717 28951 43775 28957
rect 43717 28948 43729 28951
rect 43404 28920 43729 28948
rect 43404 28908 43410 28920
rect 43717 28917 43729 28920
rect 43763 28948 43775 28951
rect 45465 28951 45523 28957
rect 45465 28948 45477 28951
rect 43763 28920 45477 28948
rect 43763 28917 43775 28920
rect 43717 28911 43775 28917
rect 45465 28917 45477 28920
rect 45511 28917 45523 28951
rect 46290 28948 46296 28960
rect 46251 28920 46296 28948
rect 45465 28911 45523 28917
rect 46290 28908 46296 28920
rect 46348 28908 46354 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 31754 28704 31760 28756
rect 31812 28744 31818 28756
rect 32490 28744 32496 28756
rect 31812 28716 32496 28744
rect 31812 28704 31818 28716
rect 32490 28704 32496 28716
rect 32548 28704 32554 28756
rect 44634 28608 44640 28620
rect 44595 28580 44640 28608
rect 44634 28568 44640 28580
rect 44692 28568 44698 28620
rect 16942 28500 16948 28552
rect 17000 28540 17006 28552
rect 17310 28549 17316 28552
rect 17037 28543 17095 28549
rect 17037 28540 17049 28543
rect 17000 28512 17049 28540
rect 17000 28500 17006 28512
rect 17037 28509 17049 28512
rect 17083 28509 17095 28543
rect 17304 28540 17316 28549
rect 17271 28512 17316 28540
rect 17037 28503 17095 28509
rect 17304 28503 17316 28512
rect 17310 28500 17316 28503
rect 17368 28500 17374 28552
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28540 24823 28543
rect 24854 28540 24860 28552
rect 24811 28512 24860 28540
rect 24811 28509 24823 28512
rect 24765 28503 24823 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 35066 28540 35072 28552
rect 34848 28512 35072 28540
rect 34848 28500 34854 28512
rect 35066 28500 35072 28512
rect 35124 28540 35130 28552
rect 35253 28543 35311 28549
rect 35253 28540 35265 28543
rect 35124 28512 35265 28540
rect 35124 28500 35130 28512
rect 35253 28509 35265 28512
rect 35299 28509 35311 28543
rect 38746 28540 38752 28552
rect 38707 28512 38752 28540
rect 35253 28503 35311 28509
rect 38746 28500 38752 28512
rect 38804 28500 38810 28552
rect 42978 28540 42984 28552
rect 42939 28512 42984 28540
rect 42978 28500 42984 28512
rect 43036 28500 43042 28552
rect 43254 28540 43260 28552
rect 43215 28512 43260 28540
rect 43254 28500 43260 28512
rect 43312 28540 43318 28552
rect 43714 28540 43720 28552
rect 43312 28512 43720 28540
rect 43312 28500 43318 28512
rect 43714 28500 43720 28512
rect 43772 28540 43778 28552
rect 44269 28543 44327 28549
rect 44269 28540 44281 28543
rect 43772 28512 44281 28540
rect 43772 28500 43778 28512
rect 44269 28509 44281 28512
rect 44315 28509 44327 28543
rect 44269 28503 44327 28509
rect 44453 28543 44511 28549
rect 44453 28509 44465 28543
rect 44499 28540 44511 28543
rect 44726 28540 44732 28552
rect 44499 28512 44732 28540
rect 44499 28509 44511 28512
rect 44453 28503 44511 28509
rect 44726 28500 44732 28512
rect 44784 28540 44790 28552
rect 44784 28512 45232 28540
rect 44784 28500 44790 28512
rect 31205 28475 31263 28481
rect 31205 28441 31217 28475
rect 31251 28441 31263 28475
rect 31205 28435 31263 28441
rect 35520 28475 35578 28481
rect 35520 28441 35532 28475
rect 35566 28472 35578 28475
rect 36170 28472 36176 28484
rect 35566 28444 36176 28472
rect 35566 28441 35578 28444
rect 35520 28435 35578 28441
rect 18417 28407 18475 28413
rect 18417 28373 18429 28407
rect 18463 28404 18475 28407
rect 20070 28404 20076 28416
rect 18463 28376 20076 28404
rect 18463 28373 18475 28376
rect 18417 28367 18475 28373
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 30650 28404 30656 28416
rect 30611 28376 30656 28404
rect 30650 28364 30656 28376
rect 30708 28404 30714 28416
rect 31220 28404 31248 28435
rect 36170 28432 36176 28444
rect 36228 28432 36234 28484
rect 43070 28432 43076 28484
rect 43128 28472 43134 28484
rect 43165 28475 43223 28481
rect 43165 28472 43177 28475
rect 43128 28444 43177 28472
rect 43128 28432 43134 28444
rect 43165 28441 43177 28444
rect 43211 28441 43223 28475
rect 43165 28435 43223 28441
rect 45204 28416 45232 28512
rect 46290 28500 46296 28552
rect 46348 28549 46354 28552
rect 46348 28540 46360 28549
rect 46348 28512 46393 28540
rect 46348 28503 46360 28512
rect 46348 28500 46354 28503
rect 46474 28500 46480 28552
rect 46532 28540 46538 28552
rect 46569 28543 46627 28549
rect 46569 28540 46581 28543
rect 46532 28512 46581 28540
rect 46532 28500 46538 28512
rect 46569 28509 46581 28512
rect 46615 28509 46627 28543
rect 46569 28503 46627 28509
rect 30708 28376 31248 28404
rect 36633 28407 36691 28413
rect 30708 28364 30714 28376
rect 36633 28373 36645 28407
rect 36679 28404 36691 28407
rect 37642 28404 37648 28416
rect 36679 28376 37648 28404
rect 36679 28373 36691 28376
rect 36633 28367 36691 28373
rect 37642 28364 37648 28376
rect 37700 28364 37706 28416
rect 42794 28404 42800 28416
rect 42755 28376 42800 28404
rect 42794 28364 42800 28376
rect 42852 28364 42858 28416
rect 45186 28404 45192 28416
rect 45147 28376 45192 28404
rect 45186 28364 45192 28376
rect 45244 28364 45250 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 19429 28203 19487 28209
rect 19429 28169 19441 28203
rect 19475 28169 19487 28203
rect 19429 28163 19487 28169
rect 36449 28203 36507 28209
rect 36449 28169 36461 28203
rect 36495 28200 36507 28203
rect 42061 28203 42119 28209
rect 36495 28172 37504 28200
rect 36495 28169 36507 28172
rect 36449 28163 36507 28169
rect 18322 28141 18328 28144
rect 18316 28132 18328 28141
rect 18283 28104 18328 28132
rect 18316 28095 18328 28104
rect 18322 28092 18328 28095
rect 18380 28092 18386 28144
rect 19444 28132 19472 28163
rect 37476 28141 37504 28172
rect 42061 28169 42073 28203
rect 42107 28169 42119 28203
rect 42061 28163 42119 28169
rect 35314 28135 35372 28141
rect 35314 28132 35326 28135
rect 19444 28104 20208 28132
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19392 28036 19901 28064
rect 19392 28024 19398 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 20070 28064 20076 28076
rect 20031 28036 20076 28064
rect 19889 28027 19947 28033
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20180 28073 20208 28104
rect 34624 28104 35326 28132
rect 34624 28073 34652 28104
rect 35314 28101 35326 28104
rect 35360 28101 35372 28135
rect 35314 28095 35372 28101
rect 37461 28135 37519 28141
rect 37461 28101 37473 28135
rect 37507 28101 37519 28135
rect 37461 28095 37519 28101
rect 38648 28135 38706 28141
rect 38648 28101 38660 28135
rect 38694 28132 38706 28135
rect 38746 28132 38752 28144
rect 38694 28104 38752 28132
rect 38694 28101 38706 28104
rect 38648 28095 38706 28101
rect 38746 28092 38752 28104
rect 38804 28092 38810 28144
rect 42076 28132 42104 28163
rect 42978 28160 42984 28212
rect 43036 28200 43042 28212
rect 43898 28200 43904 28212
rect 43036 28172 43904 28200
rect 43036 28160 43042 28172
rect 43898 28160 43904 28172
rect 43956 28200 43962 28212
rect 43993 28203 44051 28209
rect 43993 28200 44005 28203
rect 43956 28172 44005 28200
rect 43956 28160 43962 28172
rect 43993 28169 44005 28172
rect 44039 28169 44051 28203
rect 43993 28163 44051 28169
rect 45281 28203 45339 28209
rect 45281 28169 45293 28203
rect 45327 28200 45339 28203
rect 45370 28200 45376 28212
rect 45327 28172 45376 28200
rect 45327 28169 45339 28172
rect 45281 28163 45339 28169
rect 45370 28160 45376 28172
rect 45428 28160 45434 28212
rect 42858 28135 42916 28141
rect 42858 28132 42870 28135
rect 42076 28104 42870 28132
rect 42858 28101 42870 28104
rect 42904 28101 42916 28135
rect 42858 28095 42916 28101
rect 43070 28092 43076 28144
rect 43128 28132 43134 28144
rect 44910 28132 44916 28144
rect 43128 28104 44916 28132
rect 43128 28092 43134 28104
rect 44910 28092 44916 28104
rect 44968 28092 44974 28144
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28033 20223 28067
rect 23385 28067 23443 28073
rect 23385 28064 23397 28067
rect 20165 28027 20223 28033
rect 22848 28036 23397 28064
rect 16942 27956 16948 28008
rect 17000 27996 17006 28008
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 17000 27968 18061 27996
rect 17000 27956 17006 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 22848 27937 22876 28036
rect 23385 28033 23397 28036
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 34609 28067 34667 28073
rect 34609 28033 34621 28067
rect 34655 28033 34667 28067
rect 35066 28064 35072 28076
rect 35027 28036 35072 28064
rect 34609 28027 34667 28033
rect 35066 28024 35072 28036
rect 35124 28024 35130 28076
rect 37642 28064 37648 28076
rect 37603 28036 37648 28064
rect 37642 28024 37648 28036
rect 37700 28024 37706 28076
rect 37734 28024 37740 28076
rect 37792 28064 37798 28076
rect 38378 28064 38384 28076
rect 37792 28036 37837 28064
rect 38339 28036 38384 28064
rect 37792 28024 37798 28036
rect 38378 28024 38384 28036
rect 38436 28024 38442 28076
rect 41874 28064 41880 28076
rect 41835 28036 41880 28064
rect 41874 28024 41880 28036
rect 41932 28024 41938 28076
rect 42610 28064 42616 28076
rect 42571 28036 42616 28064
rect 42610 28024 42616 28036
rect 42668 28024 42674 28076
rect 45097 28067 45155 28073
rect 45097 28033 45109 28067
rect 45143 28064 45155 28067
rect 45186 28064 45192 28076
rect 45143 28036 45192 28064
rect 45143 28033 45155 28036
rect 45097 28027 45155 28033
rect 45186 28024 45192 28036
rect 45244 28064 45250 28076
rect 45370 28064 45376 28076
rect 45244 28036 45376 28064
rect 45244 28024 45250 28036
rect 45370 28024 45376 28036
rect 45428 28024 45434 28076
rect 22833 27931 22891 27937
rect 22833 27928 22845 27931
rect 6886 27900 18092 27928
rect 3418 27820 3424 27872
rect 3476 27860 3482 27872
rect 6886 27860 6914 27900
rect 3476 27832 6914 27860
rect 16301 27863 16359 27869
rect 3476 27820 3482 27832
rect 16301 27829 16313 27863
rect 16347 27860 16359 27863
rect 16758 27860 16764 27872
rect 16347 27832 16764 27860
rect 16347 27829 16359 27832
rect 16301 27823 16359 27829
rect 16758 27820 16764 27832
rect 16816 27820 16822 27872
rect 17310 27860 17316 27872
rect 17271 27832 17316 27860
rect 17310 27820 17316 27832
rect 17368 27820 17374 27872
rect 18064 27860 18092 27900
rect 19352 27900 22845 27928
rect 19352 27860 19380 27900
rect 22833 27897 22845 27900
rect 22879 27897 22891 27931
rect 30650 27928 30656 27940
rect 22833 27891 22891 27897
rect 24688 27900 30656 27928
rect 24688 27872 24716 27900
rect 30650 27888 30656 27900
rect 30708 27888 30714 27940
rect 19886 27860 19892 27872
rect 18064 27832 19380 27860
rect 19847 27832 19892 27860
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 20346 27860 20352 27872
rect 20307 27832 20352 27860
rect 20346 27820 20352 27832
rect 20404 27820 20410 27872
rect 20990 27820 20996 27872
rect 21048 27860 21054 27872
rect 21085 27863 21143 27869
rect 21085 27860 21097 27863
rect 21048 27832 21097 27860
rect 21048 27820 21054 27832
rect 21085 27829 21097 27832
rect 21131 27829 21143 27863
rect 24670 27860 24676 27872
rect 24631 27832 24676 27860
rect 21085 27823 21143 27829
rect 24670 27820 24676 27832
rect 24728 27820 24734 27872
rect 25590 27860 25596 27872
rect 25551 27832 25596 27860
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 28626 27860 28632 27872
rect 28587 27832 28632 27860
rect 28626 27820 28632 27832
rect 28684 27820 28690 27872
rect 31938 27820 31944 27872
rect 31996 27860 32002 27872
rect 32309 27863 32367 27869
rect 32309 27860 32321 27863
rect 31996 27832 32321 27860
rect 31996 27820 32002 27832
rect 32309 27829 32321 27832
rect 32355 27829 32367 27863
rect 32950 27860 32956 27872
rect 32911 27832 32956 27860
rect 32309 27823 32367 27829
rect 32950 27820 32956 27832
rect 33008 27820 33014 27872
rect 37458 27860 37464 27872
rect 37419 27832 37464 27860
rect 37458 27820 37464 27832
rect 37516 27820 37522 27872
rect 37918 27860 37924 27872
rect 37879 27832 37924 27860
rect 37918 27820 37924 27832
rect 37976 27820 37982 27872
rect 39761 27863 39819 27869
rect 39761 27829 39773 27863
rect 39807 27860 39819 27863
rect 40034 27860 40040 27872
rect 39807 27832 40040 27860
rect 39807 27829 39819 27832
rect 39761 27823 39819 27829
rect 40034 27820 40040 27832
rect 40092 27820 40098 27872
rect 40126 27820 40132 27872
rect 40184 27860 40190 27872
rect 40221 27863 40279 27869
rect 40221 27860 40233 27863
rect 40184 27832 40233 27860
rect 40184 27820 40190 27832
rect 40221 27829 40233 27832
rect 40267 27829 40279 27863
rect 40221 27823 40279 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 41874 27616 41880 27668
rect 41932 27656 41938 27668
rect 42521 27659 42579 27665
rect 42521 27656 42533 27659
rect 41932 27628 42533 27656
rect 41932 27616 41938 27628
rect 42521 27625 42533 27628
rect 42567 27625 42579 27659
rect 42521 27619 42579 27625
rect 42705 27659 42763 27665
rect 42705 27625 42717 27659
rect 42751 27656 42763 27659
rect 42886 27656 42892 27668
rect 42751 27628 42892 27656
rect 42751 27625 42763 27628
rect 42705 27619 42763 27625
rect 42886 27616 42892 27628
rect 42944 27616 42950 27668
rect 43162 27616 43168 27668
rect 43220 27656 43226 27668
rect 43717 27659 43775 27665
rect 43717 27656 43729 27659
rect 43220 27628 43729 27656
rect 43220 27616 43226 27628
rect 43717 27625 43729 27628
rect 43763 27625 43775 27659
rect 43717 27619 43775 27625
rect 18417 27591 18475 27597
rect 18417 27557 18429 27591
rect 18463 27588 18475 27591
rect 19886 27588 19892 27600
rect 18463 27560 19892 27588
rect 18463 27557 18475 27560
rect 18417 27551 18475 27557
rect 19886 27548 19892 27560
rect 19944 27548 19950 27600
rect 36541 27591 36599 27597
rect 36541 27557 36553 27591
rect 36587 27588 36599 27591
rect 37458 27588 37464 27600
rect 36587 27560 37464 27588
rect 36587 27557 36599 27560
rect 36541 27551 36599 27557
rect 37458 27548 37464 27560
rect 37516 27548 37522 27600
rect 43073 27591 43131 27597
rect 43073 27557 43085 27591
rect 43119 27588 43131 27591
rect 43533 27591 43591 27597
rect 43533 27588 43545 27591
rect 43119 27560 43545 27588
rect 43119 27557 43131 27560
rect 43073 27551 43131 27557
rect 43533 27557 43545 27560
rect 43579 27557 43591 27591
rect 45278 27588 45284 27600
rect 45239 27560 45284 27588
rect 43533 27551 43591 27557
rect 45278 27548 45284 27560
rect 45336 27548 45342 27600
rect 16942 27412 16948 27464
rect 17000 27452 17006 27464
rect 17310 27461 17316 27464
rect 17037 27455 17095 27461
rect 17037 27452 17049 27455
rect 17000 27424 17049 27452
rect 17000 27412 17006 27424
rect 17037 27421 17049 27424
rect 17083 27421 17095 27455
rect 17304 27452 17316 27461
rect 17271 27424 17316 27452
rect 17037 27415 17095 27421
rect 17304 27415 17316 27424
rect 17310 27412 17316 27415
rect 17368 27412 17374 27464
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 20990 27461 20996 27464
rect 20717 27455 20775 27461
rect 20717 27452 20729 27455
rect 20680 27424 20729 27452
rect 20680 27412 20686 27424
rect 20717 27421 20729 27424
rect 20763 27421 20775 27455
rect 20984 27452 20996 27461
rect 20951 27424 20996 27452
rect 20717 27415 20775 27421
rect 20984 27415 20996 27424
rect 20990 27412 20996 27415
rect 21048 27412 21054 27464
rect 23198 27452 23204 27464
rect 23159 27424 23204 27452
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 24029 27455 24087 27461
rect 24029 27421 24041 27455
rect 24075 27452 24087 27455
rect 25694 27455 25752 27461
rect 25694 27452 25706 27455
rect 24075 27424 25706 27452
rect 24075 27421 24087 27424
rect 24029 27415 24087 27421
rect 25694 27421 25706 27424
rect 25740 27421 25752 27455
rect 25694 27415 25752 27421
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27452 26019 27455
rect 27706 27452 27712 27464
rect 26007 27424 27712 27452
rect 26007 27421 26019 27424
rect 25961 27415 26019 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 31202 27452 31208 27464
rect 31163 27424 31208 27452
rect 31202 27412 31208 27424
rect 31260 27412 31266 27464
rect 31665 27455 31723 27461
rect 31665 27421 31677 27455
rect 31711 27452 31723 27455
rect 32306 27452 32312 27464
rect 31711 27424 32312 27452
rect 31711 27421 31723 27424
rect 31665 27415 31723 27421
rect 32306 27412 32312 27424
rect 32364 27412 32370 27464
rect 34514 27412 34520 27464
rect 34572 27452 34578 27464
rect 35434 27461 35440 27464
rect 35161 27455 35219 27461
rect 35161 27452 35173 27455
rect 34572 27424 35173 27452
rect 34572 27412 34578 27424
rect 35161 27421 35173 27424
rect 35207 27421 35219 27455
rect 35428 27452 35440 27461
rect 35395 27424 35440 27452
rect 35161 27415 35219 27421
rect 35428 27415 35440 27424
rect 35434 27412 35440 27415
rect 35492 27412 35498 27464
rect 36998 27452 37004 27464
rect 36959 27424 37004 27452
rect 36998 27412 37004 27424
rect 37056 27412 37062 27464
rect 38102 27452 38108 27464
rect 38063 27424 38108 27452
rect 38102 27412 38108 27424
rect 38160 27412 38166 27464
rect 40037 27455 40095 27461
rect 40037 27421 40049 27455
rect 40083 27452 40095 27455
rect 42058 27452 42064 27464
rect 40083 27424 42064 27452
rect 40083 27421 40095 27424
rect 40037 27415 40095 27421
rect 42058 27412 42064 27424
rect 42116 27412 42122 27464
rect 44910 27412 44916 27464
rect 44968 27452 44974 27464
rect 45189 27455 45247 27461
rect 45189 27452 45201 27455
rect 44968 27424 45201 27452
rect 44968 27412 44974 27424
rect 45189 27421 45201 27424
rect 45235 27421 45247 27455
rect 45370 27452 45376 27464
rect 45331 27424 45376 27452
rect 45189 27415 45247 27421
rect 45370 27412 45376 27424
rect 45428 27412 45434 27464
rect 27338 27344 27344 27396
rect 27396 27384 27402 27396
rect 31938 27393 31944 27396
rect 27954 27387 28012 27393
rect 27954 27384 27966 27387
rect 27396 27356 27966 27384
rect 27396 27344 27402 27356
rect 27954 27353 27966 27356
rect 28000 27353 28012 27387
rect 31932 27384 31944 27393
rect 31899 27356 31944 27384
rect 27954 27347 28012 27353
rect 31932 27347 31944 27356
rect 31938 27344 31944 27347
rect 31996 27344 32002 27396
rect 38372 27387 38430 27393
rect 38372 27353 38384 27387
rect 38418 27384 38430 27387
rect 40126 27384 40132 27396
rect 38418 27356 40132 27384
rect 38418 27353 38430 27356
rect 38372 27347 38430 27353
rect 40126 27344 40132 27356
rect 40184 27344 40190 27396
rect 40310 27393 40316 27396
rect 40304 27347 40316 27393
rect 40368 27384 40374 27396
rect 42705 27387 42763 27393
rect 40368 27356 40404 27384
rect 40310 27344 40316 27347
rect 40368 27344 40374 27356
rect 42705 27353 42717 27387
rect 42751 27384 42763 27387
rect 42794 27384 42800 27396
rect 42751 27356 42800 27384
rect 42751 27353 42763 27356
rect 42705 27347 42763 27353
rect 42794 27344 42800 27356
rect 42852 27344 42858 27396
rect 43714 27393 43720 27396
rect 43701 27387 43720 27393
rect 43701 27353 43713 27387
rect 43701 27347 43720 27353
rect 43714 27344 43720 27347
rect 43772 27344 43778 27396
rect 43898 27384 43904 27396
rect 43859 27356 43904 27384
rect 43898 27344 43904 27356
rect 43956 27344 43962 27396
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22278 27316 22284 27328
rect 22143 27288 22284 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 24581 27319 24639 27325
rect 24581 27285 24593 27319
rect 24627 27316 24639 27319
rect 25038 27316 25044 27328
rect 24627 27288 25044 27316
rect 24627 27285 24639 27288
rect 24581 27279 24639 27285
rect 25038 27276 25044 27288
rect 25096 27276 25102 27328
rect 29086 27316 29092 27328
rect 29047 27288 29092 27316
rect 29086 27276 29092 27288
rect 29144 27276 29150 27328
rect 33045 27319 33103 27325
rect 33045 27285 33057 27319
rect 33091 27316 33103 27319
rect 33410 27316 33416 27328
rect 33091 27288 33416 27316
rect 33091 27285 33103 27288
rect 33045 27279 33103 27285
rect 33410 27276 33416 27288
rect 33468 27276 33474 27328
rect 39482 27316 39488 27328
rect 39443 27288 39488 27316
rect 39482 27276 39488 27288
rect 39540 27276 39546 27328
rect 40494 27276 40500 27328
rect 40552 27316 40558 27328
rect 41417 27319 41475 27325
rect 41417 27316 41429 27319
rect 40552 27288 41429 27316
rect 40552 27276 40558 27288
rect 41417 27285 41429 27288
rect 41463 27285 41475 27319
rect 41417 27279 41475 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 18233 27115 18291 27121
rect 18233 27081 18245 27115
rect 18279 27112 18291 27115
rect 19334 27112 19340 27124
rect 18279 27084 19340 27112
rect 18279 27081 18291 27084
rect 18233 27075 18291 27081
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 31202 27072 31208 27124
rect 31260 27112 31266 27124
rect 36725 27115 36783 27121
rect 31260 27084 32444 27112
rect 31260 27072 31266 27084
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 17098 27047 17156 27053
rect 17098 27044 17110 27047
rect 16816 27016 17110 27044
rect 16816 27004 16822 27016
rect 17098 27013 17110 27016
rect 17144 27013 17156 27047
rect 17098 27007 17156 27013
rect 23008 27047 23066 27053
rect 23008 27013 23020 27047
rect 23054 27044 23066 27047
rect 23198 27044 23204 27056
rect 23054 27016 23204 27044
rect 23054 27013 23066 27016
rect 23008 27007 23066 27013
rect 23198 27004 23204 27016
rect 23256 27004 23262 27056
rect 24848 27047 24906 27053
rect 24848 27013 24860 27047
rect 24894 27044 24906 27047
rect 25590 27044 25596 27056
rect 24894 27016 25596 27044
rect 24894 27013 24906 27016
rect 24848 27007 24906 27013
rect 25590 27004 25596 27016
rect 25648 27004 25654 27056
rect 28230 27047 28288 27053
rect 28230 27044 28242 27047
rect 27540 27016 28242 27044
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26976 16911 26979
rect 16942 26976 16948 26988
rect 16899 26948 16948 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 27540 26985 27568 27016
rect 28230 27013 28242 27016
rect 28276 27013 28288 27047
rect 32306 27044 32312 27056
rect 28230 27007 28288 27013
rect 30392 27016 32312 27044
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 27706 26936 27712 26988
rect 27764 26976 27770 26988
rect 30392 26985 30420 27016
rect 32306 27004 32312 27016
rect 32364 27004 32370 27056
rect 32416 27044 32444 27084
rect 36725 27081 36737 27115
rect 36771 27112 36783 27115
rect 37734 27112 37740 27124
rect 36771 27084 37740 27112
rect 36771 27081 36783 27084
rect 36725 27075 36783 27081
rect 37734 27072 37740 27084
rect 37792 27072 37798 27124
rect 43898 27072 43904 27124
rect 43956 27112 43962 27124
rect 43993 27115 44051 27121
rect 43993 27112 44005 27115
rect 43956 27084 44005 27112
rect 43956 27072 43962 27084
rect 43993 27081 44005 27084
rect 44039 27081 44051 27115
rect 43993 27075 44051 27081
rect 32554 27047 32612 27053
rect 32554 27044 32566 27047
rect 32416 27016 32566 27044
rect 32554 27013 32566 27016
rect 32600 27013 32612 27047
rect 38102 27044 38108 27056
rect 32554 27007 32612 27013
rect 35360 27016 38108 27044
rect 27985 26979 28043 26985
rect 27985 26976 27997 26979
rect 27764 26948 27997 26976
rect 27764 26936 27770 26948
rect 27985 26945 27997 26948
rect 28031 26945 28043 26979
rect 27985 26939 28043 26945
rect 30377 26979 30435 26985
rect 30377 26945 30389 26979
rect 30423 26945 30435 26979
rect 30377 26939 30435 26945
rect 30644 26979 30702 26985
rect 30644 26945 30656 26979
rect 30690 26976 30702 26979
rect 32950 26976 32956 26988
rect 30690 26948 32956 26976
rect 30690 26945 30702 26948
rect 30644 26939 30702 26945
rect 32950 26936 32956 26948
rect 33008 26936 33014 26988
rect 35360 26985 35388 27016
rect 38102 27004 38108 27016
rect 38160 27044 38166 27056
rect 38654 27053 38660 27056
rect 38648 27044 38660 27053
rect 38160 27016 38424 27044
rect 38615 27016 38660 27044
rect 38160 27004 38166 27016
rect 35345 26979 35403 26985
rect 35345 26945 35357 26979
rect 35391 26945 35403 26979
rect 35345 26939 35403 26945
rect 35612 26979 35670 26985
rect 35612 26945 35624 26979
rect 35658 26976 35670 26979
rect 36998 26976 37004 26988
rect 35658 26948 37004 26976
rect 35658 26945 35670 26948
rect 35612 26939 35670 26945
rect 36998 26936 37004 26948
rect 37056 26936 37062 26988
rect 38396 26985 38424 27016
rect 38648 27007 38660 27016
rect 38654 27004 38660 27007
rect 38712 27004 38718 27056
rect 39482 27004 39488 27056
rect 39540 27044 39546 27056
rect 40221 27047 40279 27053
rect 40221 27044 40233 27047
rect 39540 27016 40233 27044
rect 39540 27004 39546 27016
rect 40221 27013 40233 27016
rect 40267 27013 40279 27047
rect 40221 27007 40279 27013
rect 40310 27004 40316 27056
rect 40368 27004 40374 27056
rect 43714 27004 43720 27056
rect 43772 27044 43778 27056
rect 44177 27047 44235 27053
rect 44177 27044 44189 27047
rect 43772 27016 44189 27044
rect 43772 27004 43778 27016
rect 44177 27013 44189 27016
rect 44223 27013 44235 27047
rect 44177 27007 44235 27013
rect 38381 26979 38439 26985
rect 38381 26945 38393 26979
rect 38427 26945 38439 26979
rect 40328 26976 40356 27004
rect 40494 26976 40500 26988
rect 38381 26939 38439 26945
rect 38488 26948 40356 26976
rect 40455 26948 40500 26976
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 22741 26911 22799 26917
rect 22741 26908 22753 26911
rect 20680 26880 22753 26908
rect 20680 26868 20686 26880
rect 22741 26877 22753 26880
rect 22787 26877 22799 26911
rect 24578 26908 24584 26920
rect 24539 26880 24584 26908
rect 22741 26871 22799 26877
rect 24578 26868 24584 26880
rect 24636 26868 24642 26920
rect 32306 26908 32312 26920
rect 32267 26880 32312 26908
rect 32306 26868 32312 26880
rect 32364 26868 32370 26920
rect 37921 26911 37979 26917
rect 37921 26877 37933 26911
rect 37967 26908 37979 26911
rect 38488 26908 38516 26948
rect 40494 26936 40500 26948
rect 40552 26936 40558 26988
rect 42889 26979 42947 26985
rect 42889 26976 42901 26979
rect 42812 26948 42901 26976
rect 37967 26880 38516 26908
rect 40313 26911 40371 26917
rect 37967 26877 37979 26880
rect 37921 26871 37979 26877
rect 40313 26877 40325 26911
rect 40359 26877 40371 26911
rect 40313 26871 40371 26877
rect 39761 26843 39819 26849
rect 39761 26809 39773 26843
rect 39807 26840 39819 26843
rect 40328 26840 40356 26871
rect 39807 26812 40356 26840
rect 42812 26840 42840 26948
rect 42889 26945 42901 26948
rect 42935 26945 42947 26979
rect 43070 26976 43076 26988
rect 43031 26948 43076 26976
rect 42889 26939 42947 26945
rect 43070 26936 43076 26948
rect 43128 26976 43134 26988
rect 44085 26979 44143 26985
rect 44085 26976 44097 26979
rect 43128 26948 44097 26976
rect 43128 26936 43134 26948
rect 44085 26945 44097 26948
rect 44131 26945 44143 26979
rect 58066 26976 58072 26988
rect 58027 26948 58072 26976
rect 44085 26939 44143 26945
rect 58066 26936 58072 26948
rect 58124 26936 58130 26988
rect 42978 26908 42984 26920
rect 42939 26880 42984 26908
rect 42978 26868 42984 26880
rect 43036 26868 43042 26920
rect 43165 26911 43223 26917
rect 43165 26877 43177 26911
rect 43211 26908 43223 26911
rect 43714 26908 43720 26920
rect 43211 26880 43720 26908
rect 43211 26877 43223 26880
rect 43165 26871 43223 26877
rect 43714 26868 43720 26880
rect 43772 26868 43778 26920
rect 43438 26840 43444 26852
rect 42812 26812 43444 26840
rect 39807 26809 39819 26812
rect 39761 26803 39819 26809
rect 43438 26800 43444 26812
rect 43496 26840 43502 26852
rect 43809 26843 43867 26849
rect 43809 26840 43821 26843
rect 43496 26812 43821 26840
rect 43496 26800 43502 26812
rect 43809 26809 43821 26812
rect 43855 26809 43867 26843
rect 43809 26803 43867 26809
rect 24121 26775 24179 26781
rect 24121 26741 24133 26775
rect 24167 26772 24179 26775
rect 24946 26772 24952 26784
rect 24167 26744 24952 26772
rect 24167 26741 24179 26744
rect 24121 26735 24179 26741
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 25314 26732 25320 26784
rect 25372 26772 25378 26784
rect 25961 26775 26019 26781
rect 25961 26772 25973 26775
rect 25372 26744 25973 26772
rect 25372 26732 25378 26744
rect 25961 26741 25973 26744
rect 26007 26741 26019 26775
rect 25961 26735 26019 26741
rect 26605 26775 26663 26781
rect 26605 26741 26617 26775
rect 26651 26772 26663 26775
rect 27890 26772 27896 26784
rect 26651 26744 27896 26772
rect 26651 26741 26663 26744
rect 26605 26735 26663 26741
rect 27890 26732 27896 26744
rect 27948 26732 27954 26784
rect 29365 26775 29423 26781
rect 29365 26741 29377 26775
rect 29411 26772 29423 26775
rect 29822 26772 29828 26784
rect 29411 26744 29828 26772
rect 29411 26741 29423 26744
rect 29365 26735 29423 26741
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 31757 26775 31815 26781
rect 31757 26741 31769 26775
rect 31803 26772 31815 26775
rect 33318 26772 33324 26784
rect 31803 26744 33324 26772
rect 31803 26741 31815 26744
rect 31757 26735 31815 26741
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 33594 26732 33600 26784
rect 33652 26772 33658 26784
rect 33689 26775 33747 26781
rect 33689 26772 33701 26775
rect 33652 26744 33701 26772
rect 33652 26732 33658 26744
rect 33689 26741 33701 26744
rect 33735 26741 33747 26775
rect 33689 26735 33747 26741
rect 40034 26732 40040 26784
rect 40092 26772 40098 26784
rect 40221 26775 40279 26781
rect 40221 26772 40233 26775
rect 40092 26744 40233 26772
rect 40092 26732 40098 26744
rect 40221 26741 40233 26744
rect 40267 26741 40279 26775
rect 40678 26772 40684 26784
rect 40639 26744 40684 26772
rect 40221 26735 40279 26741
rect 40678 26732 40684 26744
rect 40736 26732 40742 26784
rect 43346 26772 43352 26784
rect 43307 26744 43352 26772
rect 43346 26732 43352 26744
rect 43404 26732 43410 26784
rect 44358 26772 44364 26784
rect 44319 26744 44364 26772
rect 44358 26732 44364 26744
rect 44416 26732 44422 26784
rect 58250 26772 58256 26784
rect 58211 26744 58256 26772
rect 58250 26732 58256 26744
rect 58308 26732 58314 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 20622 26528 20628 26580
rect 20680 26568 20686 26580
rect 20717 26571 20775 26577
rect 20717 26568 20729 26571
rect 20680 26540 20729 26568
rect 20680 26528 20686 26540
rect 20717 26537 20729 26540
rect 20763 26537 20775 26571
rect 27338 26568 27344 26580
rect 27299 26540 27344 26568
rect 20717 26531 20775 26537
rect 27338 26528 27344 26540
rect 27396 26528 27402 26580
rect 38565 26571 38623 26577
rect 38565 26537 38577 26571
rect 38611 26568 38623 26571
rect 40678 26568 40684 26580
rect 38611 26540 40684 26568
rect 38611 26537 38623 26540
rect 38565 26531 38623 26537
rect 40678 26528 40684 26540
rect 40736 26528 40742 26580
rect 43162 26568 43168 26580
rect 41386 26540 43168 26568
rect 41386 26500 41414 26540
rect 43162 26528 43168 26540
rect 43220 26528 43226 26580
rect 43438 26568 43444 26580
rect 43399 26540 43444 26568
rect 43438 26528 43444 26540
rect 43496 26528 43502 26580
rect 44085 26571 44143 26577
rect 44085 26537 44097 26571
rect 44131 26568 44143 26571
rect 45554 26568 45560 26580
rect 44131 26540 45560 26568
rect 44131 26537 44143 26540
rect 44085 26531 44143 26537
rect 45554 26528 45560 26540
rect 45612 26528 45618 26580
rect 38856 26472 41414 26500
rect 24578 26432 24584 26444
rect 24539 26404 24584 26432
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 27706 26392 27712 26444
rect 27764 26432 27770 26444
rect 27801 26435 27859 26441
rect 27801 26432 27813 26435
rect 27764 26404 27813 26432
rect 27764 26392 27770 26404
rect 27801 26401 27813 26404
rect 27847 26401 27859 26435
rect 27801 26395 27859 26401
rect 37826 26392 37832 26444
rect 37884 26432 37890 26444
rect 38565 26435 38623 26441
rect 38565 26432 38577 26435
rect 37884 26404 38577 26432
rect 37884 26392 37890 26404
rect 38565 26401 38577 26404
rect 38611 26401 38623 26435
rect 38565 26395 38623 26401
rect 13538 26364 13544 26376
rect 13499 26336 13544 26364
rect 13538 26324 13544 26336
rect 13596 26324 13602 26376
rect 24854 26373 24860 26376
rect 24848 26364 24860 26373
rect 24815 26336 24860 26364
rect 24848 26327 24860 26336
rect 24854 26324 24860 26327
rect 24912 26324 24918 26376
rect 28068 26367 28126 26373
rect 28068 26333 28080 26367
rect 28114 26364 28126 26367
rect 28626 26364 28632 26376
rect 28114 26336 28632 26364
rect 28114 26333 28126 26336
rect 28068 26327 28126 26333
rect 28626 26324 28632 26336
rect 28684 26324 28690 26376
rect 30101 26367 30159 26373
rect 30101 26333 30113 26367
rect 30147 26364 30159 26367
rect 31754 26364 31760 26376
rect 30147 26336 31760 26364
rect 30147 26333 30159 26336
rect 30101 26327 30159 26333
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 31849 26367 31907 26373
rect 31849 26333 31861 26367
rect 31895 26364 31907 26367
rect 32306 26364 32312 26376
rect 31895 26336 32312 26364
rect 31895 26333 31907 26336
rect 31849 26327 31907 26333
rect 32306 26324 32312 26336
rect 32364 26364 32370 26376
rect 34514 26364 34520 26376
rect 32364 26336 34520 26364
rect 32364 26324 32370 26336
rect 34514 26324 34520 26336
rect 34572 26324 34578 26376
rect 37918 26324 37924 26376
rect 37976 26364 37982 26376
rect 38473 26367 38531 26373
rect 38473 26364 38485 26367
rect 37976 26336 38485 26364
rect 37976 26324 37982 26336
rect 38473 26333 38485 26336
rect 38519 26333 38531 26367
rect 38473 26327 38531 26333
rect 17954 26256 17960 26308
rect 18012 26296 18018 26308
rect 18877 26299 18935 26305
rect 18877 26296 18889 26299
rect 18012 26268 18889 26296
rect 18012 26256 18018 26268
rect 18877 26265 18889 26268
rect 18923 26296 18935 26299
rect 19429 26299 19487 26305
rect 19429 26296 19441 26299
rect 18923 26268 19441 26296
rect 18923 26265 18935 26268
rect 18877 26259 18935 26265
rect 19429 26265 19441 26268
rect 19475 26296 19487 26299
rect 23106 26296 23112 26308
rect 19475 26268 23112 26296
rect 19475 26265 19487 26268
rect 19429 26259 19487 26265
rect 23106 26256 23112 26268
rect 23164 26256 23170 26308
rect 32582 26305 32588 26308
rect 32576 26259 32588 26305
rect 32640 26296 32646 26308
rect 32640 26268 32676 26296
rect 32582 26256 32588 26259
rect 32640 26256 32646 26268
rect 13354 26228 13360 26240
rect 13315 26200 13360 26228
rect 13354 26188 13360 26200
rect 13412 26188 13418 26240
rect 25222 26188 25228 26240
rect 25280 26228 25286 26240
rect 25961 26231 26019 26237
rect 25961 26228 25973 26231
rect 25280 26200 25973 26228
rect 25280 26188 25286 26200
rect 25961 26197 25973 26200
rect 26007 26197 26019 26231
rect 25961 26191 26019 26197
rect 29181 26231 29239 26237
rect 29181 26197 29193 26231
rect 29227 26228 29239 26231
rect 30006 26228 30012 26240
rect 29227 26200 30012 26228
rect 29227 26197 29239 26200
rect 29181 26191 29239 26197
rect 30006 26188 30012 26200
rect 30064 26188 30070 26240
rect 33686 26228 33692 26240
rect 33647 26200 33692 26228
rect 33686 26188 33692 26200
rect 33744 26188 33750 26240
rect 38856 26237 38884 26472
rect 42058 26364 42064 26376
rect 41971 26336 42064 26364
rect 42058 26324 42064 26336
rect 42116 26364 42122 26376
rect 42702 26364 42708 26376
rect 42116 26336 42708 26364
rect 42116 26324 42122 26336
rect 42702 26324 42708 26336
rect 42760 26324 42766 26376
rect 43162 26324 43168 26376
rect 43220 26364 43226 26376
rect 43901 26367 43959 26373
rect 43901 26364 43913 26367
rect 43220 26336 43913 26364
rect 43220 26324 43226 26336
rect 43901 26333 43913 26336
rect 43947 26333 43959 26367
rect 43901 26327 43959 26333
rect 43990 26324 43996 26376
rect 44048 26364 44054 26376
rect 44048 26336 44093 26364
rect 44048 26324 44054 26336
rect 41874 26256 41880 26308
rect 41932 26296 41938 26308
rect 42306 26299 42364 26305
rect 42306 26296 42318 26299
rect 41932 26268 42318 26296
rect 41932 26256 41938 26268
rect 42306 26265 42318 26268
rect 42352 26265 42364 26299
rect 44174 26296 44180 26308
rect 44135 26268 44180 26296
rect 42306 26259 42364 26265
rect 44174 26256 44180 26268
rect 44232 26256 44238 26308
rect 38841 26231 38899 26237
rect 38841 26197 38853 26231
rect 38887 26197 38899 26231
rect 38841 26191 38899 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 24121 26027 24179 26033
rect 24121 25993 24133 26027
rect 24167 25993 24179 26027
rect 41874 26024 41880 26036
rect 41835 25996 41880 26024
rect 24121 25987 24179 25993
rect 13164 25959 13222 25965
rect 13164 25925 13176 25959
rect 13210 25956 13222 25959
rect 13354 25956 13360 25968
rect 13210 25928 13360 25956
rect 13210 25925 13222 25928
rect 13164 25919 13222 25925
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 24136 25956 24164 25987
rect 41874 25984 41880 25996
rect 41932 25984 41938 26036
rect 18892 25928 24164 25956
rect 18892 25897 18920 25928
rect 24946 25916 24952 25968
rect 25004 25956 25010 25968
rect 25041 25959 25099 25965
rect 25041 25956 25053 25959
rect 25004 25928 25053 25956
rect 25004 25916 25010 25928
rect 25041 25925 25053 25928
rect 25087 25925 25099 25959
rect 25041 25919 25099 25925
rect 27706 25916 27712 25968
rect 27764 25956 27770 25968
rect 29914 25956 29920 25968
rect 27764 25928 29920 25956
rect 27764 25916 27770 25928
rect 18877 25891 18935 25897
rect 18877 25857 18889 25891
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25888 19303 25891
rect 20346 25888 20352 25900
rect 19291 25860 20352 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 12897 25823 12955 25829
rect 12897 25789 12909 25823
rect 12943 25789 12955 25823
rect 12897 25783 12955 25789
rect 12912 25684 12940 25783
rect 15838 25780 15844 25832
rect 15896 25820 15902 25832
rect 18693 25823 18751 25829
rect 18693 25820 18705 25823
rect 15896 25792 18705 25820
rect 15896 25780 15902 25792
rect 18693 25789 18705 25792
rect 18739 25789 18751 25823
rect 19076 25820 19104 25851
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 22002 25888 22008 25900
rect 21963 25860 22008 25888
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22281 25891 22339 25897
rect 22281 25888 22293 25891
rect 22244 25860 22293 25888
rect 22244 25848 22250 25860
rect 22281 25857 22293 25860
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 24305 25891 24363 25897
rect 24305 25857 24317 25891
rect 24351 25888 24363 25891
rect 24581 25891 24639 25897
rect 24351 25860 24532 25888
rect 24351 25857 24363 25860
rect 24305 25851 24363 25857
rect 19334 25820 19340 25832
rect 19076 25792 19340 25820
rect 18693 25783 18751 25789
rect 19334 25780 19340 25792
rect 19392 25780 19398 25832
rect 22094 25820 22100 25832
rect 22055 25792 22100 25820
rect 22094 25780 22100 25792
rect 22152 25780 22158 25832
rect 24397 25823 24455 25829
rect 24397 25789 24409 25823
rect 24443 25789 24455 25823
rect 24397 25783 24455 25789
rect 22465 25755 22523 25761
rect 22465 25721 22477 25755
rect 22511 25752 22523 25755
rect 24412 25752 24440 25783
rect 22511 25724 24440 25752
rect 24504 25752 24532 25860
rect 24581 25857 24593 25891
rect 24627 25857 24639 25891
rect 24581 25851 24639 25857
rect 24596 25820 24624 25851
rect 24854 25848 24860 25900
rect 24912 25888 24918 25900
rect 25130 25888 25136 25900
rect 24912 25860 25136 25888
rect 24912 25848 24918 25860
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 25314 25888 25320 25900
rect 25275 25860 25320 25888
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 27816 25897 27844 25928
rect 29914 25916 29920 25928
rect 29972 25916 29978 25968
rect 33686 25956 33692 25968
rect 33647 25928 33692 25956
rect 33686 25916 33692 25928
rect 33744 25916 33750 25968
rect 42702 25916 42708 25968
rect 42760 25956 42766 25968
rect 45554 25965 45560 25968
rect 45548 25956 45560 25965
rect 42760 25928 45324 25956
rect 45515 25928 45560 25956
rect 42760 25916 42766 25928
rect 27801 25891 27859 25897
rect 27801 25857 27813 25891
rect 27847 25857 27859 25891
rect 27801 25851 27859 25857
rect 27890 25848 27896 25900
rect 27948 25888 27954 25900
rect 28057 25891 28115 25897
rect 28057 25888 28069 25891
rect 27948 25860 28069 25888
rect 27948 25848 27954 25860
rect 28057 25857 28069 25860
rect 28103 25857 28115 25891
rect 28057 25851 28115 25857
rect 29086 25848 29092 25900
rect 29144 25888 29150 25900
rect 29733 25891 29791 25897
rect 29733 25888 29745 25891
rect 29144 25860 29745 25888
rect 29144 25848 29150 25860
rect 29733 25857 29745 25860
rect 29779 25857 29791 25891
rect 30006 25888 30012 25900
rect 29967 25860 30012 25888
rect 29733 25851 29791 25857
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 32582 25888 32588 25900
rect 32539 25860 32588 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 32582 25848 32588 25860
rect 32640 25848 32646 25900
rect 33318 25848 33324 25900
rect 33376 25888 33382 25900
rect 33413 25891 33471 25897
rect 33413 25888 33425 25891
rect 33376 25860 33425 25888
rect 33376 25848 33382 25860
rect 33413 25857 33425 25860
rect 33459 25857 33471 25891
rect 42058 25888 42064 25900
rect 42019 25860 42064 25888
rect 33413 25851 33471 25857
rect 42058 25848 42064 25860
rect 42116 25848 42122 25900
rect 43438 25888 43444 25900
rect 43351 25860 43444 25888
rect 43438 25848 43444 25860
rect 43496 25888 43502 25900
rect 43990 25888 43996 25900
rect 43496 25860 43996 25888
rect 43496 25848 43502 25860
rect 43990 25848 43996 25860
rect 44048 25848 44054 25900
rect 44085 25891 44143 25897
rect 44085 25857 44097 25891
rect 44131 25888 44143 25891
rect 44174 25888 44180 25900
rect 44131 25860 44180 25888
rect 44131 25857 44143 25860
rect 44085 25851 44143 25857
rect 44174 25848 44180 25860
rect 44232 25848 44238 25900
rect 44358 25888 44364 25900
rect 44319 25860 44364 25888
rect 44358 25848 44364 25860
rect 44416 25848 44422 25900
rect 45296 25897 45324 25928
rect 45548 25919 45560 25928
rect 45554 25916 45560 25919
rect 45612 25916 45618 25968
rect 45281 25891 45339 25897
rect 45281 25857 45293 25891
rect 45327 25857 45339 25891
rect 45281 25851 45339 25857
rect 43168 25832 43220 25838
rect 24946 25820 24952 25832
rect 24596 25792 24952 25820
rect 24946 25780 24952 25792
rect 25004 25780 25010 25832
rect 25222 25820 25228 25832
rect 25183 25792 25228 25820
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 29822 25820 29828 25832
rect 29783 25792 29828 25820
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 33594 25820 33600 25832
rect 33555 25792 33600 25820
rect 33594 25780 33600 25792
rect 33652 25780 33658 25832
rect 43168 25774 43220 25780
rect 25501 25755 25559 25761
rect 25501 25752 25513 25755
rect 24504 25724 25513 25752
rect 22511 25721 22523 25724
rect 22465 25715 22523 25721
rect 25501 25721 25513 25724
rect 25547 25721 25559 25755
rect 25501 25715 25559 25721
rect 42886 25712 42892 25764
rect 42944 25752 42950 25764
rect 43073 25755 43131 25761
rect 43073 25752 43085 25755
rect 42944 25724 43085 25752
rect 42944 25712 42950 25724
rect 43073 25721 43085 25724
rect 43119 25721 43131 25755
rect 43073 25715 43131 25721
rect 13814 25684 13820 25696
rect 12912 25656 13820 25684
rect 13814 25644 13820 25656
rect 13872 25644 13878 25696
rect 13998 25644 14004 25696
rect 14056 25684 14062 25696
rect 14277 25687 14335 25693
rect 14277 25684 14289 25687
rect 14056 25656 14289 25684
rect 14056 25644 14062 25656
rect 14277 25653 14289 25656
rect 14323 25653 14335 25687
rect 17310 25684 17316 25696
rect 17271 25656 17316 25684
rect 14277 25647 14335 25653
rect 17310 25644 17316 25656
rect 17368 25644 17374 25696
rect 20717 25687 20775 25693
rect 20717 25653 20729 25687
rect 20763 25684 20775 25687
rect 20990 25684 20996 25696
rect 20763 25656 20996 25684
rect 20763 25653 20775 25656
rect 20717 25647 20775 25653
rect 20990 25644 20996 25656
rect 21048 25644 21054 25696
rect 21082 25644 21088 25696
rect 21140 25684 21146 25696
rect 21177 25687 21235 25693
rect 21177 25684 21189 25687
rect 21140 25656 21189 25684
rect 21140 25644 21146 25656
rect 21177 25653 21189 25656
rect 21223 25653 21235 25687
rect 22278 25684 22284 25696
rect 22239 25656 22284 25684
rect 21177 25647 21235 25653
rect 22278 25644 22284 25656
rect 22336 25644 22342 25696
rect 24581 25687 24639 25693
rect 24581 25653 24593 25687
rect 24627 25684 24639 25687
rect 24854 25684 24860 25696
rect 24627 25656 24860 25684
rect 24627 25653 24639 25656
rect 24581 25647 24639 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 25038 25684 25044 25696
rect 24999 25656 25044 25684
rect 25038 25644 25044 25656
rect 25096 25644 25102 25696
rect 29181 25687 29239 25693
rect 29181 25653 29193 25687
rect 29227 25684 29239 25687
rect 29733 25687 29791 25693
rect 29733 25684 29745 25687
rect 29227 25656 29745 25684
rect 29227 25653 29239 25656
rect 29181 25647 29239 25653
rect 29733 25653 29745 25656
rect 29779 25653 29791 25687
rect 29733 25647 29791 25653
rect 30193 25687 30251 25693
rect 30193 25653 30205 25687
rect 30239 25684 30251 25687
rect 31570 25684 31576 25696
rect 30239 25656 31576 25684
rect 30239 25653 30251 25656
rect 30193 25647 30251 25653
rect 31570 25644 31576 25656
rect 31628 25644 31634 25696
rect 31754 25684 31760 25696
rect 31715 25656 31760 25684
rect 31754 25644 31760 25656
rect 31812 25644 31818 25696
rect 33226 25684 33232 25696
rect 33187 25656 33232 25684
rect 33226 25644 33232 25656
rect 33284 25644 33290 25696
rect 33410 25684 33416 25696
rect 33371 25656 33416 25684
rect 33410 25644 33416 25656
rect 33468 25644 33474 25696
rect 40310 25684 40316 25696
rect 40271 25656 40316 25684
rect 40310 25644 40316 25656
rect 40368 25644 40374 25696
rect 46661 25687 46719 25693
rect 46661 25653 46673 25687
rect 46707 25684 46719 25687
rect 58066 25684 58072 25696
rect 46707 25656 58072 25684
rect 46707 25653 46719 25656
rect 46661 25647 46719 25653
rect 58066 25644 58072 25656
rect 58124 25644 58130 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 13265 25483 13323 25489
rect 13265 25449 13277 25483
rect 13311 25480 13323 25483
rect 13538 25480 13544 25492
rect 13311 25452 13544 25480
rect 13311 25449 13323 25452
rect 13265 25443 13323 25449
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 22186 25480 22192 25492
rect 22147 25452 22192 25480
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 33226 25480 33232 25492
rect 33187 25452 33232 25480
rect 33226 25440 33232 25452
rect 33284 25440 33290 25492
rect 44085 25483 44143 25489
rect 44085 25449 44097 25483
rect 44131 25480 44143 25483
rect 44174 25480 44180 25492
rect 44131 25452 44180 25480
rect 44131 25449 44143 25452
rect 44085 25443 44143 25449
rect 44174 25440 44180 25452
rect 44232 25440 44238 25492
rect 13446 25412 13452 25424
rect 13407 25384 13452 25412
rect 13446 25372 13452 25384
rect 13504 25372 13510 25424
rect 20622 25304 20628 25356
rect 20680 25344 20686 25356
rect 20809 25347 20867 25353
rect 20809 25344 20821 25347
rect 20680 25316 20821 25344
rect 20680 25304 20686 25316
rect 20809 25313 20821 25316
rect 20855 25313 20867 25347
rect 33134 25344 33140 25356
rect 33095 25316 33140 25344
rect 20809 25307 20867 25313
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 13725 25279 13783 25285
rect 13725 25245 13737 25279
rect 13771 25276 13783 25279
rect 13998 25276 14004 25288
rect 13771 25248 14004 25276
rect 13771 25245 13783 25248
rect 13725 25239 13783 25245
rect 13998 25236 14004 25248
rect 14056 25276 14062 25288
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 14056 25248 14473 25276
rect 14056 25236 14062 25248
rect 14461 25245 14473 25248
rect 14507 25245 14519 25279
rect 17034 25276 17040 25288
rect 16995 25248 17040 25276
rect 14461 25239 14519 25245
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 17310 25285 17316 25288
rect 17304 25276 17316 25285
rect 17271 25248 17316 25276
rect 17304 25239 17316 25248
rect 17310 25236 17316 25239
rect 17368 25236 17374 25288
rect 20346 25276 20352 25288
rect 20307 25248 20352 25276
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 21082 25285 21088 25288
rect 21076 25276 21088 25285
rect 21043 25248 21088 25276
rect 21076 25239 21088 25248
rect 21082 25236 21088 25239
rect 21140 25236 21146 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 24854 25276 24860 25288
rect 24811 25248 24860 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 30650 25276 30656 25288
rect 30611 25248 30656 25276
rect 30650 25236 30656 25248
rect 30708 25236 30714 25288
rect 31570 25236 31576 25288
rect 31628 25276 31634 25288
rect 33045 25279 33103 25285
rect 33045 25276 33057 25279
rect 31628 25248 33057 25276
rect 31628 25236 31634 25248
rect 33045 25245 33057 25248
rect 33091 25245 33103 25279
rect 33045 25239 33103 25245
rect 33321 25279 33379 25285
rect 33321 25245 33333 25279
rect 33367 25245 33379 25279
rect 33962 25276 33968 25288
rect 33923 25248 33968 25276
rect 33321 25239 33379 25245
rect 13906 25168 13912 25220
rect 13964 25208 13970 25220
rect 14277 25211 14335 25217
rect 14277 25208 14289 25211
rect 13964 25180 14289 25208
rect 13964 25168 13970 25180
rect 14277 25177 14289 25180
rect 14323 25177 14335 25211
rect 33336 25208 33364 25239
rect 33962 25236 33968 25248
rect 34020 25236 34026 25288
rect 36262 25276 36268 25288
rect 36223 25248 36268 25276
rect 36262 25236 36268 25248
rect 36320 25236 36326 25288
rect 36354 25236 36360 25288
rect 36412 25276 36418 25288
rect 36909 25279 36967 25285
rect 36909 25276 36921 25279
rect 36412 25248 36921 25276
rect 36412 25236 36418 25248
rect 36909 25245 36921 25248
rect 36955 25245 36967 25279
rect 38562 25276 38568 25288
rect 38523 25248 38568 25276
rect 36909 25239 36967 25245
rect 38562 25236 38568 25248
rect 38620 25236 38626 25288
rect 39485 25279 39543 25285
rect 39485 25245 39497 25279
rect 39531 25245 39543 25279
rect 40034 25276 40040 25288
rect 39995 25248 40040 25276
rect 39485 25239 39543 25245
rect 34698 25208 34704 25220
rect 33336 25180 34704 25208
rect 14277 25171 14335 25177
rect 34698 25168 34704 25180
rect 34756 25168 34762 25220
rect 39500 25208 39528 25239
rect 40034 25236 40040 25248
rect 40092 25236 40098 25288
rect 40310 25285 40316 25288
rect 40304 25276 40316 25285
rect 40271 25248 40316 25276
rect 40304 25239 40316 25248
rect 40310 25236 40316 25239
rect 40368 25236 40374 25288
rect 42702 25276 42708 25288
rect 42663 25248 42708 25276
rect 42702 25236 42708 25248
rect 42760 25236 42766 25288
rect 40218 25208 40224 25220
rect 39500 25180 40224 25208
rect 40218 25168 40224 25180
rect 40276 25168 40282 25220
rect 42972 25211 43030 25217
rect 42972 25177 42984 25211
rect 43018 25208 43030 25211
rect 43806 25208 43812 25220
rect 43018 25180 43812 25208
rect 43018 25177 43030 25180
rect 42972 25171 43030 25177
rect 43806 25168 43812 25180
rect 43864 25168 43870 25220
rect 14550 25100 14556 25152
rect 14608 25140 14614 25152
rect 14645 25143 14703 25149
rect 14645 25140 14657 25143
rect 14608 25112 14657 25140
rect 14608 25100 14614 25112
rect 14645 25109 14657 25112
rect 14691 25109 14703 25143
rect 14645 25103 14703 25109
rect 18417 25143 18475 25149
rect 18417 25109 18429 25143
rect 18463 25140 18475 25143
rect 18874 25140 18880 25152
rect 18463 25112 18880 25140
rect 18463 25109 18475 25112
rect 18417 25103 18475 25109
rect 18874 25100 18880 25112
rect 18932 25100 18938 25152
rect 33505 25143 33563 25149
rect 33505 25109 33517 25143
rect 33551 25140 33563 25143
rect 33870 25140 33876 25152
rect 33551 25112 33876 25140
rect 33551 25109 33563 25112
rect 33505 25103 33563 25109
rect 33870 25100 33876 25112
rect 33928 25100 33934 25152
rect 41417 25143 41475 25149
rect 41417 25109 41429 25143
rect 41463 25140 41475 25143
rect 41690 25140 41696 25152
rect 41463 25112 41696 25140
rect 41463 25109 41475 25112
rect 41417 25103 41475 25109
rect 41690 25100 41696 25112
rect 41748 25100 41754 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 13446 24896 13452 24948
rect 13504 24936 13510 24948
rect 13504 24908 14412 24936
rect 13504 24896 13510 24908
rect 13633 24871 13691 24877
rect 13633 24837 13645 24871
rect 13679 24868 13691 24871
rect 13998 24868 14004 24880
rect 13679 24840 14004 24868
rect 13679 24837 13691 24840
rect 13633 24831 13691 24837
rect 13998 24828 14004 24840
rect 14056 24828 14062 24880
rect 14384 24877 14412 24908
rect 14550 24896 14556 24948
rect 14608 24945 14614 24948
rect 14608 24939 14627 24945
rect 14615 24905 14627 24939
rect 14608 24899 14627 24905
rect 21453 24939 21511 24945
rect 21453 24905 21465 24939
rect 21499 24936 21511 24939
rect 22002 24936 22008 24948
rect 21499 24908 22008 24936
rect 21499 24905 21511 24908
rect 21453 24899 21511 24905
rect 14608 24896 14614 24899
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 42058 24896 42064 24948
rect 42116 24936 42122 24948
rect 42705 24939 42763 24945
rect 42705 24936 42717 24939
rect 42116 24908 42717 24936
rect 42116 24896 42122 24908
rect 42705 24905 42717 24908
rect 42751 24905 42763 24939
rect 42705 24899 42763 24905
rect 42886 24896 42892 24948
rect 42944 24936 42950 24948
rect 43806 24936 43812 24948
rect 42944 24908 43668 24936
rect 43767 24908 43812 24936
rect 42944 24896 42950 24908
rect 14369 24871 14427 24877
rect 14369 24837 14381 24871
rect 14415 24868 14427 24871
rect 15838 24868 15844 24880
rect 14415 24840 14504 24868
rect 14415 24837 14427 24840
rect 14369 24831 14427 24837
rect 12805 24803 12863 24809
rect 12805 24769 12817 24803
rect 12851 24800 12863 24803
rect 13170 24800 13176 24812
rect 12851 24772 13176 24800
rect 12851 24769 12863 24772
rect 12805 24763 12863 24769
rect 13170 24760 13176 24772
rect 13228 24760 13234 24812
rect 13538 24800 13544 24812
rect 13499 24772 13544 24800
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24800 13875 24803
rect 13906 24800 13912 24812
rect 13863 24772 13912 24800
rect 13863 24769 13875 24772
rect 13817 24763 13875 24769
rect 13906 24760 13912 24772
rect 13964 24760 13970 24812
rect 14476 24800 14504 24840
rect 14660 24840 15844 24868
rect 14660 24800 14688 24840
rect 15838 24828 15844 24840
rect 15896 24828 15902 24880
rect 17034 24828 17040 24880
rect 17092 24868 17098 24880
rect 20622 24868 20628 24880
rect 17092 24840 20628 24868
rect 17092 24828 17098 24840
rect 17604 24809 17632 24840
rect 20088 24809 20116 24840
rect 20622 24828 20628 24840
rect 20680 24828 20686 24880
rect 31754 24828 31760 24880
rect 31812 24868 31818 24880
rect 36078 24868 36084 24880
rect 31812 24840 36084 24868
rect 31812 24828 31818 24840
rect 36078 24828 36084 24840
rect 36136 24828 36142 24880
rect 38562 24877 38568 24880
rect 38556 24868 38568 24877
rect 38523 24840 38568 24868
rect 38556 24831 38568 24840
rect 38562 24828 38568 24831
rect 38620 24828 38626 24880
rect 40034 24828 40040 24880
rect 40092 24868 40098 24880
rect 41414 24868 41420 24880
rect 40092 24840 41420 24868
rect 40092 24828 40098 24840
rect 20346 24809 20352 24812
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 14476 24772 14688 24800
rect 14752 24772 15209 24800
rect 14752 24673 14780 24772
rect 15197 24769 15209 24772
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17856 24803 17914 24809
rect 17856 24769 17868 24803
rect 17902 24800 17914 24803
rect 19429 24803 19487 24809
rect 19429 24800 19441 24803
rect 17902 24772 19441 24800
rect 17902 24769 17914 24772
rect 17856 24763 17914 24769
rect 19429 24769 19441 24772
rect 19475 24769 19487 24803
rect 19429 24763 19487 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24769 20131 24803
rect 20340 24800 20352 24809
rect 20307 24772 20352 24800
rect 20073 24763 20131 24769
rect 20340 24763 20352 24772
rect 20346 24760 20352 24763
rect 20404 24760 20410 24812
rect 23106 24800 23112 24812
rect 23067 24772 23112 24800
rect 23106 24760 23112 24772
rect 23164 24800 23170 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23164 24772 23673 24800
rect 23164 24760 23170 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 29822 24760 29828 24812
rect 29880 24800 29886 24812
rect 30357 24803 30415 24809
rect 30357 24800 30369 24803
rect 29880 24772 30369 24800
rect 29880 24760 29886 24772
rect 30357 24769 30369 24772
rect 30403 24769 30415 24803
rect 30357 24763 30415 24769
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24800 33011 24803
rect 33669 24803 33727 24809
rect 33669 24800 33681 24803
rect 32999 24772 33681 24800
rect 32999 24769 33011 24772
rect 32953 24763 33011 24769
rect 33669 24769 33681 24772
rect 33715 24769 33727 24803
rect 33669 24763 33727 24769
rect 35796 24803 35854 24809
rect 35796 24769 35808 24803
rect 35842 24800 35854 24803
rect 36262 24800 36268 24812
rect 35842 24772 36268 24800
rect 35842 24769 35854 24772
rect 35796 24763 35854 24769
rect 36262 24760 36268 24772
rect 36320 24760 36326 24812
rect 36906 24760 36912 24812
rect 36964 24800 36970 24812
rect 37461 24803 37519 24809
rect 37461 24800 37473 24803
rect 36964 24772 37473 24800
rect 36964 24760 36970 24772
rect 37461 24769 37473 24772
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 38102 24760 38108 24812
rect 38160 24800 38166 24812
rect 40144 24809 40172 24840
rect 41414 24828 41420 24840
rect 41472 24828 41478 24880
rect 42978 24868 42984 24880
rect 42891 24840 42984 24868
rect 38289 24803 38347 24809
rect 38289 24800 38301 24803
rect 38160 24772 38301 24800
rect 38160 24760 38166 24772
rect 38289 24769 38301 24772
rect 38335 24769 38347 24803
rect 38289 24763 38347 24769
rect 40129 24803 40187 24809
rect 40129 24769 40141 24803
rect 40175 24769 40187 24803
rect 40129 24763 40187 24769
rect 40218 24760 40224 24812
rect 40276 24800 40282 24812
rect 42904 24809 42932 24840
rect 42978 24828 42984 24840
rect 43036 24868 43042 24880
rect 43438 24868 43444 24880
rect 43036 24840 43444 24868
rect 43036 24828 43042 24840
rect 43438 24828 43444 24840
rect 43496 24828 43502 24880
rect 40385 24803 40443 24809
rect 40385 24800 40397 24803
rect 40276 24772 40397 24800
rect 40276 24760 40282 24772
rect 40385 24769 40397 24772
rect 40431 24769 40443 24803
rect 40385 24763 40443 24769
rect 42889 24803 42947 24809
rect 42889 24769 42901 24803
rect 42935 24769 42947 24803
rect 43346 24800 43352 24812
rect 43307 24772 43352 24800
rect 42889 24763 42947 24769
rect 43346 24760 43352 24772
rect 43404 24760 43410 24812
rect 43640 24800 43668 24908
rect 43806 24896 43812 24908
rect 43864 24896 43870 24948
rect 43993 24803 44051 24809
rect 43993 24800 44005 24803
rect 43640 24772 44005 24800
rect 43993 24769 44005 24772
rect 44039 24769 44051 24803
rect 43993 24763 44051 24769
rect 44174 24760 44180 24812
rect 44232 24800 44238 24812
rect 44269 24803 44327 24809
rect 44269 24800 44281 24803
rect 44232 24772 44281 24800
rect 44232 24760 44238 24772
rect 44269 24769 44281 24772
rect 44315 24769 44327 24803
rect 44269 24763 44327 24769
rect 30101 24735 30159 24741
rect 30101 24701 30113 24735
rect 30147 24701 30159 24735
rect 30101 24695 30159 24701
rect 33413 24735 33471 24741
rect 33413 24701 33425 24735
rect 33459 24701 33471 24735
rect 33413 24695 33471 24701
rect 35529 24735 35587 24741
rect 35529 24701 35541 24735
rect 35575 24701 35587 24735
rect 35529 24695 35587 24701
rect 37553 24735 37611 24741
rect 37553 24701 37565 24735
rect 37599 24732 37611 24735
rect 38194 24732 38200 24744
rect 37599 24704 38200 24732
rect 37599 24701 37611 24704
rect 37553 24695 37611 24701
rect 14737 24667 14795 24673
rect 14737 24633 14749 24667
rect 14783 24633 14795 24667
rect 14737 24627 14795 24633
rect 24578 24624 24584 24676
rect 24636 24664 24642 24676
rect 24949 24667 25007 24673
rect 24949 24664 24961 24667
rect 24636 24636 24961 24664
rect 24636 24624 24642 24636
rect 24949 24633 24961 24636
rect 24995 24633 25007 24667
rect 24949 24627 25007 24633
rect 12986 24596 12992 24608
rect 12947 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 13412 24568 13553 24596
rect 13412 24556 13418 24568
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 14553 24599 14611 24605
rect 14553 24565 14565 24599
rect 14599 24596 14611 24599
rect 15194 24596 15200 24608
rect 14599 24568 15200 24596
rect 14599 24565 14611 24568
rect 14553 24559 14611 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 15378 24596 15384 24608
rect 15339 24568 15384 24596
rect 15378 24556 15384 24568
rect 15436 24556 15442 24608
rect 17126 24596 17132 24608
rect 17087 24568 17132 24596
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 18969 24599 19027 24605
rect 18969 24565 18981 24599
rect 19015 24596 19027 24599
rect 19150 24596 19156 24608
rect 19015 24568 19156 24596
rect 19015 24565 19027 24568
rect 18969 24559 19027 24565
rect 19150 24556 19156 24568
rect 19208 24556 19214 24608
rect 29638 24596 29644 24608
rect 29599 24568 29644 24596
rect 29638 24556 29644 24568
rect 29696 24556 29702 24608
rect 29914 24556 29920 24608
rect 29972 24596 29978 24608
rect 30116 24596 30144 24695
rect 33428 24664 33456 24695
rect 31036 24636 33456 24664
rect 31036 24596 31064 24636
rect 29972 24568 31064 24596
rect 31481 24599 31539 24605
rect 29972 24556 29978 24568
rect 31481 24565 31493 24599
rect 31527 24596 31539 24599
rect 31846 24596 31852 24608
rect 31527 24568 31852 24596
rect 31527 24565 31539 24568
rect 31481 24559 31539 24565
rect 31846 24556 31852 24568
rect 31904 24556 31910 24608
rect 33428 24596 33456 24636
rect 34514 24596 34520 24608
rect 33428 24568 34520 24596
rect 34514 24556 34520 24568
rect 34572 24556 34578 24608
rect 34790 24596 34796 24608
rect 34751 24568 34796 24596
rect 34790 24556 34796 24568
rect 34848 24556 34854 24608
rect 35544 24596 35572 24695
rect 38194 24692 38200 24704
rect 38252 24692 38258 24744
rect 43073 24735 43131 24741
rect 43073 24701 43085 24735
rect 43119 24701 43131 24735
rect 43073 24695 43131 24701
rect 37826 24664 37832 24676
rect 37787 24636 37832 24664
rect 37826 24624 37832 24636
rect 37884 24624 37890 24676
rect 43088 24664 43116 24695
rect 44177 24667 44235 24673
rect 44177 24664 44189 24667
rect 43088 24636 44189 24664
rect 44177 24633 44189 24636
rect 44223 24664 44235 24667
rect 44358 24664 44364 24676
rect 44223 24636 44364 24664
rect 44223 24633 44235 24636
rect 44177 24627 44235 24633
rect 44358 24624 44364 24636
rect 44416 24624 44422 24676
rect 35894 24596 35900 24608
rect 35544 24568 35900 24596
rect 35894 24556 35900 24568
rect 35952 24556 35958 24608
rect 36909 24599 36967 24605
rect 36909 24565 36921 24599
rect 36955 24596 36967 24599
rect 37461 24599 37519 24605
rect 37461 24596 37473 24599
rect 36955 24568 37473 24596
rect 36955 24565 36967 24568
rect 36909 24559 36967 24565
rect 37461 24565 37473 24568
rect 37507 24565 37519 24599
rect 37461 24559 37519 24565
rect 39669 24599 39727 24605
rect 39669 24565 39681 24599
rect 39715 24596 39727 24599
rect 40862 24596 40868 24608
rect 39715 24568 40868 24596
rect 39715 24565 39727 24568
rect 39669 24559 39727 24565
rect 40862 24556 40868 24568
rect 40920 24556 40926 24608
rect 41509 24599 41567 24605
rect 41509 24565 41521 24599
rect 41555 24596 41567 24599
rect 41598 24596 41604 24608
rect 41555 24568 41604 24596
rect 41555 24565 41567 24568
rect 41509 24559 41567 24565
rect 41598 24556 41604 24568
rect 41656 24556 41662 24608
rect 43162 24596 43168 24608
rect 43123 24568 43168 24596
rect 43162 24556 43168 24568
rect 43220 24556 43226 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 22094 24392 22100 24404
rect 22055 24364 22100 24392
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 31297 24395 31355 24401
rect 31297 24361 31309 24395
rect 31343 24392 31355 24395
rect 31757 24395 31815 24401
rect 31757 24392 31769 24395
rect 31343 24364 31769 24392
rect 31343 24361 31355 24364
rect 31297 24355 31355 24361
rect 31757 24361 31769 24364
rect 31803 24361 31815 24395
rect 31757 24355 31815 24361
rect 32217 24395 32275 24401
rect 32217 24361 32229 24395
rect 32263 24392 32275 24395
rect 33134 24392 33140 24404
rect 32263 24364 33140 24392
rect 32263 24361 32275 24364
rect 32217 24355 32275 24361
rect 33134 24352 33140 24364
rect 33192 24352 33198 24404
rect 34333 24395 34391 24401
rect 34333 24361 34345 24395
rect 34379 24392 34391 24395
rect 34885 24395 34943 24401
rect 34885 24392 34897 24395
rect 34379 24364 34897 24392
rect 34379 24361 34391 24364
rect 34333 24355 34391 24361
rect 34885 24361 34897 24364
rect 34931 24361 34943 24395
rect 34885 24355 34943 24361
rect 41414 24352 41420 24404
rect 41472 24392 41478 24404
rect 42702 24392 42708 24404
rect 41472 24364 42708 24392
rect 41472 24352 41478 24364
rect 42702 24352 42708 24364
rect 42760 24392 42766 24404
rect 42797 24395 42855 24401
rect 42797 24392 42809 24395
rect 42760 24364 42809 24392
rect 42760 24352 42766 24364
rect 42797 24361 42809 24364
rect 42843 24361 42855 24395
rect 42797 24355 42855 24361
rect 12529 24327 12587 24333
rect 12529 24293 12541 24327
rect 12575 24324 12587 24327
rect 13446 24324 13452 24336
rect 12575 24296 13452 24324
rect 12575 24293 12587 24296
rect 12529 24287 12587 24293
rect 13446 24284 13452 24296
rect 13504 24284 13510 24336
rect 34698 24284 34704 24336
rect 34756 24324 34762 24336
rect 35253 24327 35311 24333
rect 35253 24324 35265 24327
rect 34756 24296 35265 24324
rect 34756 24284 34762 24296
rect 35253 24293 35265 24296
rect 35299 24293 35311 24327
rect 35253 24287 35311 24293
rect 17034 24216 17040 24268
rect 17092 24256 17098 24268
rect 17313 24259 17371 24265
rect 17313 24256 17325 24259
rect 17092 24228 17325 24256
rect 17092 24216 17098 24228
rect 17313 24225 17325 24228
rect 17359 24225 17371 24259
rect 24578 24256 24584 24268
rect 17313 24219 17371 24225
rect 22940 24228 24584 24256
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 13449 24191 13507 24197
rect 13449 24188 13461 24191
rect 12124 24160 13461 24188
rect 12124 24148 12130 24160
rect 13449 24157 13461 24160
rect 13495 24188 13507 24191
rect 13538 24188 13544 24200
rect 13495 24160 13544 24188
rect 13495 24157 13507 24160
rect 13449 24151 13507 24157
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 12250 24080 12256 24132
rect 12308 24120 12314 24132
rect 12805 24123 12863 24129
rect 12805 24120 12817 24123
rect 12308 24092 12817 24120
rect 12308 24080 12314 24092
rect 12805 24089 12817 24092
rect 12851 24089 12863 24123
rect 13740 24120 13768 24151
rect 13814 24148 13820 24200
rect 13872 24188 13878 24200
rect 16022 24188 16028 24200
rect 13872 24160 16028 24188
rect 13872 24148 13878 24160
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 16850 24188 16856 24200
rect 16811 24160 16856 24188
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 17126 24148 17132 24200
rect 17184 24188 17190 24200
rect 17569 24191 17627 24197
rect 17569 24188 17581 24191
rect 17184 24160 17581 24188
rect 17184 24148 17190 24160
rect 17569 24157 17581 24160
rect 17615 24157 17627 24191
rect 17569 24151 17627 24157
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24188 20775 24191
rect 22940 24188 22968 24228
rect 24578 24216 24584 24228
rect 24636 24216 24642 24268
rect 29914 24256 29920 24268
rect 29875 24228 29920 24256
rect 29914 24216 29920 24228
rect 29972 24216 29978 24268
rect 31846 24256 31852 24268
rect 31807 24228 31852 24256
rect 31846 24216 31852 24228
rect 31904 24216 31910 24268
rect 34790 24216 34796 24268
rect 34848 24256 34854 24268
rect 34977 24259 35035 24265
rect 34977 24256 34989 24259
rect 34848 24228 34989 24256
rect 34848 24216 34854 24228
rect 34977 24225 34989 24228
rect 35023 24225 35035 24259
rect 34977 24219 35035 24225
rect 37829 24259 37887 24265
rect 37829 24225 37841 24259
rect 37875 24256 37887 24259
rect 38102 24256 38108 24268
rect 37875 24228 38108 24256
rect 37875 24225 37887 24228
rect 37829 24219 37887 24225
rect 38102 24216 38108 24228
rect 38160 24216 38166 24268
rect 20763 24160 22968 24188
rect 20763 24157 20775 24160
rect 20717 24151 20775 24157
rect 23014 24148 23020 24200
rect 23072 24188 23078 24200
rect 24026 24188 24032 24200
rect 23072 24160 23117 24188
rect 23987 24160 24032 24188
rect 23072 24148 23078 24160
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 29178 24188 29184 24200
rect 29139 24160 29184 24188
rect 29178 24148 29184 24160
rect 29236 24148 29242 24200
rect 29638 24148 29644 24200
rect 29696 24188 29702 24200
rect 30173 24191 30231 24197
rect 30173 24188 30185 24191
rect 29696 24160 30185 24188
rect 29696 24148 29702 24160
rect 30173 24157 30185 24160
rect 30219 24157 30231 24191
rect 30173 24151 30231 24157
rect 31662 24148 31668 24200
rect 31720 24188 31726 24200
rect 32033 24191 32091 24197
rect 32033 24188 32045 24191
rect 31720 24160 32045 24188
rect 31720 24148 31726 24160
rect 32033 24157 32045 24160
rect 32079 24157 32091 24191
rect 32950 24188 32956 24200
rect 32911 24160 32956 24188
rect 32033 24151 32091 24157
rect 32950 24148 32956 24160
rect 33008 24148 33014 24200
rect 33220 24191 33278 24197
rect 33220 24157 33232 24191
rect 33266 24188 33278 24191
rect 33962 24188 33968 24200
rect 33266 24160 33968 24188
rect 33266 24157 33278 24160
rect 33220 24151 33278 24157
rect 33962 24148 33968 24160
rect 34020 24148 34026 24200
rect 34606 24148 34612 24200
rect 34664 24188 34670 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34664 24160 34897 24188
rect 34664 24148 34670 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 13906 24120 13912 24132
rect 13740 24092 13912 24120
rect 12805 24083 12863 24089
rect 13906 24080 13912 24092
rect 13964 24120 13970 24132
rect 13964 24092 14688 24120
rect 13964 24080 13970 24092
rect 14660 24064 14688 24092
rect 15378 24080 15384 24132
rect 15436 24120 15442 24132
rect 15758 24123 15816 24129
rect 15758 24120 15770 24123
rect 15436 24092 15770 24120
rect 15436 24080 15442 24092
rect 15758 24089 15770 24092
rect 15804 24089 15816 24123
rect 15758 24083 15816 24089
rect 16206 24080 16212 24132
rect 16264 24120 16270 24132
rect 20990 24129 20996 24132
rect 20984 24120 20996 24129
rect 16264 24092 18920 24120
rect 20951 24092 20996 24120
rect 16264 24080 16270 24092
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 13262 24052 13268 24064
rect 13223 24024 13268 24052
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 13998 24052 14004 24064
rect 13679 24024 14004 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13998 24012 14004 24024
rect 14056 24052 14062 24064
rect 14458 24052 14464 24064
rect 14056 24024 14464 24052
rect 14056 24012 14062 24024
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 14642 24052 14648 24064
rect 14603 24024 14648 24052
rect 14642 24012 14648 24024
rect 14700 24012 14706 24064
rect 18690 24012 18696 24064
rect 18748 24052 18754 24064
rect 18892 24052 18920 24092
rect 20984 24083 20996 24092
rect 20990 24080 20996 24083
rect 21048 24080 21054 24132
rect 24670 24120 24676 24132
rect 21100 24092 24676 24120
rect 21100 24052 21128 24092
rect 24670 24080 24676 24092
rect 24728 24080 24734 24132
rect 24848 24123 24906 24129
rect 24848 24089 24860 24123
rect 24894 24089 24906 24123
rect 24848 24083 24906 24089
rect 31757 24123 31815 24129
rect 31757 24089 31769 24123
rect 31803 24120 31815 24123
rect 31846 24120 31852 24132
rect 31803 24092 31852 24120
rect 31803 24089 31815 24092
rect 31757 24083 31815 24089
rect 18748 24024 18793 24052
rect 18892 24024 21128 24052
rect 18748 24012 18754 24024
rect 23290 24012 23296 24064
rect 23348 24052 23354 24064
rect 24863 24052 24891 24083
rect 31846 24080 31852 24092
rect 31904 24080 31910 24132
rect 36078 24120 36084 24132
rect 35991 24092 36084 24120
rect 36078 24080 36084 24092
rect 36136 24080 36142 24132
rect 41509 24123 41567 24129
rect 41509 24120 41521 24123
rect 41156 24092 41521 24120
rect 23348 24024 24891 24052
rect 23348 24012 23354 24024
rect 25774 24012 25780 24064
rect 25832 24052 25838 24064
rect 25961 24055 26019 24061
rect 25961 24052 25973 24055
rect 25832 24024 25973 24052
rect 25832 24012 25838 24024
rect 25961 24021 25973 24024
rect 26007 24021 26019 24055
rect 36096 24052 36124 24080
rect 41156 24064 41184 24092
rect 41509 24089 41521 24092
rect 41555 24089 41567 24123
rect 41509 24083 41567 24089
rect 38381 24055 38439 24061
rect 38381 24052 38393 24055
rect 36096 24024 38393 24052
rect 25961 24015 26019 24021
rect 38381 24021 38393 24024
rect 38427 24052 38439 24055
rect 41049 24055 41107 24061
rect 41049 24052 41061 24055
rect 38427 24024 41061 24052
rect 38427 24021 38439 24024
rect 38381 24015 38439 24021
rect 41049 24021 41061 24024
rect 41095 24052 41107 24055
rect 41138 24052 41144 24064
rect 41095 24024 41144 24052
rect 41095 24021 41107 24024
rect 41049 24015 41107 24021
rect 41138 24012 41144 24024
rect 41196 24012 41202 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 18417 23851 18475 23857
rect 18417 23817 18429 23851
rect 18463 23817 18475 23851
rect 19334 23848 19340 23860
rect 19295 23820 19340 23848
rect 18417 23811 18475 23817
rect 12250 23780 12256 23792
rect 11900 23752 12256 23780
rect 11900 23721 11928 23752
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 14737 23783 14795 23789
rect 14737 23749 14749 23783
rect 14783 23780 14795 23783
rect 16206 23780 16212 23792
rect 14783 23752 16212 23780
rect 14783 23749 14795 23752
rect 14737 23743 14795 23749
rect 16206 23740 16212 23752
rect 16264 23740 16270 23792
rect 16850 23740 16856 23792
rect 16908 23780 16914 23792
rect 17282 23783 17340 23789
rect 17282 23780 17294 23783
rect 16908 23752 17294 23780
rect 16908 23740 16914 23752
rect 17282 23749 17294 23752
rect 17328 23749 17340 23783
rect 18432 23780 18460 23811
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 24946 23808 24952 23860
rect 25004 23848 25010 23860
rect 26053 23851 26111 23857
rect 26053 23848 26065 23851
rect 25004 23820 26065 23848
rect 25004 23808 25010 23820
rect 26053 23817 26065 23820
rect 26099 23817 26111 23851
rect 31662 23848 31668 23860
rect 31623 23820 31668 23848
rect 26053 23811 26111 23817
rect 31662 23808 31668 23820
rect 31720 23808 31726 23860
rect 34606 23848 34612 23860
rect 34567 23820 34612 23848
rect 34606 23808 34612 23820
rect 34664 23808 34670 23860
rect 36906 23848 36912 23860
rect 36867 23820 36912 23848
rect 36906 23808 36912 23820
rect 36964 23808 36970 23860
rect 38102 23808 38108 23860
rect 38160 23808 38166 23860
rect 38194 23808 38200 23860
rect 38252 23848 38258 23860
rect 39209 23851 39267 23857
rect 39209 23848 39221 23851
rect 38252 23820 39221 23848
rect 38252 23808 38258 23820
rect 39209 23817 39221 23820
rect 39255 23817 39267 23851
rect 42978 23848 42984 23860
rect 42939 23820 42984 23848
rect 39209 23811 39267 23817
rect 42978 23808 42984 23820
rect 43036 23808 43042 23860
rect 18877 23783 18935 23789
rect 18877 23780 18889 23783
rect 18432 23752 18889 23780
rect 17282 23743 17340 23749
rect 18877 23749 18889 23752
rect 18923 23749 18935 23783
rect 24578 23780 24584 23792
rect 18877 23743 18935 23749
rect 23768 23752 24584 23780
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23681 11943 23715
rect 12066 23712 12072 23724
rect 12027 23684 12072 23712
rect 11885 23675 11943 23681
rect 12066 23672 12072 23684
rect 12124 23672 12130 23724
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15470 23712 15476 23724
rect 15252 23684 15476 23712
rect 15252 23672 15258 23684
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 11977 23647 12035 23653
rect 11977 23613 11989 23647
rect 12023 23644 12035 23647
rect 15580 23644 15608 23675
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 15712 23684 15757 23712
rect 15712 23672 15718 23684
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 15896 23684 15941 23712
rect 15896 23672 15902 23684
rect 16022 23672 16028 23724
rect 16080 23712 16086 23724
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 16080 23684 17049 23712
rect 16080 23672 16086 23684
rect 17037 23681 17049 23684
rect 17083 23681 17095 23715
rect 19150 23712 19156 23724
rect 19111 23684 19156 23712
rect 17037 23675 17095 23681
rect 19150 23672 19156 23684
rect 19208 23672 19214 23724
rect 23290 23712 23296 23724
rect 23251 23684 23296 23712
rect 23290 23672 23296 23684
rect 23348 23672 23354 23724
rect 23768 23721 23796 23752
rect 24578 23740 24584 23752
rect 24636 23740 24642 23792
rect 30552 23783 30610 23789
rect 30552 23749 30564 23783
rect 30598 23780 30610 23783
rect 30650 23780 30656 23792
rect 30598 23752 30656 23780
rect 30598 23749 30610 23752
rect 30552 23743 30610 23749
rect 30650 23740 30656 23752
rect 30708 23740 30714 23792
rect 35894 23780 35900 23792
rect 33244 23752 35900 23780
rect 24026 23721 24032 23724
rect 23753 23715 23811 23721
rect 23753 23681 23765 23715
rect 23799 23681 23811 23715
rect 24020 23712 24032 23721
rect 23987 23684 24032 23712
rect 23753 23675 23811 23681
rect 24020 23675 24032 23684
rect 24026 23672 24032 23675
rect 24084 23672 24090 23724
rect 25590 23712 25596 23724
rect 25551 23684 25596 23712
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 25866 23712 25872 23724
rect 25827 23684 25872 23712
rect 25866 23672 25872 23684
rect 25924 23672 25930 23724
rect 29822 23712 29828 23724
rect 29783 23684 29828 23712
rect 29822 23672 29828 23684
rect 29880 23672 29886 23724
rect 29914 23672 29920 23724
rect 29972 23712 29978 23724
rect 30285 23715 30343 23721
rect 30285 23712 30297 23715
rect 29972 23684 30297 23712
rect 29972 23672 29978 23684
rect 30285 23681 30297 23684
rect 30331 23681 30343 23715
rect 30285 23675 30343 23681
rect 32950 23672 32956 23724
rect 33008 23712 33014 23724
rect 33244 23721 33272 23752
rect 33502 23721 33508 23724
rect 33229 23715 33287 23721
rect 33229 23712 33241 23715
rect 33008 23684 33241 23712
rect 33008 23672 33014 23684
rect 33229 23681 33241 23684
rect 33275 23681 33287 23715
rect 33229 23675 33287 23681
rect 33496 23675 33508 23721
rect 33560 23712 33566 23724
rect 35544 23721 35572 23752
rect 35894 23740 35900 23752
rect 35952 23780 35958 23792
rect 38120 23780 38148 23808
rect 35952 23752 38148 23780
rect 35952 23740 35958 23752
rect 35529 23715 35587 23721
rect 33560 23684 33596 23712
rect 33502 23672 33508 23675
rect 33560 23672 33566 23684
rect 35529 23681 35541 23715
rect 35575 23681 35587 23715
rect 35529 23675 35587 23681
rect 35796 23715 35854 23721
rect 35796 23681 35808 23715
rect 35842 23712 35854 23715
rect 36354 23712 36360 23724
rect 35842 23684 36360 23712
rect 35842 23681 35854 23684
rect 35796 23675 35854 23681
rect 36354 23672 36360 23684
rect 36412 23672 36418 23724
rect 37844 23721 37872 23752
rect 37829 23715 37887 23721
rect 37829 23681 37841 23715
rect 37875 23681 37887 23715
rect 37829 23675 37887 23681
rect 37918 23672 37924 23724
rect 37976 23712 37982 23724
rect 38085 23715 38143 23721
rect 38085 23712 38097 23715
rect 37976 23684 38097 23712
rect 37976 23672 37982 23684
rect 38085 23681 38097 23684
rect 38131 23681 38143 23715
rect 40034 23712 40040 23724
rect 39995 23684 40040 23712
rect 38085 23675 38143 23681
rect 40034 23672 40040 23684
rect 40092 23672 40098 23724
rect 40310 23721 40316 23724
rect 40304 23675 40316 23721
rect 40368 23712 40374 23724
rect 42610 23712 42616 23724
rect 40368 23684 40404 23712
rect 42571 23684 42616 23712
rect 40310 23672 40316 23675
rect 40368 23672 40374 23684
rect 42610 23672 42616 23684
rect 42668 23672 42674 23724
rect 42797 23715 42855 23721
rect 42797 23681 42809 23715
rect 42843 23712 42855 23715
rect 43622 23712 43628 23724
rect 42843 23684 43628 23712
rect 42843 23681 42855 23684
rect 42797 23675 42855 23681
rect 43622 23672 43628 23684
rect 43680 23672 43686 23724
rect 12023 23616 15608 23644
rect 12023 23613 12035 23616
rect 11977 23607 12035 23613
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 18748 23616 18981 23644
rect 18748 23604 18754 23616
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 25774 23644 25780 23656
rect 25735 23616 25780 23644
rect 18969 23607 19027 23613
rect 25774 23604 25780 23616
rect 25832 23604 25838 23656
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11112 23548 13492 23576
rect 11112 23536 11118 23548
rect 13464 23517 13492 23548
rect 13449 23511 13507 23517
rect 13449 23477 13461 23511
rect 13495 23508 13507 23511
rect 13998 23508 14004 23520
rect 13495 23480 14004 23508
rect 13495 23477 13507 23480
rect 13449 23471 13507 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15194 23508 15200 23520
rect 15155 23480 15200 23508
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 18874 23508 18880 23520
rect 18835 23480 18880 23508
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 25133 23511 25191 23517
rect 25133 23477 25145 23511
rect 25179 23508 25191 23511
rect 25593 23511 25651 23517
rect 25593 23508 25605 23511
rect 25179 23480 25605 23508
rect 25179 23477 25191 23480
rect 25133 23471 25191 23477
rect 25593 23477 25605 23480
rect 25639 23477 25651 23511
rect 25593 23471 25651 23477
rect 41417 23511 41475 23517
rect 41417 23477 41429 23511
rect 41463 23508 41475 23511
rect 41506 23508 41512 23520
rect 41463 23480 41512 23508
rect 41463 23477 41475 23480
rect 41417 23471 41475 23477
rect 41506 23468 41512 23480
rect 41564 23468 41570 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 12345 23307 12403 23313
rect 12345 23304 12357 23307
rect 12308 23276 12357 23304
rect 12308 23264 12314 23276
rect 12345 23273 12357 23276
rect 12391 23304 12403 23307
rect 14829 23307 14887 23313
rect 12391 23276 14412 23304
rect 12391 23273 12403 23276
rect 12345 23267 12403 23273
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 13814 23168 13820 23180
rect 13771 23140 13820 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 13814 23128 13820 23140
rect 13872 23128 13878 23180
rect 14384 23177 14412 23276
rect 14829 23273 14841 23307
rect 14875 23304 14887 23307
rect 15654 23304 15660 23316
rect 14875 23276 15660 23304
rect 14875 23273 14887 23276
rect 14829 23267 14887 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16206 23304 16212 23316
rect 16167 23276 16212 23304
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 24029 23307 24087 23313
rect 24029 23273 24041 23307
rect 24075 23304 24087 23307
rect 25590 23304 25596 23316
rect 24075 23276 25596 23304
rect 24075 23273 24087 23276
rect 24029 23267 24087 23273
rect 25590 23264 25596 23276
rect 25648 23264 25654 23316
rect 25866 23264 25872 23316
rect 25924 23304 25930 23316
rect 25961 23307 26019 23313
rect 25961 23304 25973 23307
rect 25924 23276 25973 23304
rect 25924 23264 25930 23276
rect 25961 23273 25973 23276
rect 26007 23273 26019 23307
rect 25961 23267 26019 23273
rect 31113 23307 31171 23313
rect 31113 23273 31125 23307
rect 31159 23304 31171 23307
rect 31846 23304 31852 23316
rect 31159 23276 31852 23304
rect 31159 23273 31171 23276
rect 31113 23267 31171 23273
rect 31846 23264 31852 23276
rect 31904 23264 31910 23316
rect 33502 23264 33508 23316
rect 33560 23304 33566 23316
rect 33597 23307 33655 23313
rect 33597 23304 33609 23307
rect 33560 23276 33609 23304
rect 33560 23264 33566 23276
rect 33597 23273 33609 23276
rect 33643 23273 33655 23307
rect 33597 23267 33655 23273
rect 36541 23307 36599 23313
rect 36541 23273 36553 23307
rect 36587 23304 36599 23307
rect 37918 23304 37924 23316
rect 36587 23276 37924 23304
rect 36587 23273 36599 23276
rect 36541 23267 36599 23273
rect 37918 23264 37924 23276
rect 37976 23264 37982 23316
rect 40221 23307 40279 23313
rect 40221 23273 40233 23307
rect 40267 23304 40279 23307
rect 40310 23304 40316 23316
rect 40267 23276 40316 23304
rect 40267 23273 40279 23276
rect 40221 23267 40279 23273
rect 40310 23264 40316 23276
rect 40368 23264 40374 23316
rect 41141 23307 41199 23313
rect 41141 23273 41153 23307
rect 41187 23304 41199 23307
rect 41506 23304 41512 23316
rect 41187 23276 41512 23304
rect 41187 23273 41199 23276
rect 41141 23267 41199 23273
rect 41506 23264 41512 23276
rect 41564 23264 41570 23316
rect 15470 23196 15476 23248
rect 15528 23236 15534 23248
rect 15565 23239 15623 23245
rect 15565 23236 15577 23239
rect 15528 23208 15577 23236
rect 15528 23196 15534 23208
rect 15565 23205 15577 23208
rect 15611 23205 15623 23239
rect 15565 23199 15623 23205
rect 41325 23239 41383 23245
rect 41325 23205 41337 23239
rect 41371 23236 41383 23239
rect 42610 23236 42616 23248
rect 41371 23208 42616 23236
rect 41371 23205 41383 23208
rect 41325 23199 41383 23205
rect 42610 23196 42616 23208
rect 42668 23196 42674 23248
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23137 14427 23171
rect 14642 23168 14648 23180
rect 14555 23140 14648 23168
rect 14369 23131 14427 23137
rect 14642 23128 14648 23140
rect 14700 23168 14706 23180
rect 24578 23168 24584 23180
rect 14700 23140 15700 23168
rect 24539 23140 24584 23168
rect 14700 23128 14706 23140
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23100 3111 23103
rect 12342 23100 12348 23112
rect 3099 23072 12348 23100
rect 3099 23069 3111 23072
rect 3053 23063 3111 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 13188 23072 14473 23100
rect 12066 22992 12072 23044
rect 12124 23032 12130 23044
rect 13188 23032 13216 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14550 23060 14556 23112
rect 14608 23100 14614 23112
rect 15672 23109 15700 23140
rect 24578 23128 24584 23140
rect 24636 23128 24642 23180
rect 41049 23171 41107 23177
rect 41049 23137 41061 23171
rect 41095 23168 41107 23171
rect 41598 23168 41604 23180
rect 41095 23140 41604 23168
rect 41095 23137 41107 23140
rect 41049 23131 41107 23137
rect 41598 23128 41604 23140
rect 41656 23128 41662 23180
rect 15473 23103 15531 23109
rect 15473 23100 15485 23103
rect 14608 23072 15485 23100
rect 14608 23060 14614 23072
rect 15473 23069 15485 23072
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 24596 23100 24624 23128
rect 24854 23109 24860 23112
rect 24848 23100 24860 23109
rect 22695 23072 24624 23100
rect 24815 23072 24860 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 24848 23063 24860 23072
rect 24854 23060 24860 23063
rect 24912 23060 24918 23112
rect 28902 23060 28908 23112
rect 28960 23100 28966 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 28960 23072 29745 23100
rect 28960 23060 28966 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 40862 23100 40868 23112
rect 40823 23072 40868 23100
rect 29733 23063 29791 23069
rect 40862 23060 40868 23072
rect 40920 23060 40926 23112
rect 41141 23103 41199 23109
rect 41141 23069 41153 23103
rect 41187 23100 41199 23103
rect 41690 23100 41696 23112
rect 41187 23072 41696 23100
rect 41187 23069 41199 23072
rect 41141 23063 41199 23069
rect 41690 23060 41696 23072
rect 41748 23060 41754 23112
rect 12124 23004 13216 23032
rect 13480 23035 13538 23041
rect 12124 22992 12130 23004
rect 13480 23001 13492 23035
rect 13526 23032 13538 23035
rect 15194 23032 15200 23044
rect 13526 23004 15200 23032
rect 13526 23001 13538 23004
rect 13480 22995 13538 23001
rect 15194 22992 15200 23004
rect 15252 22992 15258 23044
rect 22916 23035 22974 23041
rect 22916 23001 22928 23035
rect 22962 23032 22974 23035
rect 23014 23032 23020 23044
rect 22962 23004 23020 23032
rect 22962 23001 22974 23004
rect 22916 22995 22974 23001
rect 23014 22992 23020 23004
rect 23072 22992 23078 23044
rect 29178 22992 29184 23044
rect 29236 23032 29242 23044
rect 29978 23035 30036 23041
rect 29978 23032 29990 23035
rect 29236 23004 29990 23032
rect 29236 22992 29242 23004
rect 29978 23001 29990 23004
rect 30024 23001 30036 23035
rect 29978 22995 30036 23001
rect 2866 22964 2872 22976
rect 2827 22936 2872 22964
rect 2866 22924 2872 22936
rect 2924 22924 2930 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12161 22763 12219 22769
rect 12161 22760 12173 22763
rect 12124 22732 12173 22760
rect 12124 22720 12130 22732
rect 12161 22729 12173 22732
rect 12207 22729 12219 22763
rect 12161 22723 12219 22729
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 13872 22732 15301 22760
rect 13872 22720 13878 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 2716 22695 2774 22701
rect 2716 22661 2728 22695
rect 2762 22692 2774 22695
rect 2866 22692 2872 22704
rect 2762 22664 2872 22692
rect 2762 22661 2774 22664
rect 2716 22655 2774 22661
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13274 22695 13332 22701
rect 13274 22692 13286 22695
rect 13044 22664 13286 22692
rect 13044 22652 13050 22664
rect 13274 22661 13286 22664
rect 13320 22661 13332 22695
rect 13274 22655 13332 22661
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 13814 22624 13820 22636
rect 13587 22596 13820 22624
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 13998 22624 14004 22636
rect 13959 22596 14004 22624
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37608 22596 37841 22624
rect 37608 22584 37614 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 38013 22627 38071 22633
rect 38013 22593 38025 22627
rect 38059 22624 38071 22627
rect 38194 22624 38200 22636
rect 38059 22596 38200 22624
rect 38059 22593 38071 22596
rect 38013 22587 38071 22593
rect 38194 22584 38200 22596
rect 38252 22584 38258 22636
rect 2958 22556 2964 22568
rect 2919 22528 2964 22556
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16724 22392 16865 22420
rect 16724 22380 16730 22392
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 37918 22420 37924 22432
rect 37879 22392 37924 22420
rect 16853 22383 16911 22389
rect 37918 22380 37924 22392
rect 37976 22380 37982 22432
rect 41598 22420 41604 22432
rect 41559 22392 41604 22420
rect 41598 22380 41604 22392
rect 41656 22380 41662 22432
rect 42610 22420 42616 22432
rect 42571 22392 42616 22420
rect 42610 22380 42616 22392
rect 42668 22380 42674 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1762 22216 1768 22228
rect 1723 22188 1768 22216
rect 1762 22176 1768 22188
rect 1820 22176 1826 22228
rect 13354 22216 13360 22228
rect 13315 22188 13360 22216
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 40865 22219 40923 22225
rect 40865 22185 40877 22219
rect 40911 22216 40923 22219
rect 42705 22219 42763 22225
rect 40911 22188 42288 22216
rect 40911 22185 40923 22188
rect 40865 22179 40923 22185
rect 2866 22148 2872 22160
rect 2827 22120 2872 22148
rect 2866 22108 2872 22120
rect 2924 22108 2930 22160
rect 32858 22148 32864 22160
rect 32819 22120 32864 22148
rect 32858 22108 32864 22120
rect 32916 22108 32922 22160
rect 42260 22148 42288 22188
rect 42705 22185 42717 22219
rect 42751 22216 42763 22219
rect 43165 22219 43223 22225
rect 43165 22216 43177 22219
rect 42751 22188 43177 22216
rect 42751 22185 42763 22188
rect 42705 22179 42763 22185
rect 43165 22185 43177 22188
rect 43211 22185 43223 22219
rect 43165 22179 43223 22185
rect 42886 22148 42892 22160
rect 42260 22120 42892 22148
rect 42886 22108 42892 22120
rect 42944 22108 42950 22160
rect 35894 22040 35900 22092
rect 35952 22080 35958 22092
rect 36173 22083 36231 22089
rect 36173 22080 36185 22083
rect 35952 22052 36185 22080
rect 35952 22040 35958 22052
rect 36173 22049 36185 22052
rect 36219 22049 36231 22083
rect 36173 22043 36231 22049
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 13262 21972 13268 22024
rect 13320 21987 13326 22024
rect 16945 22015 17003 22021
rect 13320 21981 13369 21987
rect 13320 21972 13323 21981
rect 13289 21950 13323 21972
rect 13311 21947 13323 21950
rect 13357 21947 13369 21981
rect 16945 21981 16957 22015
rect 16991 22012 17003 22015
rect 17034 22012 17040 22024
rect 16991 21984 17040 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 17034 21972 17040 21984
rect 17092 21972 17098 22024
rect 17586 22012 17592 22024
rect 17547 21984 17592 22012
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 20346 22012 20352 22024
rect 20307 21984 20352 22012
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 20990 22012 20996 22024
rect 20951 21984 20996 22012
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 33870 22012 33876 22024
rect 33831 21984 33876 22012
rect 33870 21972 33876 21984
rect 33928 21972 33934 22024
rect 34054 22012 34060 22024
rect 34015 21984 34060 22012
rect 34054 21972 34060 21984
rect 34112 21972 34118 22024
rect 38838 22012 38844 22024
rect 38799 21984 38844 22012
rect 38838 21972 38844 21984
rect 38896 21972 38902 22024
rect 39022 22012 39028 22024
rect 38983 21984 39028 22012
rect 39022 21972 39028 21984
rect 39080 21972 39086 22024
rect 41325 22015 41383 22021
rect 41325 21981 41337 22015
rect 41371 22012 41383 22015
rect 41414 22012 41420 22024
rect 41371 21984 41420 22012
rect 41371 21981 41383 21984
rect 41325 21975 41383 21981
rect 41414 21972 41420 21984
rect 41472 21972 41478 22024
rect 41598 22021 41604 22024
rect 41592 22012 41604 22021
rect 41559 21984 41604 22012
rect 41592 21975 41604 21984
rect 41598 21972 41604 21975
rect 41656 21972 41662 22024
rect 43346 22012 43352 22024
rect 43307 21984 43352 22012
rect 43346 21972 43352 21984
rect 43404 21972 43410 22024
rect 43441 22015 43499 22021
rect 43441 21981 43453 22015
rect 43487 22012 43499 22015
rect 43714 22012 43720 22024
rect 43487 21984 43720 22012
rect 43487 21981 43499 21984
rect 43441 21975 43499 21981
rect 43714 21972 43720 21984
rect 43772 21972 43778 22024
rect 13311 21941 13369 21947
rect 13446 21904 13452 21956
rect 13504 21944 13510 21956
rect 13541 21947 13599 21953
rect 13541 21944 13553 21947
rect 13504 21916 13553 21944
rect 13504 21904 13510 21916
rect 13541 21913 13553 21916
rect 13587 21913 13599 21947
rect 13541 21907 13599 21913
rect 36440 21947 36498 21953
rect 36440 21913 36452 21947
rect 36486 21944 36498 21947
rect 36630 21944 36636 21956
rect 36486 21916 36636 21944
rect 36486 21913 36498 21916
rect 36440 21907 36498 21913
rect 36630 21904 36636 21916
rect 36688 21904 36694 21956
rect 38013 21947 38071 21953
rect 38013 21913 38025 21947
rect 38059 21913 38071 21947
rect 38194 21944 38200 21956
rect 38155 21916 38200 21944
rect 38013 21907 38071 21913
rect 4525 21879 4583 21885
rect 4525 21845 4537 21879
rect 4571 21876 4583 21879
rect 4614 21876 4620 21888
rect 4571 21848 4620 21876
rect 4571 21845 4583 21848
rect 4525 21839 4583 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 13170 21876 13176 21888
rect 13131 21848 13176 21876
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 14366 21876 14372 21888
rect 14327 21848 14372 21876
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 33965 21879 34023 21885
rect 33965 21845 33977 21879
rect 34011 21876 34023 21879
rect 37366 21876 37372 21888
rect 34011 21848 37372 21876
rect 34011 21845 34023 21848
rect 33965 21839 34023 21845
rect 37366 21836 37372 21848
rect 37424 21836 37430 21888
rect 37550 21876 37556 21888
rect 37511 21848 37556 21876
rect 37550 21836 37556 21848
rect 37608 21876 37614 21888
rect 38028 21876 38056 21907
rect 38194 21904 38200 21916
rect 38252 21904 38258 21956
rect 41874 21904 41880 21956
rect 41932 21944 41938 21956
rect 43165 21947 43223 21953
rect 43165 21944 43177 21947
rect 41932 21916 43177 21944
rect 41932 21904 41938 21916
rect 43165 21913 43177 21916
rect 43211 21913 43223 21947
rect 43165 21907 43223 21913
rect 38378 21876 38384 21888
rect 37608 21848 38056 21876
rect 38339 21848 38384 21876
rect 37608 21836 37614 21848
rect 38378 21836 38384 21848
rect 38436 21836 38442 21888
rect 39206 21876 39212 21888
rect 39167 21848 39212 21876
rect 39206 21836 39212 21848
rect 39264 21836 39270 21888
rect 43622 21876 43628 21888
rect 43583 21848 43628 21876
rect 43622 21836 43628 21848
rect 43680 21836 43686 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2590 21632 2596 21684
rect 2648 21672 2654 21684
rect 2869 21675 2927 21681
rect 2869 21672 2881 21675
rect 2648 21644 2881 21672
rect 2648 21632 2654 21644
rect 2869 21641 2881 21644
rect 2915 21672 2927 21675
rect 2958 21672 2964 21684
rect 2915 21644 2964 21672
rect 2915 21641 2927 21644
rect 2869 21635 2927 21641
rect 2958 21632 2964 21644
rect 3016 21632 3022 21684
rect 38194 21632 38200 21684
rect 38252 21672 38258 21684
rect 38841 21675 38899 21681
rect 38841 21672 38853 21675
rect 38252 21644 38853 21672
rect 38252 21632 38258 21644
rect 38841 21641 38853 21644
rect 38887 21641 38899 21675
rect 38841 21635 38899 21641
rect 43346 21632 43352 21684
rect 43404 21672 43410 21684
rect 43993 21675 44051 21681
rect 43993 21672 44005 21675
rect 43404 21644 44005 21672
rect 43404 21632 43410 21644
rect 43993 21641 44005 21644
rect 44039 21641 44051 21675
rect 43993 21635 44051 21641
rect 17120 21607 17178 21613
rect 17120 21573 17132 21607
rect 17166 21604 17178 21607
rect 17586 21604 17592 21616
rect 17166 21576 17592 21604
rect 17166 21573 17178 21576
rect 17120 21567 17178 21573
rect 17586 21564 17592 21576
rect 17644 21564 17650 21616
rect 20346 21613 20352 21616
rect 20340 21604 20352 21613
rect 20307 21576 20352 21604
rect 20340 21567 20352 21576
rect 20346 21564 20352 21567
rect 20404 21564 20410 21616
rect 35894 21604 35900 21616
rect 33428 21576 35900 21604
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21536 4399 21539
rect 4614 21536 4620 21548
rect 4387 21508 4620 21536
rect 4387 21505 4399 21508
rect 4341 21499 4399 21505
rect 4614 21496 4620 21508
rect 4672 21536 4678 21548
rect 13998 21536 14004 21548
rect 4672 21508 14004 21536
rect 4672 21496 4678 21508
rect 13998 21496 14004 21508
rect 14056 21536 14062 21548
rect 14366 21536 14372 21548
rect 14056 21508 14372 21536
rect 14056 21496 14062 21508
rect 14366 21496 14372 21508
rect 14424 21536 14430 21548
rect 14826 21536 14832 21548
rect 14424 21508 14832 21536
rect 14424 21496 14430 21508
rect 14826 21496 14832 21508
rect 14884 21496 14890 21548
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 16942 21536 16948 21548
rect 16899 21508 16948 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18104 21508 18705 21536
rect 18104 21496 18110 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 28445 21539 28503 21545
rect 28445 21505 28457 21539
rect 28491 21536 28503 21539
rect 29161 21539 29219 21545
rect 29161 21536 29173 21539
rect 28491 21508 29173 21536
rect 28491 21505 28503 21508
rect 28445 21499 28503 21505
rect 29161 21505 29173 21508
rect 29207 21505 29219 21539
rect 30742 21536 30748 21548
rect 30703 21508 30748 21536
rect 29161 21499 29219 21505
rect 18782 21468 18788 21480
rect 18743 21440 18788 21468
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 18233 21403 18291 21409
rect 18233 21369 18245 21403
rect 18279 21400 18291 21403
rect 18984 21400 19012 21499
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 31018 21536 31024 21548
rect 30979 21508 31024 21536
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 33428 21545 33456 21576
rect 35894 21564 35900 21576
rect 35952 21564 35958 21616
rect 36909 21607 36967 21613
rect 36909 21573 36921 21607
rect 36955 21604 36967 21607
rect 37550 21604 37556 21616
rect 36955 21576 37556 21604
rect 36955 21573 36967 21576
rect 36909 21567 36967 21573
rect 37550 21564 37556 21576
rect 37608 21564 37614 21616
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 33680 21539 33738 21545
rect 33680 21505 33692 21539
rect 33726 21536 33738 21539
rect 34146 21536 34152 21548
rect 33726 21508 34152 21536
rect 33726 21505 33738 21508
rect 33680 21499 33738 21505
rect 34146 21496 34152 21508
rect 34204 21496 34210 21548
rect 35434 21536 35440 21548
rect 35395 21508 35440 21536
rect 35434 21496 35440 21508
rect 35492 21496 35498 21548
rect 35526 21496 35532 21548
rect 35584 21536 35590 21548
rect 35713 21539 35771 21545
rect 35713 21536 35725 21539
rect 35584 21508 35725 21536
rect 35584 21496 35590 21508
rect 35713 21505 35725 21508
rect 35759 21505 35771 21539
rect 35912 21536 35940 21564
rect 37734 21545 37740 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 35912 21508 37473 21536
rect 35713 21499 35771 21505
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 37461 21499 37519 21505
rect 37728 21499 37740 21545
rect 37792 21536 37798 21548
rect 37792 21508 37828 21536
rect 37734 21496 37740 21499
rect 37792 21496 37798 21508
rect 39390 21496 39396 21548
rect 39448 21536 39454 21548
rect 40414 21539 40472 21545
rect 40414 21536 40426 21539
rect 39448 21508 40426 21536
rect 39448 21496 39454 21508
rect 40414 21505 40426 21508
rect 40460 21505 40472 21539
rect 40414 21499 40472 21505
rect 40681 21539 40739 21545
rect 40681 21505 40693 21539
rect 40727 21536 40739 21539
rect 41414 21536 41420 21548
rect 40727 21508 41420 21536
rect 40727 21505 40739 21508
rect 40681 21499 40739 21505
rect 41414 21496 41420 21508
rect 41472 21536 41478 21548
rect 42334 21536 42340 21548
rect 41472 21508 42340 21536
rect 41472 21496 41478 21508
rect 42334 21496 42340 21508
rect 42392 21536 42398 21548
rect 42886 21545 42892 21548
rect 42613 21539 42671 21545
rect 42613 21536 42625 21539
rect 42392 21508 42625 21536
rect 42392 21496 42398 21508
rect 42613 21505 42625 21508
rect 42659 21505 42671 21539
rect 42880 21536 42892 21545
rect 42847 21508 42892 21536
rect 42613 21499 42671 21505
rect 42880 21499 42892 21508
rect 42886 21496 42892 21499
rect 42944 21496 42950 21548
rect 20070 21468 20076 21480
rect 20031 21440 20076 21468
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 28902 21468 28908 21480
rect 28863 21440 28908 21468
rect 28902 21428 28908 21440
rect 28960 21428 28966 21480
rect 30834 21468 30840 21480
rect 30795 21440 30840 21468
rect 30834 21428 30840 21440
rect 30892 21428 30898 21480
rect 35621 21471 35679 21477
rect 35621 21437 35633 21471
rect 35667 21468 35679 21471
rect 36262 21468 36268 21480
rect 35667 21440 36268 21468
rect 35667 21437 35679 21440
rect 35621 21431 35679 21437
rect 36262 21428 36268 21440
rect 36320 21428 36326 21480
rect 18279 21372 19012 21400
rect 31205 21403 31263 21409
rect 18279 21369 18291 21372
rect 18233 21363 18291 21369
rect 31205 21369 31217 21403
rect 31251 21400 31263 21403
rect 33226 21400 33232 21412
rect 31251 21372 33232 21400
rect 31251 21369 31263 21372
rect 31205 21363 31263 21369
rect 33226 21360 33232 21372
rect 33284 21360 33290 21412
rect 34793 21403 34851 21409
rect 34793 21369 34805 21403
rect 34839 21400 34851 21403
rect 36633 21403 36691 21409
rect 34839 21372 35480 21400
rect 34839 21369 34851 21372
rect 34793 21363 34851 21369
rect 2133 21335 2191 21341
rect 2133 21301 2145 21335
rect 2179 21332 2191 21335
rect 2314 21332 2320 21344
rect 2179 21304 2320 21332
rect 2179 21301 2191 21304
rect 2133 21295 2191 21301
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 4985 21335 5043 21341
rect 4985 21301 4997 21335
rect 5031 21332 5043 21335
rect 5534 21332 5540 21344
rect 5031 21304 5540 21332
rect 5031 21301 5043 21304
rect 4985 21295 5043 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16574 21332 16580 21344
rect 16347 21304 16580 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 18690 21332 18696 21344
rect 18651 21304 18696 21332
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 19153 21335 19211 21341
rect 19153 21332 19165 21335
rect 19116 21304 19165 21332
rect 19116 21292 19122 21304
rect 19153 21301 19165 21304
rect 19199 21301 19211 21335
rect 21450 21332 21456 21344
rect 21411 21304 21456 21332
rect 19153 21295 19211 21301
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 22002 21332 22008 21344
rect 21963 21304 22008 21332
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 30285 21335 30343 21341
rect 30285 21301 30297 21335
rect 30331 21332 30343 21335
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30331 21304 30757 21332
rect 30331 21301 30343 21304
rect 30285 21295 30343 21301
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 31754 21332 31760 21344
rect 31715 21304 31760 21332
rect 30745 21295 30803 21301
rect 31754 21292 31760 21304
rect 31812 21292 31818 21344
rect 32493 21335 32551 21341
rect 32493 21301 32505 21335
rect 32539 21332 32551 21335
rect 32582 21332 32588 21344
rect 32539 21304 32588 21332
rect 32539 21301 32551 21304
rect 32493 21295 32551 21301
rect 32582 21292 32588 21304
rect 32640 21292 32646 21344
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 35452 21341 35480 21372
rect 36633 21369 36645 21403
rect 36679 21400 36691 21403
rect 37366 21400 37372 21412
rect 36679 21372 37372 21400
rect 36679 21369 36691 21372
rect 36633 21363 36691 21369
rect 37366 21360 37372 21372
rect 37424 21360 37430 21412
rect 35253 21335 35311 21341
rect 35253 21332 35265 21335
rect 34572 21304 35265 21332
rect 34572 21292 34578 21304
rect 35253 21301 35265 21304
rect 35299 21301 35311 21335
rect 35253 21295 35311 21301
rect 35437 21335 35495 21341
rect 35437 21301 35449 21335
rect 35483 21301 35495 21335
rect 35437 21295 35495 21301
rect 36449 21335 36507 21341
rect 36449 21301 36461 21335
rect 36495 21332 36507 21335
rect 36814 21332 36820 21344
rect 36495 21304 36820 21332
rect 36495 21301 36507 21304
rect 36449 21295 36507 21301
rect 36814 21292 36820 21304
rect 36872 21292 36878 21344
rect 39114 21292 39120 21344
rect 39172 21332 39178 21344
rect 39301 21335 39359 21341
rect 39301 21332 39313 21335
rect 39172 21304 39313 21332
rect 39172 21292 39178 21304
rect 39301 21301 39313 21304
rect 39347 21301 39359 21335
rect 39301 21295 39359 21301
rect 40770 21292 40776 21344
rect 40828 21332 40834 21344
rect 41141 21335 41199 21341
rect 41141 21332 41153 21335
rect 40828 21304 41153 21332
rect 40828 21292 40834 21304
rect 41141 21301 41153 21304
rect 41187 21301 41199 21335
rect 41141 21295 41199 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 3970 21128 3976 21140
rect 3931 21100 3976 21128
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 18049 21131 18107 21137
rect 18049 21097 18061 21131
rect 18095 21128 18107 21131
rect 18690 21128 18696 21140
rect 18095 21100 18696 21128
rect 18095 21097 18107 21100
rect 18049 21091 18107 21097
rect 18690 21088 18696 21100
rect 18748 21088 18754 21140
rect 21450 21088 21456 21140
rect 21508 21128 21514 21140
rect 22097 21131 22155 21137
rect 22097 21128 22109 21131
rect 21508 21100 22109 21128
rect 21508 21088 21514 21100
rect 22097 21097 22109 21100
rect 22143 21097 22155 21131
rect 22097 21091 22155 21097
rect 29181 21131 29239 21137
rect 29181 21097 29193 21131
rect 29227 21128 29239 21131
rect 30834 21128 30840 21140
rect 29227 21100 30840 21128
rect 29227 21097 29239 21100
rect 29181 21091 29239 21097
rect 30834 21088 30840 21100
rect 30892 21088 30898 21140
rect 34146 21128 34152 21140
rect 34107 21100 34152 21128
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 36262 21128 36268 21140
rect 36223 21100 36268 21128
rect 36262 21088 36268 21100
rect 36320 21088 36326 21140
rect 37553 21131 37611 21137
rect 37553 21097 37565 21131
rect 37599 21128 37611 21131
rect 38378 21128 38384 21140
rect 37599 21100 38384 21128
rect 37599 21097 37611 21100
rect 37553 21091 37611 21097
rect 38378 21088 38384 21100
rect 38436 21088 38442 21140
rect 38657 21131 38715 21137
rect 38657 21097 38669 21131
rect 38703 21128 38715 21131
rect 39022 21128 39028 21140
rect 38703 21100 39028 21128
rect 38703 21097 38715 21100
rect 38657 21091 38715 21097
rect 39022 21088 39028 21100
rect 39080 21088 39086 21140
rect 39390 21128 39396 21140
rect 39351 21100 39396 21128
rect 39390 21088 39396 21100
rect 39448 21088 39454 21140
rect 41414 21128 41420 21140
rect 40512 21100 41420 21128
rect 3421 21063 3479 21069
rect 3421 21029 3433 21063
rect 3467 21060 3479 21063
rect 21637 21063 21695 21069
rect 3467 21032 4108 21060
rect 3467 21029 3479 21032
rect 3421 21023 3479 21029
rect 4080 21001 4108 21032
rect 21637 21029 21649 21063
rect 21683 21060 21695 21063
rect 37366 21060 37372 21072
rect 21683 21032 22232 21060
rect 37279 21032 37372 21060
rect 21683 21029 21695 21032
rect 21637 21023 21695 21029
rect 22204 21001 22232 21032
rect 37366 21020 37372 21032
rect 37424 21060 37430 21072
rect 38838 21060 38844 21072
rect 37424 21032 38844 21060
rect 37424 21020 37430 21032
rect 38838 21020 38844 21032
rect 38896 21020 38902 21072
rect 4065 20995 4123 21001
rect 4065 20961 4077 20995
rect 4111 20961 4123 20995
rect 4065 20955 4123 20961
rect 22189 20995 22247 21001
rect 22189 20961 22201 20995
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2590 20924 2596 20936
rect 2087 20896 2596 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 4246 20924 4252 20936
rect 4207 20896 4252 20924
rect 4246 20884 4252 20896
rect 4304 20884 4310 20936
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20924 13599 20927
rect 13630 20924 13636 20936
rect 13587 20896 13636 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 13630 20884 13636 20896
rect 13688 20884 13694 20936
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 13964 20896 14289 20924
rect 13964 20884 13970 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20924 16727 20927
rect 16758 20924 16764 20936
rect 16715 20896 16764 20924
rect 16715 20893 16727 20896
rect 16669 20887 16727 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 19978 20924 19984 20936
rect 19843 20896 19984 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20070 20884 20076 20936
rect 20128 20924 20134 20936
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 20128 20896 20269 20924
rect 20128 20884 20134 20896
rect 20257 20893 20269 20896
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20524 20927 20582 20933
rect 20524 20893 20536 20927
rect 20570 20924 20582 20927
rect 20990 20924 20996 20936
rect 20570 20896 20996 20924
rect 20570 20893 20582 20896
rect 20524 20887 20582 20893
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 22370 20924 22376 20936
rect 22331 20896 22376 20924
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20924 27859 20927
rect 27890 20924 27896 20936
rect 27847 20896 27896 20924
rect 27847 20893 27859 20896
rect 27801 20887 27859 20893
rect 27890 20884 27896 20896
rect 27948 20924 27954 20936
rect 28902 20924 28908 20936
rect 27948 20896 28908 20924
rect 27948 20884 27954 20896
rect 28902 20884 28908 20896
rect 28960 20924 28966 20936
rect 29914 20924 29920 20936
rect 28960 20896 29920 20924
rect 28960 20884 28966 20896
rect 29914 20884 29920 20896
rect 29972 20924 29978 20936
rect 31849 20927 31907 20933
rect 31849 20924 31861 20927
rect 29972 20896 31861 20924
rect 29972 20884 29978 20896
rect 31849 20893 31861 20896
rect 31895 20924 31907 20927
rect 32306 20924 32312 20936
rect 31895 20896 32312 20924
rect 31895 20893 31907 20896
rect 31849 20887 31907 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 32582 20933 32588 20936
rect 32576 20924 32588 20933
rect 32543 20896 32588 20924
rect 32576 20887 32588 20896
rect 32582 20884 32588 20887
rect 32640 20884 32646 20936
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20924 34943 20927
rect 35894 20924 35900 20936
rect 34931 20896 35900 20924
rect 34931 20893 34943 20896
rect 34885 20887 34943 20893
rect 35894 20884 35900 20896
rect 35952 20884 35958 20936
rect 36722 20924 36728 20936
rect 36683 20896 36728 20924
rect 36722 20884 36728 20896
rect 36780 20884 36786 20936
rect 2130 20816 2136 20868
rect 2188 20856 2194 20868
rect 2286 20859 2344 20865
rect 2286 20856 2298 20859
rect 2188 20828 2298 20856
rect 2188 20816 2194 20828
rect 2286 20825 2298 20828
rect 2332 20825 2344 20859
rect 2286 20819 2344 20825
rect 3418 20816 3424 20868
rect 3476 20856 3482 20868
rect 3973 20859 4031 20865
rect 3973 20856 3985 20859
rect 3476 20828 3985 20856
rect 3476 20816 3482 20828
rect 3973 20825 3985 20828
rect 4019 20825 4031 20859
rect 3973 20819 4031 20825
rect 16936 20859 16994 20865
rect 16936 20825 16948 20859
rect 16982 20856 16994 20859
rect 17034 20856 17040 20868
rect 16982 20828 17040 20856
rect 16982 20825 16994 20828
rect 16936 20819 16994 20825
rect 17034 20816 17040 20828
rect 17092 20816 17098 20868
rect 22094 20856 22100 20868
rect 22055 20828 22100 20856
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 28068 20859 28126 20865
rect 28068 20825 28080 20859
rect 28114 20825 28126 20859
rect 28068 20819 28126 20825
rect 30101 20859 30159 20865
rect 30101 20825 30113 20859
rect 30147 20856 30159 20859
rect 31754 20856 31760 20868
rect 30147 20828 31760 20856
rect 30147 20825 30159 20828
rect 30101 20819 30159 20825
rect 4433 20791 4491 20797
rect 4433 20757 4445 20791
rect 4479 20788 4491 20791
rect 4706 20788 4712 20800
rect 4479 20760 4712 20788
rect 4479 20757 4491 20760
rect 4433 20751 4491 20757
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 22554 20788 22560 20800
rect 22515 20760 22560 20788
rect 22554 20748 22560 20760
rect 22612 20748 22618 20800
rect 28083 20788 28111 20819
rect 31754 20816 31760 20828
rect 31812 20816 31818 20868
rect 35152 20859 35210 20865
rect 35152 20825 35164 20859
rect 35198 20856 35210 20859
rect 35342 20856 35348 20868
rect 35198 20828 35348 20856
rect 35198 20825 35210 20828
rect 35152 20819 35210 20825
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 37384 20865 37412 21020
rect 37918 20952 37924 21004
rect 37976 20992 37982 21004
rect 38289 20995 38347 21001
rect 38289 20992 38301 20995
rect 37976 20964 38301 20992
rect 37976 20952 37982 20964
rect 38289 20961 38301 20964
rect 38335 20961 38347 20995
rect 39114 20992 39120 21004
rect 38289 20955 38347 20961
rect 38396 20964 39120 20992
rect 37369 20859 37427 20865
rect 37369 20825 37381 20859
rect 37415 20825 37427 20859
rect 37369 20819 37427 20825
rect 37585 20859 37643 20865
rect 37585 20825 37597 20859
rect 37631 20856 37643 20859
rect 37936 20856 37964 20952
rect 38396 20933 38424 20964
rect 39114 20952 39120 20964
rect 39172 20952 39178 21004
rect 40512 21001 40540 21100
rect 41414 21088 41420 21100
rect 41472 21088 41478 21140
rect 41874 21128 41880 21140
rect 41835 21100 41880 21128
rect 41874 21088 41880 21100
rect 41932 21088 41938 21140
rect 43714 21128 43720 21140
rect 43675 21100 43720 21128
rect 43714 21088 43720 21100
rect 43772 21088 43778 21140
rect 40497 20995 40555 21001
rect 40497 20961 40509 20995
rect 40543 20961 40555 20995
rect 42334 20992 42340 21004
rect 42295 20964 42340 20992
rect 40497 20955 40555 20961
rect 42334 20952 42340 20964
rect 42392 20952 42398 21004
rect 38381 20927 38439 20933
rect 38381 20893 38393 20927
rect 38427 20893 38439 20927
rect 39206 20924 39212 20936
rect 39167 20896 39212 20924
rect 38381 20887 38439 20893
rect 39206 20884 39212 20896
rect 39264 20884 39270 20936
rect 40770 20933 40776 20936
rect 40764 20924 40776 20933
rect 40731 20896 40776 20924
rect 40764 20887 40776 20896
rect 40770 20884 40776 20887
rect 40828 20884 40834 20936
rect 42610 20933 42616 20936
rect 42604 20924 42616 20933
rect 42571 20896 42616 20924
rect 42604 20887 42616 20896
rect 42610 20884 42616 20887
rect 42668 20884 42674 20936
rect 37631 20828 37964 20856
rect 37631 20825 37643 20828
rect 37585 20819 37643 20825
rect 30466 20788 30472 20800
rect 28083 20760 30472 20788
rect 30466 20748 30472 20760
rect 30524 20748 30530 20800
rect 33502 20748 33508 20800
rect 33560 20788 33566 20800
rect 33689 20791 33747 20797
rect 33689 20788 33701 20791
rect 33560 20760 33701 20788
rect 33560 20748 33566 20760
rect 33689 20757 33701 20760
rect 33735 20757 33747 20791
rect 33689 20751 33747 20757
rect 37737 20791 37795 20797
rect 37737 20757 37749 20791
rect 37783 20788 37795 20791
rect 37918 20788 37924 20800
rect 37783 20760 37924 20788
rect 37783 20757 37795 20760
rect 37737 20751 37795 20757
rect 37918 20748 37924 20760
rect 37976 20748 37982 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 3970 20584 3976 20596
rect 3931 20556 3976 20584
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 4433 20587 4491 20593
rect 4433 20584 4445 20587
rect 4304 20556 4445 20584
rect 4304 20544 4310 20556
rect 4433 20553 4445 20556
rect 4479 20553 4491 20587
rect 4433 20547 4491 20553
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20584 15715 20587
rect 21453 20587 21511 20593
rect 15703 20556 18828 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 2866 20525 2872 20528
rect 2860 20516 2872 20525
rect 2827 20488 2872 20516
rect 2860 20479 2872 20488
rect 2866 20476 2872 20479
rect 2924 20476 2930 20528
rect 5534 20476 5540 20528
rect 5592 20525 5598 20528
rect 5592 20516 5604 20525
rect 13814 20516 13820 20528
rect 5592 20488 5637 20516
rect 13372 20488 13820 20516
rect 5592 20479 5604 20488
rect 5592 20476 5598 20479
rect 2130 20448 2136 20460
rect 2091 20420 2136 20448
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2590 20448 2596 20460
rect 2551 20420 2596 20448
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 13372 20457 13400 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 16574 20476 16580 20528
rect 16632 20516 16638 20528
rect 18800 20525 18828 20556
rect 21453 20553 21465 20587
rect 21499 20584 21511 20587
rect 22370 20584 22376 20596
rect 21499 20556 22376 20584
rect 21499 20553 21511 20556
rect 21453 20547 21511 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 29365 20587 29423 20593
rect 29365 20553 29377 20587
rect 29411 20584 29423 20587
rect 30742 20584 30748 20596
rect 29411 20556 30748 20584
rect 29411 20553 29423 20556
rect 29365 20547 29423 20553
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 31018 20544 31024 20596
rect 31076 20584 31082 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 31076 20556 31309 20584
rect 31076 20544 31082 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 33965 20587 34023 20593
rect 33965 20553 33977 20587
rect 34011 20553 34023 20587
rect 33965 20547 34023 20553
rect 34609 20587 34667 20593
rect 34609 20553 34621 20587
rect 34655 20584 34667 20587
rect 35434 20584 35440 20596
rect 34655 20556 35440 20584
rect 34655 20553 34667 20556
rect 34609 20547 34667 20553
rect 32858 20525 32864 20528
rect 17098 20519 17156 20525
rect 17098 20516 17110 20519
rect 16632 20488 17110 20516
rect 16632 20476 16638 20488
rect 17098 20485 17110 20488
rect 17144 20485 17156 20519
rect 17098 20479 17156 20485
rect 18785 20519 18843 20525
rect 18785 20485 18797 20519
rect 18831 20485 18843 20519
rect 32852 20516 32864 20525
rect 18785 20479 18843 20485
rect 19076 20488 22094 20516
rect 32819 20488 32864 20516
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 13624 20451 13682 20457
rect 13624 20417 13636 20451
rect 13670 20448 13682 20451
rect 13906 20448 13912 20460
rect 13670 20420 13912 20448
rect 13670 20417 13682 20420
rect 13624 20411 13682 20417
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 15194 20448 15200 20460
rect 15155 20420 15200 20448
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 15654 20448 15660 20460
rect 15519 20420 15660 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20448 16911 20451
rect 16942 20448 16948 20460
rect 16899 20420 16948 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 19076 20457 19104 20488
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20329 20451 20387 20457
rect 20329 20448 20341 20451
rect 20036 20420 20341 20448
rect 20036 20408 20042 20420
rect 20329 20417 20341 20420
rect 20375 20417 20387 20451
rect 22066 20448 22094 20488
rect 32852 20479 32864 20488
rect 32858 20476 32864 20479
rect 32916 20476 32922 20528
rect 33980 20516 34008 20547
rect 35434 20544 35440 20556
rect 35492 20544 35498 20596
rect 36630 20584 36636 20596
rect 36591 20556 36636 20584
rect 36630 20544 36636 20556
rect 36688 20544 36694 20596
rect 37734 20584 37740 20596
rect 37695 20556 37740 20584
rect 37734 20544 37740 20556
rect 37792 20544 37798 20596
rect 35526 20516 35532 20528
rect 33980 20488 35532 20516
rect 35526 20476 35532 20488
rect 35584 20476 35590 20528
rect 35744 20519 35802 20525
rect 35744 20485 35756 20519
rect 35790 20516 35802 20519
rect 36722 20516 36728 20528
rect 35790 20488 36728 20516
rect 35790 20485 35802 20488
rect 35744 20479 35802 20485
rect 36722 20476 36728 20488
rect 36780 20476 36786 20528
rect 39114 20516 39120 20528
rect 39075 20488 39120 20516
rect 39114 20476 39120 20488
rect 39172 20476 39178 20528
rect 22554 20448 22560 20460
rect 22066 20420 22560 20448
rect 20329 20411 20387 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 27890 20408 27896 20460
rect 27948 20448 27954 20460
rect 28258 20457 28264 20460
rect 27985 20451 28043 20457
rect 27985 20448 27997 20451
rect 27948 20420 27997 20448
rect 27948 20408 27954 20420
rect 27985 20417 27997 20420
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28252 20411 28264 20457
rect 28316 20448 28322 20460
rect 29914 20448 29920 20460
rect 28316 20420 28352 20448
rect 29875 20420 29920 20448
rect 28258 20408 28264 20411
rect 28316 20408 28322 20420
rect 29914 20408 29920 20420
rect 29972 20408 29978 20460
rect 30006 20408 30012 20460
rect 30064 20448 30070 20460
rect 30173 20451 30231 20457
rect 30173 20448 30185 20451
rect 30064 20420 30185 20448
rect 30064 20408 30070 20420
rect 30173 20417 30185 20420
rect 30219 20417 30231 20451
rect 30173 20411 30231 20417
rect 35894 20408 35900 20460
rect 35952 20448 35958 20460
rect 35989 20451 36047 20457
rect 35989 20448 36001 20451
rect 35952 20420 36001 20448
rect 35952 20408 35958 20420
rect 35989 20417 36001 20420
rect 36035 20417 36047 20451
rect 36814 20448 36820 20460
rect 36775 20420 36820 20448
rect 35989 20411 36047 20417
rect 36814 20408 36820 20420
rect 36872 20408 36878 20460
rect 37918 20448 37924 20460
rect 37879 20420 37924 20448
rect 37918 20408 37924 20420
rect 37976 20408 37982 20460
rect 5810 20380 5816 20392
rect 5771 20352 5816 20380
rect 5810 20340 5816 20352
rect 5868 20340 5874 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15289 20383 15347 20389
rect 15289 20380 15301 20383
rect 14792 20352 15301 20380
rect 14792 20340 14798 20352
rect 15289 20349 15301 20352
rect 15335 20349 15347 20383
rect 18966 20380 18972 20392
rect 18927 20352 18972 20380
rect 15289 20343 15347 20349
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 20070 20380 20076 20392
rect 20031 20352 20076 20380
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 32306 20340 32312 20392
rect 32364 20380 32370 20392
rect 32585 20383 32643 20389
rect 32585 20380 32597 20383
rect 32364 20352 32597 20380
rect 32364 20340 32370 20352
rect 32585 20349 32597 20352
rect 32631 20349 32643 20383
rect 32585 20343 32643 20349
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20312 18291 20315
rect 18782 20312 18788 20324
rect 18279 20284 18788 20312
rect 18279 20281 18291 20284
rect 18233 20275 18291 20281
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 38838 20272 38844 20324
rect 38896 20312 38902 20324
rect 39393 20315 39451 20321
rect 39393 20312 39405 20315
rect 38896 20284 39405 20312
rect 38896 20272 38902 20284
rect 39393 20281 39405 20284
rect 39439 20281 39451 20315
rect 39393 20275 39451 20281
rect 12710 20244 12716 20256
rect 12671 20216 12716 20244
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 14737 20247 14795 20253
rect 14737 20213 14749 20247
rect 14783 20244 14795 20247
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 14783 20216 15209 20244
rect 14783 20213 14795 20216
rect 14737 20207 14795 20213
rect 15197 20213 15209 20216
rect 15243 20213 15255 20247
rect 19058 20244 19064 20256
rect 19019 20216 19064 20244
rect 15197 20207 15255 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19245 20247 19303 20253
rect 19245 20213 19257 20247
rect 19291 20244 19303 20247
rect 19334 20244 19340 20256
rect 19291 20216 19340 20244
rect 19291 20213 19303 20216
rect 19245 20207 19303 20213
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 39577 20247 39635 20253
rect 39577 20213 39589 20247
rect 39623 20244 39635 20247
rect 40126 20244 40132 20256
rect 39623 20216 40132 20244
rect 39623 20213 39635 20216
rect 39577 20207 39635 20213
rect 40126 20204 40132 20216
rect 40184 20204 40190 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 3418 20040 3424 20052
rect 3379 20012 3424 20040
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20040 13783 20043
rect 15194 20040 15200 20052
rect 13771 20012 15200 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15654 20040 15660 20052
rect 15615 20012 15660 20040
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 17957 20043 18015 20049
rect 17957 20009 17969 20043
rect 18003 20040 18015 20043
rect 18046 20040 18052 20052
rect 18003 20012 18052 20040
rect 18003 20009 18015 20012
rect 17957 20003 18015 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 21545 20043 21603 20049
rect 21545 20009 21557 20043
rect 21591 20040 21603 20043
rect 22094 20040 22100 20052
rect 21591 20012 22100 20040
rect 21591 20009 21603 20012
rect 21545 20003 21603 20009
rect 22094 20000 22100 20012
rect 22152 20000 22158 20052
rect 28258 20040 28264 20052
rect 28219 20012 28264 20040
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 30006 20040 30012 20052
rect 29967 20012 30012 20040
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 30466 20040 30472 20052
rect 30427 20012 30472 20040
rect 30466 20000 30472 20012
rect 30524 20000 30530 20052
rect 33502 20040 33508 20052
rect 33463 20012 33508 20040
rect 33502 20000 33508 20012
rect 33560 20000 33566 20052
rect 33689 20043 33747 20049
rect 33689 20009 33701 20043
rect 33735 20040 33747 20043
rect 34054 20040 34060 20052
rect 33735 20012 34060 20040
rect 33735 20009 33747 20012
rect 33689 20003 33747 20009
rect 34054 20000 34060 20012
rect 34112 20000 34118 20052
rect 35069 20043 35127 20049
rect 35069 20009 35081 20043
rect 35115 20040 35127 20043
rect 35342 20040 35348 20052
rect 35115 20012 35348 20040
rect 35115 20009 35127 20012
rect 35069 20003 35127 20009
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 13872 19876 14289 19904
rect 13872 19864 13878 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 33413 19907 33471 19913
rect 33413 19873 33425 19907
rect 33459 19904 33471 19907
rect 34514 19904 34520 19916
rect 33459 19876 34520 19904
rect 33459 19873 33471 19876
rect 33413 19867 33471 19873
rect 34514 19864 34520 19876
rect 34572 19864 34578 19916
rect 2038 19836 2044 19848
rect 1999 19808 2044 19836
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2314 19845 2320 19848
rect 2308 19836 2320 19845
rect 2275 19808 2320 19836
rect 2308 19799 2320 19808
rect 2314 19796 2320 19799
rect 2372 19796 2378 19848
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 13832 19836 13860 19864
rect 12391 19808 13860 19836
rect 16577 19839 16635 19845
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 16577 19805 16589 19839
rect 16623 19836 16635 19839
rect 16623 19808 16988 19836
rect 16623 19805 16635 19808
rect 16577 19799 16635 19805
rect 16960 19780 16988 19808
rect 20070 19796 20076 19848
rect 20128 19836 20134 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 20128 19808 20177 19836
rect 20128 19796 20134 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20432 19839 20490 19845
rect 20432 19805 20444 19839
rect 20478 19836 20490 19839
rect 22002 19836 22008 19848
rect 20478 19808 22008 19836
rect 20478 19805 20490 19808
rect 20432 19799 20490 19805
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 32122 19836 32128 19848
rect 32083 19808 32128 19836
rect 32122 19796 32128 19808
rect 32180 19796 32186 19848
rect 33226 19836 33232 19848
rect 33187 19808 33232 19836
rect 33226 19796 33232 19808
rect 33284 19796 33290 19848
rect 33505 19839 33563 19845
rect 33505 19805 33517 19839
rect 33551 19836 33563 19839
rect 33686 19836 33692 19848
rect 33551 19808 33692 19836
rect 33551 19805 33563 19808
rect 33505 19799 33563 19805
rect 33686 19796 33692 19808
rect 33744 19796 33750 19848
rect 12612 19771 12670 19777
rect 12612 19737 12624 19771
rect 12658 19768 12670 19771
rect 12710 19768 12716 19780
rect 12658 19740 12716 19768
rect 12658 19737 12670 19740
rect 12612 19731 12670 19737
rect 12710 19728 12716 19740
rect 12768 19728 12774 19780
rect 14550 19777 14556 19780
rect 14544 19731 14556 19777
rect 14608 19768 14614 19780
rect 14608 19740 14644 19768
rect 14550 19728 14556 19731
rect 14608 19728 14614 19740
rect 16666 19728 16672 19780
rect 16724 19768 16730 19780
rect 16822 19771 16880 19777
rect 16822 19768 16834 19771
rect 16724 19740 16834 19768
rect 16724 19728 16730 19740
rect 16822 19737 16834 19740
rect 16868 19737 16880 19771
rect 16822 19731 16880 19737
rect 16942 19728 16948 19780
rect 17000 19728 17006 19780
rect 18414 19700 18420 19712
rect 18375 19672 18420 19700
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 14734 19496 14740 19508
rect 14695 19468 14740 19496
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 33686 19496 33692 19508
rect 33647 19468 33692 19496
rect 33686 19456 33692 19468
rect 33744 19456 33750 19508
rect 13814 19428 13820 19440
rect 13372 19400 13820 19428
rect 5810 19320 5816 19372
rect 5868 19360 5874 19372
rect 6546 19360 6552 19372
rect 5868 19332 6552 19360
rect 5868 19320 5874 19332
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 13372 19369 13400 19400
rect 13814 19388 13820 19400
rect 13872 19388 13878 19440
rect 32122 19388 32128 19440
rect 32180 19428 32186 19440
rect 32554 19431 32612 19437
rect 32554 19428 32566 19431
rect 32180 19400 32566 19428
rect 32180 19388 32186 19400
rect 32554 19397 32566 19400
rect 32600 19397 32612 19431
rect 32554 19391 32612 19397
rect 13630 19369 13636 19372
rect 6805 19363 6863 19369
rect 6805 19360 6817 19363
rect 6656 19332 6817 19360
rect 5997 19295 6055 19301
rect 5997 19261 6009 19295
rect 6043 19292 6055 19295
rect 6656 19292 6684 19332
rect 6805 19329 6817 19332
rect 6851 19329 6863 19363
rect 6805 19323 6863 19329
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19329 13415 19363
rect 13624 19360 13636 19369
rect 13591 19332 13636 19360
rect 13357 19323 13415 19329
rect 13624 19323 13636 19332
rect 13630 19320 13636 19323
rect 13688 19320 13694 19372
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 17954 19360 17960 19372
rect 14884 19332 17960 19360
rect 14884 19320 14890 19332
rect 17954 19320 17960 19332
rect 18012 19360 18018 19372
rect 18414 19360 18420 19372
rect 18012 19332 18420 19360
rect 18012 19320 18018 19332
rect 18414 19320 18420 19332
rect 18472 19360 18478 19372
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 18472 19332 18521 19360
rect 18472 19320 18478 19332
rect 18509 19329 18521 19332
rect 18555 19329 18567 19363
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 18509 19323 18567 19329
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 6043 19264 6684 19292
rect 6043 19261 6055 19264
rect 5997 19255 6055 19261
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 2501 19159 2559 19165
rect 2501 19156 2513 19159
rect 2372 19128 2513 19156
rect 2372 19116 2378 19128
rect 2501 19125 2513 19128
rect 2547 19125 2559 19159
rect 7926 19156 7932 19168
rect 7887 19128 7932 19156
rect 2501 19119 2559 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 17402 19156 17408 19168
rect 17363 19128 17408 19156
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 19981 19159 20039 19165
rect 19981 19125 19993 19159
rect 20027 19156 20039 19159
rect 20070 19156 20076 19168
rect 20027 19128 20076 19156
rect 20027 19125 20039 19128
rect 19981 19119 20039 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 37826 19156 37832 19168
rect 37787 19128 37832 19156
rect 37826 19116 37832 19128
rect 37884 19116 37890 19168
rect 40954 19156 40960 19168
rect 40915 19128 40960 19156
rect 40954 19116 40960 19128
rect 41012 19116 41018 19168
rect 41785 19159 41843 19165
rect 41785 19125 41797 19159
rect 41831 19156 41843 19159
rect 42794 19156 42800 19168
rect 41831 19128 42800 19156
rect 41831 19125 41843 19128
rect 41785 19119 41843 19125
rect 42794 19116 42800 19128
rect 42852 19116 42858 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3973 18955 4031 18961
rect 3973 18952 3985 18955
rect 3467 18924 3985 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3973 18921 3985 18924
rect 4019 18921 4031 18955
rect 3973 18915 4031 18921
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18952 7435 18955
rect 7926 18952 7932 18964
rect 7423 18924 7932 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 14461 18955 14519 18961
rect 14461 18921 14473 18955
rect 14507 18952 14519 18955
rect 14550 18952 14556 18964
rect 14507 18924 14556 18952
rect 14507 18921 14519 18924
rect 14461 18915 14519 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 2038 18816 2044 18828
rect 1999 18788 2044 18816
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 3878 18776 3884 18828
rect 3936 18816 3942 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3936 18788 4077 18816
rect 3936 18776 3942 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 2314 18757 2320 18760
rect 2308 18748 2320 18757
rect 2275 18720 2320 18748
rect 2308 18711 2320 18720
rect 2314 18708 2320 18711
rect 2372 18708 2378 18760
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 4249 18751 4307 18757
rect 4249 18748 4261 18751
rect 4212 18720 4261 18748
rect 4212 18708 4218 18720
rect 4249 18717 4261 18720
rect 4295 18717 4307 18751
rect 5626 18748 5632 18760
rect 5587 18720 5632 18748
rect 4249 18711 4307 18717
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 7006 18708 7012 18760
rect 7064 18748 7070 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 7064 18720 7113 18748
rect 7064 18708 7070 18720
rect 7101 18717 7113 18720
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7926 18748 7932 18760
rect 7239 18720 7932 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 16850 18748 16856 18760
rect 16807 18720 16856 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 18598 18748 18604 18760
rect 18559 18720 18604 18748
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 21082 18748 21088 18760
rect 21043 18720 21088 18748
rect 20901 18711 20959 18717
rect 21082 18708 21088 18720
rect 21140 18708 21146 18760
rect 37093 18751 37151 18757
rect 37093 18717 37105 18751
rect 37139 18748 37151 18751
rect 37366 18748 37372 18760
rect 37139 18720 37372 18748
rect 37139 18717 37151 18720
rect 37093 18711 37151 18717
rect 37366 18708 37372 18720
rect 37424 18708 37430 18760
rect 37458 18708 37464 18760
rect 37516 18748 37522 18760
rect 37553 18751 37611 18757
rect 37553 18748 37565 18751
rect 37516 18720 37565 18748
rect 37516 18708 37522 18720
rect 37553 18717 37565 18720
rect 37599 18748 37611 18751
rect 40681 18751 40739 18757
rect 40681 18748 40693 18751
rect 37599 18720 40693 18748
rect 37599 18717 37611 18720
rect 37553 18711 37611 18717
rect 40681 18717 40693 18720
rect 40727 18748 40739 18751
rect 40770 18748 40776 18760
rect 40727 18720 40776 18748
rect 40727 18717 40739 18720
rect 40681 18711 40739 18717
rect 40770 18708 40776 18720
rect 40828 18708 40834 18760
rect 40954 18757 40960 18760
rect 40948 18748 40960 18757
rect 40915 18720 40960 18748
rect 40948 18711 40960 18720
rect 40954 18708 40960 18711
rect 41012 18708 41018 18760
rect 44450 18748 44456 18760
rect 44411 18720 44456 18748
rect 44450 18708 44456 18720
rect 44508 18708 44514 18760
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3973 18683 4031 18689
rect 3973 18680 3985 18683
rect 3568 18652 3985 18680
rect 3568 18640 3574 18652
rect 3973 18649 3985 18652
rect 4019 18649 4031 18683
rect 7374 18680 7380 18692
rect 7335 18652 7380 18680
rect 3973 18643 4031 18649
rect 7374 18640 7380 18652
rect 7432 18640 7438 18692
rect 16298 18640 16304 18692
rect 16356 18680 16362 18692
rect 37826 18689 37832 18692
rect 17006 18683 17064 18689
rect 17006 18680 17018 18683
rect 16356 18652 17018 18680
rect 16356 18640 16362 18652
rect 17006 18649 17018 18652
rect 17052 18649 17064 18683
rect 37820 18680 37832 18689
rect 37787 18652 37832 18680
rect 17006 18643 17064 18649
rect 37820 18643 37832 18652
rect 37826 18640 37832 18643
rect 37884 18640 37890 18692
rect 4430 18612 4436 18624
rect 4391 18584 4436 18612
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 6917 18615 6975 18621
rect 6917 18612 6929 18615
rect 4856 18584 6929 18612
rect 4856 18572 4862 18584
rect 6917 18581 6929 18584
rect 6963 18581 6975 18615
rect 6917 18575 6975 18581
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18782 18612 18788 18624
rect 18187 18584 18788 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 20990 18612 20996 18624
rect 20951 18584 20996 18612
rect 20990 18572 20996 18584
rect 21048 18572 21054 18624
rect 38930 18612 38936 18624
rect 38891 18584 38936 18612
rect 38930 18572 38936 18584
rect 38988 18572 38994 18624
rect 42061 18615 42119 18621
rect 42061 18581 42073 18615
rect 42107 18612 42119 18615
rect 42610 18612 42616 18624
rect 42107 18584 42616 18612
rect 42107 18581 42119 18584
rect 42061 18575 42119 18581
rect 42610 18572 42616 18584
rect 42668 18572 42674 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 3510 18408 3516 18420
rect 3471 18380 3516 18408
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 7926 18408 7932 18420
rect 7887 18380 7932 18408
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 19245 18411 19303 18417
rect 19245 18408 19257 18411
rect 19024 18380 19257 18408
rect 19024 18368 19030 18380
rect 19245 18377 19257 18380
rect 19291 18377 19303 18411
rect 19245 18371 19303 18377
rect 4706 18340 4712 18352
rect 4632 18312 4712 18340
rect 2038 18232 2044 18284
rect 2096 18272 2102 18284
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 2096 18244 2145 18272
rect 2096 18232 2102 18244
rect 2133 18241 2145 18244
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2222 18232 2228 18284
rect 2280 18272 2286 18284
rect 4632 18281 4660 18312
rect 4706 18300 4712 18312
rect 4764 18300 4770 18352
rect 7098 18340 7104 18352
rect 6564 18312 7104 18340
rect 6564 18284 6592 18312
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 18782 18340 18788 18352
rect 18743 18312 18788 18340
rect 18782 18300 18788 18312
rect 18840 18300 18846 18352
rect 44450 18349 44456 18352
rect 44444 18340 44456 18349
rect 44411 18312 44456 18340
rect 44444 18303 44456 18312
rect 44450 18300 44456 18303
rect 44508 18300 44514 18352
rect 2389 18275 2447 18281
rect 2389 18272 2401 18275
rect 2280 18244 2401 18272
rect 2280 18232 2286 18244
rect 2389 18241 2401 18244
rect 2435 18241 2447 18275
rect 2389 18235 2447 18241
rect 4617 18275 4675 18281
rect 4617 18241 4629 18275
rect 4663 18241 4675 18275
rect 4798 18272 4804 18284
rect 4759 18244 4804 18272
rect 4617 18235 4675 18241
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 6546 18272 6552 18284
rect 6507 18244 6552 18272
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 6805 18275 6863 18281
rect 6805 18272 6817 18275
rect 6656 18244 6817 18272
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18204 6055 18207
rect 6656 18204 6684 18244
rect 6805 18241 6817 18244
rect 6851 18241 6863 18275
rect 16298 18272 16304 18284
rect 16259 18244 16304 18272
rect 6805 18235 6863 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17201 18275 17259 18281
rect 17201 18272 17213 18275
rect 17092 18244 17213 18272
rect 17092 18232 17098 18244
rect 17201 18241 17213 18244
rect 17247 18241 17259 18275
rect 19058 18272 19064 18284
rect 19019 18244 19064 18272
rect 17201 18235 17259 18241
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 20340 18275 20398 18281
rect 20340 18241 20352 18275
rect 20386 18272 20398 18275
rect 20714 18272 20720 18284
rect 20386 18244 20720 18272
rect 20386 18241 20398 18244
rect 20340 18235 20398 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21450 18232 21456 18284
rect 21508 18272 21514 18284
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21508 18244 22017 18272
rect 21508 18232 21514 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22281 18275 22339 18281
rect 22152 18244 22197 18272
rect 22152 18232 22158 18244
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22922 18272 22928 18284
rect 22327 18244 22928 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 37728 18275 37786 18281
rect 37728 18241 37740 18275
rect 37774 18272 37786 18275
rect 39301 18275 39359 18281
rect 39301 18272 39313 18275
rect 37774 18244 39313 18272
rect 37774 18241 37786 18244
rect 37728 18235 37786 18241
rect 39301 18241 39313 18244
rect 39347 18241 39359 18275
rect 39301 18235 39359 18241
rect 40681 18275 40739 18281
rect 40681 18241 40693 18275
rect 40727 18272 40739 18275
rect 40770 18272 40776 18284
rect 40727 18244 40776 18272
rect 40727 18241 40739 18244
rect 40681 18235 40739 18241
rect 40770 18232 40776 18244
rect 40828 18232 40834 18284
rect 40954 18281 40960 18284
rect 40948 18235 40960 18281
rect 41012 18272 41018 18284
rect 41012 18244 41048 18272
rect 40954 18232 40960 18235
rect 41012 18232 41018 18244
rect 41966 18232 41972 18284
rect 42024 18272 42030 18284
rect 42613 18275 42671 18281
rect 42613 18272 42625 18275
rect 42024 18244 42625 18272
rect 42024 18232 42030 18244
rect 42613 18241 42625 18244
rect 42659 18241 42671 18275
rect 42613 18235 42671 18241
rect 42889 18275 42947 18281
rect 42889 18241 42901 18275
rect 42935 18272 42947 18275
rect 43990 18272 43996 18284
rect 42935 18244 43996 18272
rect 42935 18241 42947 18244
rect 42889 18235 42947 18241
rect 43990 18232 43996 18244
rect 44048 18232 44054 18284
rect 16942 18204 16948 18216
rect 6043 18176 6684 18204
rect 16903 18176 16948 18204
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 18874 18204 18880 18216
rect 18835 18176 18880 18204
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 20070 18204 20076 18216
rect 20031 18176 20076 18204
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 37458 18204 37464 18216
rect 37419 18176 37464 18204
rect 37458 18164 37464 18176
rect 37516 18164 37522 18216
rect 42705 18207 42763 18213
rect 42705 18173 42717 18207
rect 42751 18173 42763 18207
rect 42705 18167 42763 18173
rect 44177 18207 44235 18213
rect 44177 18173 44189 18207
rect 44223 18173 44235 18207
rect 44177 18167 44235 18173
rect 42061 18139 42119 18145
rect 42061 18105 42073 18139
rect 42107 18136 42119 18139
rect 42720 18136 42748 18167
rect 42107 18108 42748 18136
rect 42107 18105 42119 18108
rect 42061 18099 42119 18105
rect 3970 18068 3976 18080
rect 3931 18040 3976 18068
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4617 18071 4675 18077
rect 4617 18068 4629 18071
rect 4488 18040 4629 18068
rect 4488 18028 4494 18040
rect 4617 18037 4629 18040
rect 4663 18037 4675 18071
rect 4617 18031 4675 18037
rect 4985 18071 5043 18077
rect 4985 18037 4997 18071
rect 5031 18068 5043 18071
rect 5074 18068 5080 18080
rect 5031 18040 5080 18068
rect 5031 18037 5043 18040
rect 4985 18031 5043 18037
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 8386 18068 8392 18080
rect 8347 18040 8392 18068
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 18325 18071 18383 18077
rect 18325 18037 18337 18071
rect 18371 18068 18383 18071
rect 18785 18071 18843 18077
rect 18785 18068 18797 18071
rect 18371 18040 18797 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 18785 18037 18797 18040
rect 18831 18037 18843 18071
rect 21450 18068 21456 18080
rect 21411 18040 21456 18068
rect 18785 18031 18843 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22281 18071 22339 18077
rect 22281 18068 22293 18071
rect 22244 18040 22293 18068
rect 22244 18028 22250 18040
rect 22281 18037 22293 18040
rect 22327 18037 22339 18071
rect 36906 18068 36912 18080
rect 36867 18040 36912 18068
rect 22281 18031 22339 18037
rect 36906 18028 36912 18040
rect 36964 18028 36970 18080
rect 38838 18068 38844 18080
rect 38799 18040 38844 18068
rect 38838 18028 38844 18040
rect 38896 18028 38902 18080
rect 40221 18071 40279 18077
rect 40221 18037 40233 18071
rect 40267 18068 40279 18071
rect 40310 18068 40316 18080
rect 40267 18040 40316 18068
rect 40267 18037 40279 18040
rect 40221 18031 40279 18037
rect 40310 18028 40316 18040
rect 40368 18028 40374 18080
rect 42610 18068 42616 18080
rect 42571 18040 42616 18068
rect 42610 18028 42616 18040
rect 42668 18028 42674 18080
rect 43073 18071 43131 18077
rect 43073 18037 43085 18071
rect 43119 18068 43131 18071
rect 43346 18068 43352 18080
rect 43119 18040 43352 18068
rect 43119 18037 43131 18040
rect 43073 18031 43131 18037
rect 43346 18028 43352 18040
rect 43404 18028 43410 18080
rect 44192 18068 44220 18167
rect 44542 18068 44548 18080
rect 44192 18040 44548 18068
rect 44542 18028 44548 18040
rect 44600 18028 44606 18080
rect 45557 18071 45615 18077
rect 45557 18037 45569 18071
rect 45603 18068 45615 18071
rect 46290 18068 46296 18080
rect 45603 18040 46296 18068
rect 45603 18037 45615 18040
rect 45557 18031 45615 18037
rect 46290 18028 46296 18040
rect 46348 18028 46354 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 3421 17867 3479 17873
rect 3421 17833 3433 17867
rect 3467 17864 3479 17867
rect 3878 17864 3884 17876
rect 3467 17836 3884 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 7006 17864 7012 17876
rect 6595 17836 7012 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 17034 17864 17040 17876
rect 16995 17836 17040 17864
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 18877 17867 18935 17873
rect 18877 17833 18889 17867
rect 18923 17864 18935 17867
rect 19058 17864 19064 17876
rect 18923 17836 19064 17864
rect 18923 17833 18935 17836
rect 18877 17827 18935 17833
rect 19058 17824 19064 17836
rect 19116 17824 19122 17876
rect 38746 17864 38752 17876
rect 38707 17836 38752 17864
rect 38746 17824 38752 17836
rect 38804 17824 38810 17876
rect 43346 17864 43352 17876
rect 43307 17836 43352 17864
rect 43346 17824 43352 17836
rect 43404 17824 43410 17876
rect 22922 17796 22928 17808
rect 22883 17768 22928 17796
rect 22922 17756 22928 17768
rect 22980 17756 22986 17808
rect 2038 17728 2044 17740
rect 1999 17700 2044 17728
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 38838 17728 38844 17740
rect 17000 17700 17540 17728
rect 38799 17700 38844 17728
rect 17000 17688 17006 17700
rect 2308 17663 2366 17669
rect 2308 17629 2320 17663
rect 2354 17660 2366 17663
rect 3970 17660 3976 17672
rect 2354 17632 3976 17660
rect 2354 17629 2366 17632
rect 2308 17623 2366 17629
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4614 17660 4620 17672
rect 4203 17632 4620 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 6546 17660 6552 17672
rect 4672 17632 6552 17660
rect 4672 17620 4678 17632
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7116 17632 7941 17660
rect 7116 17604 7144 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 14642 17660 14648 17672
rect 14603 17632 14648 17660
rect 7929 17623 7987 17629
rect 14642 17620 14648 17632
rect 14700 17620 14706 17672
rect 17512 17669 17540 17700
rect 38838 17688 38844 17700
rect 38896 17688 38902 17740
rect 43438 17728 43444 17740
rect 43399 17700 43444 17728
rect 43438 17688 43444 17700
rect 43496 17688 43502 17740
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 17543 17632 19717 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 19705 17629 19717 17632
rect 19751 17660 19763 17663
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 19751 17632 21557 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 20088 17604 20116 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 36633 17663 36691 17669
rect 36633 17629 36645 17663
rect 36679 17660 36691 17663
rect 37458 17660 37464 17672
rect 36679 17632 37464 17660
rect 36679 17629 36691 17632
rect 36633 17623 36691 17629
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 38930 17660 38936 17672
rect 38891 17632 38936 17660
rect 38930 17620 38936 17632
rect 38988 17620 38994 17672
rect 43622 17660 43628 17672
rect 43583 17632 43628 17660
rect 43622 17620 43628 17632
rect 43680 17620 43686 17672
rect 44634 17660 44640 17672
rect 44595 17632 44640 17660
rect 44634 17620 44640 17632
rect 44692 17620 44698 17672
rect 45186 17660 45192 17672
rect 45147 17632 45192 17660
rect 45186 17620 45192 17632
rect 45244 17620 45250 17672
rect 7098 17592 7104 17604
rect 5460 17564 7104 17592
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5460 17533 5488 17564
rect 7098 17552 7104 17564
rect 7156 17552 7162 17604
rect 7684 17595 7742 17601
rect 7684 17561 7696 17595
rect 7730 17592 7742 17595
rect 8386 17592 8392 17604
rect 7730 17564 8392 17592
rect 7730 17561 7742 17564
rect 7684 17555 7742 17561
rect 8386 17552 8392 17564
rect 8444 17552 8450 17604
rect 17764 17595 17822 17601
rect 17764 17561 17776 17595
rect 17810 17592 17822 17595
rect 18598 17592 18604 17604
rect 17810 17564 18604 17592
rect 17810 17561 17822 17564
rect 17764 17555 17822 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 19972 17595 20030 17601
rect 19972 17561 19984 17595
rect 20018 17561 20030 17595
rect 19972 17555 20030 17561
rect 5445 17527 5503 17533
rect 5445 17524 5457 17527
rect 4672 17496 5457 17524
rect 4672 17484 4678 17496
rect 5445 17493 5457 17496
rect 5491 17493 5503 17527
rect 19996 17524 20024 17555
rect 20070 17552 20076 17604
rect 20128 17552 20134 17604
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 36906 17601 36912 17604
rect 21790 17595 21848 17601
rect 21790 17592 21802 17595
rect 21692 17564 21802 17592
rect 21692 17552 21698 17564
rect 21790 17561 21802 17564
rect 21836 17561 21848 17595
rect 36900 17592 36912 17601
rect 36867 17564 36912 17592
rect 21790 17555 21848 17561
rect 36900 17555 36912 17564
rect 36906 17552 36912 17555
rect 36964 17552 36970 17604
rect 38657 17595 38715 17601
rect 38657 17561 38669 17595
rect 38703 17561 38715 17595
rect 38657 17555 38715 17561
rect 40681 17595 40739 17601
rect 40681 17561 40693 17595
rect 40727 17592 40739 17595
rect 41138 17592 41144 17604
rect 40727 17564 41144 17592
rect 40727 17561 40739 17564
rect 40681 17555 40739 17561
rect 20990 17524 20996 17536
rect 19996 17496 20996 17524
rect 5445 17487 5503 17493
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21085 17527 21143 17533
rect 21085 17493 21097 17527
rect 21131 17524 21143 17527
rect 22094 17524 22100 17536
rect 21131 17496 22100 17524
rect 21131 17493 21143 17496
rect 21085 17487 21143 17493
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 38013 17527 38071 17533
rect 38013 17493 38025 17527
rect 38059 17524 38071 17527
rect 38672 17524 38700 17555
rect 41138 17552 41144 17564
rect 41196 17552 41202 17604
rect 42886 17592 42892 17604
rect 42847 17564 42892 17592
rect 42886 17552 42892 17564
rect 42944 17552 42950 17604
rect 43349 17595 43407 17601
rect 43349 17561 43361 17595
rect 43395 17561 43407 17595
rect 43349 17555 43407 17561
rect 38059 17496 38700 17524
rect 39117 17527 39175 17533
rect 38059 17493 38071 17496
rect 38013 17487 38071 17493
rect 39117 17493 39129 17527
rect 39163 17524 39175 17527
rect 43364 17524 43392 17555
rect 39163 17496 43392 17524
rect 43809 17527 43867 17533
rect 39163 17493 39175 17496
rect 39117 17487 39175 17493
rect 43809 17493 43821 17527
rect 43855 17524 43867 17527
rect 43898 17524 43904 17536
rect 43855 17496 43904 17524
rect 43855 17493 43867 17496
rect 43809 17487 43867 17493
rect 43898 17484 43904 17496
rect 43956 17484 43962 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4154 17320 4160 17332
rect 4019 17292 4160 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 18417 17323 18475 17329
rect 18417 17289 18429 17323
rect 18463 17320 18475 17323
rect 18874 17320 18880 17332
rect 18463 17292 18880 17320
rect 18463 17289 18475 17292
rect 18417 17283 18475 17289
rect 18874 17280 18880 17292
rect 18932 17280 18938 17332
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 21082 17320 21088 17332
rect 20855 17292 21088 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 22215 17323 22273 17329
rect 22215 17289 22227 17323
rect 22261 17320 22273 17323
rect 22922 17320 22928 17332
rect 22261 17292 22928 17320
rect 22261 17289 22273 17292
rect 22215 17283 22273 17289
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 38746 17280 38752 17332
rect 38804 17320 38810 17332
rect 38841 17323 38899 17329
rect 38841 17320 38853 17323
rect 38804 17292 38853 17320
rect 38804 17280 38810 17292
rect 38841 17289 38853 17292
rect 38887 17289 38899 17323
rect 38841 17283 38899 17289
rect 41601 17323 41659 17329
rect 41601 17289 41613 17323
rect 41647 17320 41659 17323
rect 41966 17320 41972 17332
rect 41647 17292 41972 17320
rect 41647 17289 41659 17292
rect 41601 17283 41659 17289
rect 41966 17280 41972 17292
rect 42024 17280 42030 17332
rect 42794 17280 42800 17332
rect 42852 17320 42858 17332
rect 42852 17292 42932 17320
rect 42852 17280 42858 17292
rect 4884 17255 4942 17261
rect 2608 17224 4660 17252
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 2608 17193 2636 17224
rect 4632 17196 4660 17224
rect 4884 17221 4896 17255
rect 4930 17252 4942 17255
rect 5626 17252 5632 17264
rect 4930 17224 5632 17252
rect 4930 17221 4942 17224
rect 4884 17215 4942 17221
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 14642 17261 14648 17264
rect 14636 17252 14648 17261
rect 14603 17224 14648 17252
rect 14636 17215 14648 17224
rect 14642 17212 14648 17215
rect 14700 17212 14706 17264
rect 17304 17255 17362 17261
rect 17304 17221 17316 17255
rect 17350 17252 17362 17255
rect 17402 17252 17408 17264
rect 17350 17224 17408 17252
rect 17350 17221 17362 17224
rect 17304 17215 17362 17221
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 22005 17255 22063 17261
rect 22005 17221 22017 17255
rect 22051 17252 22063 17255
rect 22094 17252 22100 17264
rect 22051 17224 22100 17252
rect 22051 17221 22063 17224
rect 22005 17215 22063 17221
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 2096 17156 2605 17184
rect 2096 17144 2102 17156
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 2860 17187 2918 17193
rect 2860 17153 2872 17187
rect 2906 17184 2918 17187
rect 3970 17184 3976 17196
rect 2906 17156 3976 17184
rect 2906 17153 2918 17156
rect 2860 17147 2918 17153
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 4614 17184 4620 17196
rect 4527 17156 4620 17184
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 17000 17156 17049 17184
rect 17000 17144 17006 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 22020 17184 22048 17215
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 37366 17212 37372 17264
rect 37424 17252 37430 17264
rect 42904 17261 42932 17292
rect 43622 17280 43628 17332
rect 43680 17320 43686 17332
rect 46753 17323 46811 17329
rect 46753 17320 46765 17323
rect 43680 17292 46765 17320
rect 43680 17280 43686 17292
rect 46753 17289 46765 17292
rect 46799 17289 46811 17323
rect 46753 17283 46811 17289
rect 37706 17255 37764 17261
rect 37706 17252 37718 17255
rect 37424 17224 37718 17252
rect 37424 17212 37430 17224
rect 37706 17221 37718 17224
rect 37752 17221 37764 17255
rect 42880 17255 42938 17261
rect 37706 17215 37764 17221
rect 40236 17224 40816 17252
rect 37458 17184 37464 17196
rect 21223 17156 22048 17184
rect 37419 17156 37464 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 37458 17144 37464 17156
rect 37516 17144 37522 17196
rect 40034 17144 40040 17196
rect 40092 17184 40098 17196
rect 40236 17193 40264 17224
rect 40788 17196 40816 17224
rect 42880 17221 42892 17255
rect 42926 17221 42938 17255
rect 42880 17215 42938 17221
rect 44720 17255 44778 17261
rect 44720 17221 44732 17255
rect 44766 17252 44778 17255
rect 45186 17252 45192 17264
rect 44766 17224 45192 17252
rect 44766 17221 44778 17224
rect 44720 17215 44778 17221
rect 45186 17212 45192 17224
rect 45244 17212 45250 17264
rect 40221 17187 40279 17193
rect 40221 17184 40233 17187
rect 40092 17156 40233 17184
rect 40092 17144 40098 17156
rect 40221 17153 40233 17156
rect 40267 17153 40279 17187
rect 40221 17147 40279 17153
rect 40310 17144 40316 17196
rect 40368 17184 40374 17196
rect 40477 17187 40535 17193
rect 40477 17184 40489 17187
rect 40368 17156 40489 17184
rect 40368 17144 40374 17156
rect 40477 17153 40489 17156
rect 40523 17153 40535 17187
rect 40477 17147 40535 17153
rect 40770 17144 40776 17196
rect 40828 17184 40834 17196
rect 44453 17187 44511 17193
rect 40828 17156 42656 17184
rect 40828 17144 40834 17156
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17116 2191 17119
rect 2222 17116 2228 17128
rect 2179 17088 2228 17116
rect 2179 17085 2191 17088
rect 2133 17079 2191 17085
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 14332 17088 14381 17116
rect 14332 17076 14338 17088
rect 14369 17085 14381 17088
rect 14415 17085 14427 17119
rect 21082 17116 21088 17128
rect 21043 17088 21088 17116
rect 14369 17079 14427 17085
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 42628 17125 42656 17156
rect 44453 17153 44465 17187
rect 44499 17184 44511 17187
rect 44542 17184 44548 17196
rect 44499 17156 44548 17184
rect 44499 17153 44511 17156
rect 44453 17147 44511 17153
rect 44542 17144 44548 17156
rect 44600 17144 44606 17196
rect 45554 17144 45560 17196
rect 45612 17184 45618 17196
rect 46293 17187 46351 17193
rect 46293 17184 46305 17187
rect 45612 17156 46305 17184
rect 45612 17144 45618 17156
rect 46293 17153 46305 17156
rect 46339 17153 46351 17187
rect 46566 17184 46572 17196
rect 46527 17156 46572 17184
rect 46293 17147 46351 17153
rect 46566 17144 46572 17156
rect 46624 17144 46630 17196
rect 42613 17119 42671 17125
rect 42613 17085 42625 17119
rect 42659 17085 42671 17119
rect 42613 17079 42671 17085
rect 46385 17119 46443 17125
rect 46385 17085 46397 17119
rect 46431 17085 46443 17119
rect 46385 17079 46443 17085
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 7374 17048 7380 17060
rect 6043 17020 7380 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 6546 16980 6552 16992
rect 6507 16952 6552 16980
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 15749 16983 15807 16989
rect 15749 16949 15761 16983
rect 15795 16980 15807 16983
rect 16114 16980 16120 16992
rect 15795 16952 16120 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 21082 16940 21088 16992
rect 21140 16980 21146 16992
rect 21450 16980 21456 16992
rect 21140 16952 21456 16980
rect 21140 16940 21146 16952
rect 21450 16940 21456 16952
rect 21508 16980 21514 16992
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 21508 16952 22201 16980
rect 21508 16940 21514 16952
rect 22189 16949 22201 16952
rect 22235 16949 22247 16983
rect 22370 16980 22376 16992
rect 22331 16952 22376 16980
rect 22189 16943 22247 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 42628 16980 42656 17079
rect 43990 17048 43996 17060
rect 43951 17020 43996 17048
rect 43990 17008 43996 17020
rect 44048 17008 44054 17060
rect 45833 17051 45891 17057
rect 45833 17017 45845 17051
rect 45879 17048 45891 17051
rect 46400 17048 46428 17079
rect 45879 17020 46428 17048
rect 45879 17017 45891 17020
rect 45833 17011 45891 17017
rect 42794 16980 42800 16992
rect 42628 16952 42800 16980
rect 42794 16940 42800 16952
rect 42852 16940 42858 16992
rect 46290 16980 46296 16992
rect 46251 16952 46296 16980
rect 46290 16940 46296 16952
rect 46348 16940 46354 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 3970 16776 3976 16788
rect 3931 16748 3976 16776
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 16114 16776 16120 16788
rect 16075 16748 16120 16776
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 21545 16779 21603 16785
rect 21545 16745 21557 16779
rect 21591 16776 21603 16779
rect 21634 16776 21640 16788
rect 21591 16748 21640 16776
rect 21591 16745 21603 16748
rect 21545 16739 21603 16745
rect 21634 16736 21640 16748
rect 21692 16736 21698 16788
rect 40954 16776 40960 16788
rect 40915 16748 40960 16776
rect 40954 16736 40960 16748
rect 41012 16736 41018 16788
rect 46566 16776 46572 16788
rect 46527 16748 46572 16776
rect 46566 16736 46572 16748
rect 46624 16736 46630 16788
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21453 16711 21511 16717
rect 21453 16708 21465 16711
rect 20864 16680 21465 16708
rect 20864 16668 20870 16680
rect 21453 16677 21465 16680
rect 21499 16677 21511 16711
rect 21453 16671 21511 16677
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14182 16640 14188 16652
rect 13771 16612 14188 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 16206 16640 16212 16652
rect 16167 16612 16212 16640
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 21082 16640 21088 16652
rect 20916 16612 21088 16640
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16572 16451 16575
rect 16482 16572 16488 16584
rect 16439 16544 16488 16572
rect 16439 16541 16451 16544
rect 16393 16535 16451 16541
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16572 20775 16575
rect 20806 16572 20812 16584
rect 20763 16544 20812 16572
rect 20763 16541 20775 16544
rect 20717 16535 20775 16541
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 20916 16581 20944 16612
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 42794 16600 42800 16652
rect 42852 16640 42858 16652
rect 43165 16643 43223 16649
rect 43165 16640 43177 16643
rect 42852 16612 43177 16640
rect 42852 16600 42858 16612
rect 43165 16609 43177 16612
rect 43211 16640 43223 16643
rect 44542 16640 44548 16652
rect 43211 16612 44548 16640
rect 43211 16609 43223 16612
rect 43165 16603 43223 16609
rect 44542 16600 44548 16612
rect 44600 16640 44606 16652
rect 45189 16643 45247 16649
rect 45189 16640 45201 16643
rect 44600 16612 45201 16640
rect 44600 16600 44606 16612
rect 45189 16609 45201 16612
rect 45235 16609 45247 16643
rect 45189 16603 45247 16609
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 22186 16572 22192 16584
rect 21361 16535 21419 16541
rect 21560 16544 22192 16572
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 14522 16507 14580 16513
rect 14522 16504 14534 16507
rect 14148 16476 14534 16504
rect 14148 16464 14154 16476
rect 14522 16473 14534 16476
rect 14568 16473 14580 16507
rect 14522 16467 14580 16473
rect 16117 16507 16175 16513
rect 16117 16473 16129 16507
rect 16163 16473 16175 16507
rect 21376 16504 21404 16535
rect 21560 16504 21588 16544
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 41138 16532 41144 16584
rect 41196 16572 41202 16584
rect 41417 16575 41475 16581
rect 41417 16572 41429 16575
rect 41196 16544 41429 16572
rect 41196 16532 41202 16544
rect 41417 16541 41429 16544
rect 41463 16541 41475 16575
rect 44450 16572 44456 16584
rect 44411 16544 44456 16572
rect 41417 16535 41475 16541
rect 44450 16532 44456 16544
rect 44508 16532 44514 16584
rect 44634 16532 44640 16584
rect 44692 16572 44698 16584
rect 45445 16575 45503 16581
rect 45445 16572 45457 16575
rect 44692 16544 45457 16572
rect 44692 16532 44698 16544
rect 45445 16541 45457 16544
rect 45491 16541 45503 16575
rect 45445 16535 45503 16541
rect 21376 16476 21588 16504
rect 21637 16507 21695 16513
rect 16117 16467 16175 16473
rect 21637 16473 21649 16507
rect 21683 16504 21695 16507
rect 22370 16504 22376 16516
rect 21683 16476 22376 16504
rect 21683 16473 21695 16476
rect 21637 16467 21695 16473
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16436 15715 16439
rect 16132 16436 16160 16467
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 15703 16408 16160 16436
rect 16577 16439 16635 16445
rect 15703 16405 15715 16408
rect 15657 16399 15715 16405
rect 16577 16405 16589 16439
rect 16623 16436 16635 16439
rect 17770 16436 17776 16448
rect 16623 16408 17776 16436
rect 16623 16405 16635 16408
rect 16577 16399 16635 16405
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 15933 16235 15991 16241
rect 15933 16201 15945 16235
rect 15979 16232 15991 16235
rect 16206 16232 16212 16244
rect 15979 16204 16212 16232
rect 15979 16201 15991 16204
rect 15933 16195 15991 16201
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 20806 16232 20812 16244
rect 19444 16204 20812 16232
rect 14182 16124 14188 16176
rect 14240 16164 14246 16176
rect 19444 16173 19472 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 41138 16192 41144 16244
rect 41196 16232 41202 16244
rect 41233 16235 41291 16241
rect 41233 16232 41245 16235
rect 41196 16204 41245 16232
rect 41196 16192 41202 16204
rect 41233 16201 41245 16204
rect 41279 16201 41291 16235
rect 41233 16195 41291 16201
rect 45465 16235 45523 16241
rect 45465 16201 45477 16235
rect 45511 16232 45523 16235
rect 45554 16232 45560 16244
rect 45511 16204 45560 16232
rect 45511 16201 45523 16204
rect 45465 16195 45523 16201
rect 45554 16192 45560 16204
rect 45612 16192 45618 16244
rect 14798 16167 14856 16173
rect 14798 16164 14810 16167
rect 14240 16136 14810 16164
rect 14240 16124 14246 16136
rect 14798 16133 14810 16136
rect 14844 16133 14856 16167
rect 14798 16127 14856 16133
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 19613 16167 19671 16173
rect 19613 16133 19625 16167
rect 19659 16164 19671 16167
rect 20254 16164 20260 16176
rect 19659 16136 20260 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20254 16124 20260 16136
rect 20312 16124 20318 16176
rect 44352 16167 44410 16173
rect 44352 16133 44364 16167
rect 44398 16164 44410 16167
rect 44450 16164 44456 16176
rect 44398 16136 44456 16164
rect 44398 16133 44410 16136
rect 44352 16127 44410 16133
rect 44450 16124 44456 16136
rect 44508 16124 44514 16176
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16096 8815 16099
rect 9122 16096 9128 16108
rect 8803 16068 9128 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 14090 16096 14096 16108
rect 14051 16068 14096 16096
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 20070 16096 20076 16108
rect 19751 16068 20076 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16096 20407 16099
rect 20898 16096 20904 16108
rect 20395 16068 20904 16096
rect 20395 16065 20407 16068
rect 20349 16059 20407 16065
rect 14274 15988 14280 16040
rect 14332 16028 14338 16040
rect 14550 16028 14556 16040
rect 14332 16000 14556 16028
rect 14332 15988 14338 16000
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 19978 15988 19984 16040
rect 20036 16028 20042 16040
rect 20180 16028 20208 16059
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 42794 16056 42800 16108
rect 42852 16096 42858 16108
rect 43806 16096 43812 16108
rect 42852 16068 43812 16096
rect 42852 16056 42858 16068
rect 43806 16056 43812 16068
rect 43864 16096 43870 16108
rect 44085 16099 44143 16105
rect 44085 16096 44097 16099
rect 43864 16068 44097 16096
rect 43864 16056 43870 16068
rect 44085 16065 44097 16068
rect 44131 16065 44143 16099
rect 44085 16059 44143 16065
rect 20036 16000 20208 16028
rect 20036 15988 20042 16000
rect 8938 15892 8944 15904
rect 8899 15864 8944 15892
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 16850 15892 16856 15904
rect 16811 15864 16856 15892
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 20257 15895 20315 15901
rect 20257 15892 20269 15895
rect 20128 15864 20269 15892
rect 20128 15852 20134 15864
rect 20257 15861 20269 15864
rect 20303 15861 20315 15895
rect 20257 15855 20315 15861
rect 40129 15895 40187 15901
rect 40129 15861 40141 15895
rect 40175 15892 40187 15895
rect 40310 15892 40316 15904
rect 40175 15864 40316 15892
rect 40175 15861 40187 15864
rect 40129 15855 40187 15861
rect 40310 15852 40316 15864
rect 40368 15852 40374 15904
rect 40586 15892 40592 15904
rect 40547 15864 40592 15892
rect 40586 15852 40592 15864
rect 40644 15852 40650 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 8202 15688 8208 15700
rect 7883 15660 8208 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 20073 15691 20131 15697
rect 20073 15657 20085 15691
rect 20119 15688 20131 15691
rect 20806 15688 20812 15700
rect 20119 15660 20812 15688
rect 20119 15657 20131 15660
rect 20073 15651 20131 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 41417 15691 41475 15697
rect 41417 15657 41429 15691
rect 41463 15688 41475 15691
rect 41877 15691 41935 15697
rect 41877 15688 41889 15691
rect 41463 15660 41889 15688
rect 41463 15657 41475 15660
rect 41417 15651 41475 15657
rect 41877 15657 41889 15660
rect 41923 15657 41935 15691
rect 41877 15651 41935 15657
rect 42337 15691 42395 15697
rect 42337 15657 42349 15691
rect 42383 15688 42395 15691
rect 43438 15688 43444 15700
rect 42383 15660 43444 15688
rect 42383 15657 42395 15660
rect 42337 15651 42395 15657
rect 43438 15648 43444 15660
rect 43496 15648 43502 15700
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 22278 15552 22284 15564
rect 19392 15524 19564 15552
rect 19392 15512 19398 15524
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 10238 15487 10296 15493
rect 10238 15484 10250 15487
rect 8996 15456 10250 15484
rect 8996 15444 9002 15456
rect 10238 15453 10250 15456
rect 10284 15453 10296 15487
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10238 15447 10296 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15372 15487 15430 15493
rect 15372 15453 15384 15487
rect 15418 15484 15430 15487
rect 16850 15484 16856 15496
rect 15418 15456 16856 15484
rect 15418 15453 15430 15456
rect 15372 15447 15430 15453
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 19536 15493 19564 15524
rect 22020 15524 22284 15552
rect 22020 15493 22048 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 40034 15552 40040 15564
rect 39995 15524 40040 15552
rect 40034 15512 40040 15524
rect 40092 15512 40098 15564
rect 41966 15552 41972 15564
rect 41927 15524 41972 15552
rect 41966 15512 41972 15524
rect 42024 15512 42030 15564
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19300 15456 19441 15484
rect 19300 15444 19306 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 22005 15487 22063 15493
rect 19935 15456 20944 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20916 15428 20944 15456
rect 22005 15453 22017 15487
rect 22051 15453 22063 15487
rect 22186 15484 22192 15496
rect 22147 15456 22192 15484
rect 22005 15447 22063 15453
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15453 22891 15487
rect 22833 15447 22891 15453
rect 39485 15487 39543 15493
rect 39485 15453 39497 15487
rect 39531 15484 39543 15487
rect 39574 15484 39580 15496
rect 39531 15456 39580 15484
rect 39531 15453 39543 15456
rect 39485 15447 39543 15453
rect 8018 15416 8024 15428
rect 7979 15388 8024 15416
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19392 15388 19717 15416
rect 19392 15376 19398 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 19705 15379 19763 15385
rect 19797 15419 19855 15425
rect 19797 15385 19809 15419
rect 19843 15416 19855 15419
rect 19978 15416 19984 15428
rect 19843 15388 19984 15416
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 19978 15376 19984 15388
rect 20036 15416 20042 15428
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 20036 15388 20729 15416
rect 20036 15376 20042 15388
rect 20717 15385 20729 15388
rect 20763 15385 20775 15419
rect 20717 15379 20775 15385
rect 20898 15376 20904 15428
rect 20956 15416 20962 15428
rect 21821 15419 21879 15425
rect 21821 15416 21833 15419
rect 20956 15388 21833 15416
rect 20956 15376 20962 15388
rect 21821 15385 21833 15388
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 22848 15416 22876 15447
rect 39574 15444 39580 15456
rect 39632 15444 39638 15496
rect 40304 15487 40362 15493
rect 40304 15453 40316 15487
rect 40350 15484 40362 15487
rect 40586 15484 40592 15496
rect 40350 15456 40592 15484
rect 40350 15453 40362 15456
rect 40304 15447 40362 15453
rect 40586 15444 40592 15456
rect 40644 15444 40650 15496
rect 42150 15484 42156 15496
rect 42111 15456 42156 15484
rect 42150 15444 42156 15456
rect 42208 15444 42214 15496
rect 43714 15484 43720 15496
rect 43675 15456 43720 15484
rect 43714 15444 43720 15456
rect 43772 15444 43778 15496
rect 41874 15416 41880 15428
rect 22152 15388 22876 15416
rect 41835 15388 41880 15416
rect 22152 15376 22158 15388
rect 41874 15376 41880 15388
rect 41932 15376 41938 15428
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 7821 15351 7879 15357
rect 7821 15317 7833 15351
rect 7867 15348 7879 15351
rect 8938 15348 8944 15360
rect 7867 15320 8944 15348
rect 7867 15317 7879 15320
rect 7821 15311 7879 15317
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 20530 15348 20536 15360
rect 20491 15320 20536 15348
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 22646 15348 22652 15360
rect 22607 15320 22652 15348
rect 22646 15308 22652 15320
rect 22704 15308 22710 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 8938 15144 8944 15156
rect 8899 15116 8944 15144
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 19334 15144 19340 15156
rect 18739 15116 19340 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 4614 15076 4620 15088
rect 3528 15048 4620 15076
rect 3528 15017 3556 15048
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 9306 15076 9312 15088
rect 9219 15048 9312 15076
rect 9306 15036 9312 15048
rect 9364 15076 9370 15088
rect 10045 15079 10103 15085
rect 10045 15076 10057 15079
rect 9364 15048 10057 15076
rect 9364 15036 9370 15048
rect 10045 15045 10057 15048
rect 10091 15045 10103 15079
rect 10045 15039 10103 15045
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 11204 15048 11713 15076
rect 11204 15036 11210 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 11790 15036 11796 15088
rect 11848 15076 11854 15088
rect 11901 15079 11959 15085
rect 11901 15076 11913 15079
rect 11848 15048 11913 15076
rect 11848 15036 11854 15048
rect 11901 15045 11913 15048
rect 11947 15045 11959 15079
rect 11901 15039 11959 15045
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 3769 15011 3827 15017
rect 3769 15008 3781 15011
rect 3660 14980 3781 15008
rect 3660 14968 3666 14980
rect 3769 14977 3781 14980
rect 3815 14977 3827 15011
rect 7098 15008 7104 15020
rect 7059 14980 7104 15008
rect 3769 14971 3827 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7374 15017 7380 15020
rect 7368 14971 7380 15017
rect 7432 15008 7438 15020
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 7432 14980 7468 15008
rect 8496 14980 9137 15008
rect 7374 14968 7380 14971
rect 7432 14968 7438 14980
rect 8496 14881 8524 14980
rect 9125 14977 9137 14980
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 9447 14980 10241 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 10229 14977 10241 14980
rect 10275 15008 10287 15011
rect 10962 15008 10968 15020
rect 10275 14980 10968 15008
rect 10275 14977 10287 14980
rect 10229 14971 10287 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 14826 15008 14832 15020
rect 12575 14980 14832 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18708 15008 18736 15107
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 21453 15147 21511 15153
rect 21453 15113 21465 15147
rect 21499 15144 21511 15147
rect 22094 15144 22100 15156
rect 21499 15116 22100 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 23385 15147 23443 15153
rect 23385 15144 23397 15147
rect 22244 15116 23397 15144
rect 22244 15104 22250 15116
rect 23385 15113 23397 15116
rect 23431 15113 23443 15147
rect 23385 15107 23443 15113
rect 40681 15147 40739 15153
rect 40681 15113 40693 15147
rect 40727 15144 40739 15147
rect 41874 15144 41880 15156
rect 40727 15116 41880 15144
rect 40727 15113 40739 15116
rect 40681 15107 40739 15113
rect 41874 15104 41880 15116
rect 41932 15104 41938 15156
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 19806 15079 19864 15085
rect 19806 15076 19818 15079
rect 19484 15048 19818 15076
rect 19484 15036 19490 15048
rect 19806 15045 19818 15048
rect 19852 15045 19864 15079
rect 19806 15039 19864 15045
rect 20438 15036 20444 15088
rect 20496 15076 20502 15088
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 20496 15048 21281 15076
rect 20496 15036 20502 15048
rect 21269 15045 21281 15048
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 22272 15079 22330 15085
rect 22272 15045 22284 15079
rect 22318 15076 22330 15079
rect 22646 15076 22652 15088
rect 22318 15048 22652 15076
rect 22318 15045 22330 15048
rect 22272 15039 22330 15045
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 20898 15008 20904 15020
rect 18279 14980 18736 15008
rect 20859 14980 20904 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 39574 15017 39580 15020
rect 39568 15008 39580 15017
rect 39535 14980 39580 15008
rect 39568 14971 39580 14980
rect 39574 14968 39580 14971
rect 39632 14968 39638 15020
rect 43806 15008 43812 15020
rect 43767 14980 43812 15008
rect 43806 14968 43812 14980
rect 43864 14968 43870 15020
rect 44076 15011 44134 15017
rect 44076 14977 44088 15011
rect 44122 15008 44134 15011
rect 45830 15008 45836 15020
rect 44122 14980 45836 15008
rect 44122 14977 44134 14980
rect 44076 14971 44134 14977
rect 45830 14968 45836 14980
rect 45888 14968 45894 15020
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20622 14940 20628 14952
rect 20119 14912 20628 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20622 14900 20628 14912
rect 20680 14940 20686 14952
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 20680 14912 22017 14940
rect 20680 14900 20686 14912
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 39114 14900 39120 14952
rect 39172 14940 39178 14952
rect 39301 14943 39359 14949
rect 39301 14940 39313 14943
rect 39172 14912 39313 14940
rect 39172 14900 39178 14912
rect 39301 14909 39313 14912
rect 39347 14909 39359 14943
rect 39301 14903 39359 14909
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14872 8539 14875
rect 8570 14872 8576 14884
rect 8527 14844 8576 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 12069 14875 12127 14881
rect 12069 14841 12081 14875
rect 12115 14872 12127 14875
rect 13722 14872 13728 14884
rect 12115 14844 13728 14872
rect 12115 14841 12127 14844
rect 12069 14835 12127 14841
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 4893 14807 4951 14813
rect 4893 14773 4905 14807
rect 4939 14804 4951 14807
rect 5626 14804 5632 14816
rect 4939 14776 5632 14804
rect 4939 14773 4951 14776
rect 4893 14767 4951 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9364 14776 9873 14804
rect 9364 14764 9370 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9861 14767 9919 14773
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11756 14776 11897 14804
rect 11756 14764 11762 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 11885 14767 11943 14773
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 13136 14776 13829 14804
rect 13136 14764 13142 14776
rect 13817 14773 13829 14776
rect 13863 14804 13875 14807
rect 14550 14804 14556 14816
rect 13863 14776 14556 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14826 14804 14832 14816
rect 14787 14776 14832 14804
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 18141 14807 18199 14813
rect 18141 14773 18153 14807
rect 18187 14804 18199 14807
rect 20254 14804 20260 14816
rect 18187 14776 20260 14804
rect 18187 14773 18199 14776
rect 18141 14767 18199 14773
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14804 21327 14807
rect 21910 14804 21916 14816
rect 21315 14776 21916 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 21910 14764 21916 14776
rect 21968 14764 21974 14816
rect 41138 14804 41144 14816
rect 41099 14776 41144 14804
rect 41138 14764 41144 14776
rect 41196 14764 41202 14816
rect 45189 14807 45247 14813
rect 45189 14773 45201 14807
rect 45235 14804 45247 14807
rect 45554 14804 45560 14816
rect 45235 14776 45560 14804
rect 45235 14773 45247 14776
rect 45189 14767 45247 14773
rect 45554 14764 45560 14776
rect 45612 14764 45618 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3602 14600 3608 14612
rect 3467 14572 3608 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7432 14572 7573 14600
rect 7432 14560 7438 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 8904 14572 9321 14600
rect 8904 14560 8910 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 11790 14600 11796 14612
rect 10827 14572 11796 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 17126 14560 17132 14612
rect 17184 14600 17190 14612
rect 17773 14603 17831 14609
rect 17773 14600 17785 14603
rect 17184 14572 17785 14600
rect 17184 14560 17190 14572
rect 17773 14569 17785 14572
rect 17819 14569 17831 14603
rect 17773 14563 17831 14569
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 20438 14600 20444 14612
rect 18923 14572 20444 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20622 14560 20628 14612
rect 20680 14600 20686 14612
rect 21910 14600 21916 14612
rect 20680 14572 20852 14600
rect 21871 14572 21916 14600
rect 20680 14560 20686 14572
rect 9122 14532 9128 14544
rect 9083 14504 9128 14532
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 17313 14535 17371 14541
rect 17313 14501 17325 14535
rect 17359 14532 17371 14535
rect 18141 14535 18199 14541
rect 17359 14504 17908 14532
rect 17359 14501 17371 14504
rect 17313 14495 17371 14501
rect 8202 14464 8208 14476
rect 6886 14436 8208 14464
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14396 4491 14399
rect 4522 14396 4528 14408
rect 4479 14368 4528 14396
rect 4479 14365 4491 14368
rect 4433 14359 4491 14365
rect 3252 14328 3280 14359
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4706 14396 4712 14408
rect 4667 14368 4712 14396
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14396 5779 14399
rect 6886 14396 6914 14436
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8570 14464 8576 14476
rect 8531 14436 8576 14464
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 9214 14424 9220 14476
rect 9272 14424 9278 14476
rect 11790 14464 11796 14476
rect 10980 14436 11796 14464
rect 5767 14368 6914 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7708 14368 7757 14396
rect 7708 14356 7714 14368
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 9232 14396 9260 14424
rect 10980 14405 11008 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 15102 14424 15108 14476
rect 15160 14464 15166 14476
rect 17880 14473 17908 14504
rect 18141 14501 18153 14535
rect 18187 14501 18199 14535
rect 18141 14495 18199 14501
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14532 19487 14535
rect 19794 14532 19800 14544
rect 19475 14504 19800 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 17865 14467 17923 14473
rect 15160 14436 15792 14464
rect 15160 14424 15166 14436
rect 15764 14408 15792 14436
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 18156 14464 18184 14495
rect 19794 14492 19800 14504
rect 19852 14492 19858 14544
rect 19334 14464 19340 14476
rect 18156 14436 19340 14464
rect 17865 14427 17923 14433
rect 8435 14368 9260 14396
rect 10965 14399 11023 14405
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 10965 14365 10977 14399
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14396 11299 14399
rect 11330 14396 11336 14408
rect 11287 14368 11336 14396
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 13078 14396 13084 14408
rect 12406 14368 13084 14396
rect 9306 14337 9312 14340
rect 5353 14331 5411 14337
rect 5353 14328 5365 14331
rect 3252 14300 5365 14328
rect 5353 14297 5365 14300
rect 5399 14297 5411 14331
rect 5353 14291 5411 14297
rect 9293 14331 9312 14337
rect 9293 14297 9305 14331
rect 9293 14291 9312 14297
rect 9306 14288 9312 14291
rect 9364 14288 9370 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9582 14328 9588 14340
rect 9539 14300 9588 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10502 14288 10508 14340
rect 10560 14328 10566 14340
rect 12406 14328 12434 14368
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13722 14396 13728 14408
rect 13683 14368 13728 14396
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 14458 14396 14464 14408
rect 14419 14368 14464 14396
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 10560 14300 12434 14328
rect 12836 14331 12894 14337
rect 10560 14288 10566 14300
rect 12836 14297 12848 14331
rect 12882 14328 12894 14331
rect 15488 14328 15516 14359
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15804 14368 15945 14396
rect 15804 14356 15810 14368
rect 15933 14365 15945 14368
rect 15979 14396 15991 14399
rect 15979 14368 17724 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16178 14331 16236 14337
rect 16178 14328 16190 14331
rect 12882 14300 13584 14328
rect 15488 14300 16190 14328
rect 12882 14297 12894 14300
rect 12836 14291 12894 14297
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 8168 14232 8217 14260
rect 8168 14220 8174 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 8205 14223 8263 14229
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11238 14260 11244 14272
rect 11195 14232 11244 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 11790 14260 11796 14272
rect 11747 14232 11796 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 13556 14269 13584 14300
rect 16178 14297 16190 14300
rect 16224 14297 16236 14331
rect 17696 14328 17724 14368
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 18708 14405 18736 14436
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 20824 14473 20852 14572
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 41417 14603 41475 14609
rect 41417 14569 41429 14603
rect 41463 14600 41475 14603
rect 41966 14600 41972 14612
rect 41463 14572 41972 14600
rect 41463 14569 41475 14572
rect 41417 14563 41475 14569
rect 41966 14560 41972 14572
rect 42024 14560 42030 14612
rect 45830 14600 45836 14612
rect 45791 14572 45836 14600
rect 45830 14560 45836 14572
rect 45888 14560 45894 14612
rect 20809 14467 20867 14473
rect 20809 14433 20821 14467
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 18693 14399 18751 14405
rect 17828 14368 17873 14396
rect 17828 14356 17834 14368
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19150 14396 19156 14408
rect 18923 14368 19156 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 21450 14396 21456 14408
rect 21411 14368 21456 14396
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22186 14396 22192 14408
rect 22143 14368 22192 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22336 14368 22381 14396
rect 22336 14356 22342 14368
rect 39942 14356 39948 14408
rect 40000 14396 40006 14408
rect 40310 14405 40316 14408
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 40000 14368 40049 14396
rect 40000 14356 40006 14368
rect 40037 14365 40049 14368
rect 40083 14365 40095 14399
rect 40304 14396 40316 14405
rect 40271 14368 40316 14396
rect 40037 14359 40095 14365
rect 40304 14359 40316 14368
rect 40310 14356 40316 14359
rect 40368 14356 40374 14408
rect 43257 14399 43315 14405
rect 43257 14365 43269 14399
rect 43303 14396 43315 14399
rect 43346 14396 43352 14408
rect 43303 14368 43352 14396
rect 43303 14365 43315 14368
rect 43257 14359 43315 14365
rect 43346 14356 43352 14368
rect 43404 14396 43410 14408
rect 43806 14396 43812 14408
rect 43404 14368 43812 14396
rect 43404 14356 43410 14368
rect 43806 14356 43812 14368
rect 43864 14356 43870 14408
rect 45186 14396 45192 14408
rect 45147 14368 45192 14396
rect 45186 14356 45192 14368
rect 45244 14356 45250 14408
rect 19978 14328 19984 14340
rect 17696 14300 19984 14328
rect 16178 14291 16236 14297
rect 19978 14288 19984 14300
rect 20036 14288 20042 14340
rect 20564 14331 20622 14337
rect 20564 14297 20576 14331
rect 20610 14328 20622 14331
rect 43524 14331 43582 14337
rect 20610 14300 21312 14328
rect 20610 14297 20622 14300
rect 20564 14291 20622 14297
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14229 13599 14263
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 13541 14223 13599 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 21284 14269 21312 14300
rect 43524 14297 43536 14331
rect 43570 14328 43582 14331
rect 43714 14328 43720 14340
rect 43570 14300 43720 14328
rect 43570 14297 43582 14300
rect 43524 14291 43582 14297
rect 43714 14288 43720 14300
rect 43772 14288 43778 14340
rect 21269 14263 21327 14269
rect 21269 14229 21281 14263
rect 21315 14229 21327 14263
rect 21269 14223 21327 14229
rect 44637 14263 44695 14269
rect 44637 14229 44649 14263
rect 44683 14260 44695 14263
rect 45278 14260 45284 14272
rect 44683 14232 45284 14260
rect 44683 14229 44695 14232
rect 44637 14223 44695 14229
rect 45278 14220 45284 14232
rect 45336 14220 45342 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 4890 14056 4896 14068
rect 4847 14028 4896 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 4890 14016 4896 14028
rect 4948 14056 4954 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 4948 14028 5365 14056
rect 4948 14016 4954 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 5353 14019 5411 14025
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5592 14028 5733 14056
rect 5592 14016 5598 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 5721 14019 5779 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8846 14056 8852 14068
rect 8807 14028 8852 14056
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12069 14059 12127 14065
rect 12069 14025 12081 14059
rect 12115 14056 12127 14059
rect 14458 14056 14464 14068
rect 12115 14028 14464 14056
rect 12115 14025 12127 14028
rect 12069 14019 12127 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 41417 14059 41475 14065
rect 20312 14028 20944 14056
rect 20312 14016 20318 14028
rect 4614 13988 4620 14000
rect 3436 13960 4620 13988
rect 3436 13929 3464 13960
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 10962 13988 10968 14000
rect 7944 13960 10968 13988
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3688 13923 3746 13929
rect 3688 13889 3700 13923
rect 3734 13920 3746 13923
rect 4246 13920 4252 13932
rect 3734 13892 4252 13920
rect 3734 13889 3746 13892
rect 3688 13883 3746 13889
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4856 13892 5273 13920
rect 4856 13880 4862 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5261 13883 5319 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 7944 13929 7972 13960
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 8110 13920 8116 13932
rect 8071 13892 8116 13920
rect 7929 13883 7987 13889
rect 7944 13852 7972 13883
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8680 13929 8708 13960
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11057 13991 11115 13997
rect 11057 13957 11069 13991
rect 11103 13988 11115 13991
rect 11330 13988 11336 14000
rect 11103 13960 11336 13988
rect 11103 13957 11115 13960
rect 11057 13951 11115 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 11701 13991 11759 13997
rect 11701 13957 11713 13991
rect 11747 13957 11759 13991
rect 11701 13951 11759 13957
rect 11917 13991 11975 13997
rect 11917 13957 11929 13991
rect 11963 13988 11975 13991
rect 12618 13988 12624 14000
rect 11963 13960 12624 13988
rect 11963 13957 11975 13960
rect 11917 13951 11975 13957
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 8849 13923 8907 13929
rect 8849 13889 8861 13923
rect 8895 13920 8907 13923
rect 9214 13920 9220 13932
rect 8895 13892 9220 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11238 13920 11244 13932
rect 11195 13892 11244 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 8018 13852 8024 13864
rect 7944 13824 8024 13852
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 10888 13852 10916 13883
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 11716 13920 11744 13951
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 13664 13991 13722 13997
rect 13664 13957 13676 13991
rect 13710 13988 13722 13991
rect 14274 13988 14280 14000
rect 13710 13960 14280 13988
rect 13710 13957 13722 13960
rect 13664 13951 13722 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14826 13948 14832 14000
rect 14884 13988 14890 14000
rect 17681 13991 17739 13997
rect 17681 13988 17693 13991
rect 14884 13960 17693 13988
rect 14884 13948 14890 13960
rect 17681 13957 17693 13960
rect 17727 13988 17739 13991
rect 18141 13991 18199 13997
rect 18141 13988 18153 13991
rect 17727 13960 18153 13988
rect 17727 13957 17739 13960
rect 17681 13951 17739 13957
rect 18141 13957 18153 13960
rect 18187 13957 18199 13991
rect 18141 13951 18199 13957
rect 19889 13991 19947 13997
rect 19889 13957 19901 13991
rect 19935 13988 19947 13991
rect 19978 13988 19984 14000
rect 19935 13960 19984 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 19978 13948 19984 13960
rect 20036 13988 20042 14000
rect 20622 13988 20628 14000
rect 20036 13960 20628 13988
rect 20036 13948 20042 13960
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 12802 13920 12808 13932
rect 11716 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 15102 13920 15108 13932
rect 13955 13892 15108 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20916 13929 20944 14028
rect 41417 14025 41429 14059
rect 41463 14056 41475 14059
rect 42150 14056 42156 14068
rect 41463 14028 42156 14056
rect 41463 14025 41475 14028
rect 41417 14019 41475 14025
rect 42150 14016 42156 14028
rect 42208 14016 42214 14068
rect 44174 14016 44180 14068
rect 44232 14056 44238 14068
rect 45741 14059 45799 14065
rect 45741 14056 45753 14059
rect 44232 14028 45753 14056
rect 44232 14016 44238 14028
rect 45741 14025 45753 14028
rect 45787 14025 45799 14059
rect 45741 14019 45799 14025
rect 40304 13991 40362 13997
rect 40304 13957 40316 13991
rect 40350 13988 40362 13991
rect 41138 13988 41144 14000
rect 40350 13960 41144 13988
rect 40350 13957 40362 13960
rect 40304 13951 40362 13957
rect 41138 13948 41144 13960
rect 41196 13948 41202 14000
rect 43708 13991 43766 13997
rect 43708 13957 43720 13991
rect 43754 13988 43766 13991
rect 45186 13988 45192 14000
rect 43754 13960 45192 13988
rect 43754 13957 43766 13960
rect 43708 13951 43766 13957
rect 45186 13948 45192 13960
rect 45244 13948 45250 14000
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20496 13892 20821 13920
rect 20496 13880 20502 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 43346 13880 43352 13932
rect 43404 13920 43410 13932
rect 43441 13923 43499 13929
rect 43441 13920 43453 13923
rect 43404 13892 43453 13920
rect 43404 13880 43410 13892
rect 43441 13889 43453 13892
rect 43487 13889 43499 13923
rect 43441 13883 43499 13889
rect 44450 13880 44456 13932
rect 44508 13920 44514 13932
rect 45281 13923 45339 13929
rect 45281 13920 45293 13923
rect 44508 13892 45293 13920
rect 44508 13880 44514 13892
rect 45281 13889 45293 13892
rect 45327 13889 45339 13923
rect 45281 13883 45339 13889
rect 45554 13880 45560 13932
rect 45612 13920 45618 13932
rect 45612 13892 45657 13920
rect 45612 13880 45618 13892
rect 11790 13852 11796 13864
rect 10888 13824 11796 13852
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20404 13824 20637 13852
rect 20404 13812 20410 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 39114 13812 39120 13864
rect 39172 13852 39178 13864
rect 39942 13852 39948 13864
rect 39172 13824 39948 13852
rect 39172 13812 39178 13824
rect 39942 13812 39948 13824
rect 40000 13852 40006 13864
rect 40037 13855 40095 13861
rect 40037 13852 40049 13855
rect 40000 13824 40049 13852
rect 40000 13812 40006 13824
rect 40037 13821 40049 13824
rect 40083 13821 40095 13855
rect 45373 13855 45431 13861
rect 45373 13852 45385 13855
rect 40037 13815 40095 13821
rect 44836 13824 45385 13852
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 44836 13793 44864 13824
rect 45373 13821 45385 13824
rect 45419 13821 45431 13855
rect 45373 13815 45431 13821
rect 44821 13787 44879 13793
rect 11296 13756 12572 13784
rect 11296 13744 11302 13756
rect 12544 13728 12572 13756
rect 44821 13753 44833 13787
rect 44867 13753 44879 13787
rect 44821 13747 44879 13753
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11756 13688 11897 13716
rect 11756 13676 11762 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 12526 13716 12532 13728
rect 12487 13688 12532 13716
rect 11885 13679 11943 13685
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 16022 13716 16028 13728
rect 15983 13688 16028 13716
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 45278 13716 45284 13728
rect 45239 13688 45284 13716
rect 45278 13676 45284 13688
rect 45336 13676 45342 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 12618 13512 12624 13524
rect 12579 13484 12624 13512
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 17126 13512 17132 13524
rect 17087 13484 17132 13512
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 19981 13515 20039 13521
rect 19981 13481 19993 13515
rect 20027 13512 20039 13515
rect 20070 13512 20076 13524
rect 20027 13484 20076 13512
rect 20027 13481 20039 13484
rect 19981 13475 20039 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20165 13515 20223 13521
rect 20165 13481 20177 13515
rect 20211 13512 20223 13515
rect 21450 13512 21456 13524
rect 20211 13484 21456 13512
rect 20211 13481 20223 13484
rect 20165 13475 20223 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 43346 13512 43352 13524
rect 42996 13484 43352 13512
rect 4157 13447 4215 13453
rect 4157 13413 4169 13447
rect 4203 13444 4215 13447
rect 5626 13444 5632 13456
rect 4203 13416 5632 13444
rect 4203 13413 4215 13416
rect 4157 13407 4215 13413
rect 5626 13404 5632 13416
rect 5684 13444 5690 13456
rect 12161 13447 12219 13453
rect 5684 13416 6592 13444
rect 5684 13404 5690 13416
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13376 4031 13379
rect 5534 13376 5540 13388
rect 4019 13348 5540 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 5534 13336 5540 13348
rect 5592 13376 5598 13388
rect 5592 13348 5672 13376
rect 5592 13336 5598 13348
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4249 13271 4307 13277
rect 4264 13240 4292 13271
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5644 13317 5672 13348
rect 6564 13317 6592 13416
rect 12161 13413 12173 13447
rect 12207 13444 12219 13447
rect 12526 13444 12532 13456
rect 12207 13416 12532 13444
rect 12207 13413 12219 13416
rect 12161 13407 12219 13413
rect 12526 13404 12532 13416
rect 12584 13444 12590 13456
rect 12894 13444 12900 13456
rect 12584 13416 12900 13444
rect 12584 13404 12590 13416
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 15746 13376 15752 13388
rect 15707 13348 15752 13376
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 42996 13385 43024 13484
rect 43346 13472 43352 13484
rect 43404 13472 43410 13524
rect 44361 13515 44419 13521
rect 44361 13481 44373 13515
rect 44407 13512 44419 13515
rect 44450 13512 44456 13524
rect 44407 13484 44456 13512
rect 44407 13481 44419 13484
rect 44361 13475 44419 13481
rect 44450 13472 44456 13484
rect 44508 13472 44514 13524
rect 42981 13379 43039 13385
rect 42981 13345 42993 13379
rect 43027 13345 43039 13379
rect 42981 13339 43039 13345
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4948 13280 5089 13308
rect 4948 13268 4954 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 6638 13308 6644 13320
rect 6595 13280 6644 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 5166 13240 5172 13252
rect 4264 13212 5172 13240
rect 5166 13200 5172 13212
rect 5224 13240 5230 13252
rect 5828 13240 5856 13271
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13308 7987 13311
rect 8110 13308 8116 13320
rect 7975 13280 8116 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8570 13308 8576 13320
rect 8251 13280 8576 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11054 13308 11060 13320
rect 11011 13280 11060 13308
rect 11011 13277 11023 13280
rect 10965 13271 11023 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 16022 13317 16028 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12406 13280 13001 13308
rect 8018 13240 8024 13252
rect 5224 13212 5856 13240
rect 7979 13212 8024 13240
rect 5224 13200 5230 13212
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 11388 13212 11989 13240
rect 11388 13200 11394 13212
rect 11977 13209 11989 13212
rect 12023 13240 12035 13243
rect 12250 13240 12256 13252
rect 12023 13212 12256 13240
rect 12023 13209 12035 13212
rect 11977 13203 12035 13209
rect 12250 13200 12256 13212
rect 12308 13240 12314 13252
rect 12406 13240 12434 13280
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 16016 13308 16028 13317
rect 15983 13280 16028 13308
rect 12989 13271 13047 13277
rect 16016 13271 16028 13280
rect 16022 13268 16028 13271
rect 16080 13268 16086 13320
rect 20438 13308 20444 13320
rect 19812 13280 20444 13308
rect 12308 13212 12434 13240
rect 12805 13243 12863 13249
rect 12308 13200 12314 13212
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 12894 13240 12900 13252
rect 12851 13212 12900 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 19812 13249 19840 13280
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 40034 13308 40040 13320
rect 39995 13280 40040 13308
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 19797 13243 19855 13249
rect 19797 13209 19809 13243
rect 19843 13209 19855 13243
rect 19797 13203 19855 13209
rect 20013 13243 20071 13249
rect 20013 13209 20025 13243
rect 20059 13240 20071 13243
rect 20530 13240 20536 13252
rect 20059 13212 20536 13240
rect 20059 13209 20071 13212
rect 20013 13203 20071 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 43254 13249 43260 13252
rect 43248 13203 43260 13249
rect 43312 13240 43318 13252
rect 43312 13212 43348 13240
rect 43254 13200 43260 13203
rect 43312 13200 43318 13212
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 4982 13172 4988 13184
rect 4295 13144 4988 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 8202 13172 8208 13184
rect 6595 13144 8208 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 11020 13144 11621 13172
rect 11020 13132 11026 13144
rect 11609 13141 11621 13144
rect 11655 13141 11667 13175
rect 11790 13172 11796 13184
rect 11751 13144 11796 13172
rect 11609 13135 11667 13141
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 11940 13144 11985 13172
rect 11940 13132 11946 13144
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5166 12968 5172 12980
rect 5092 12940 5172 12968
rect 4798 12832 4804 12844
rect 4711 12804 4804 12832
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 5092 12841 5120 12940
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 7403 12971 7461 12977
rect 7403 12937 7415 12971
rect 7449 12968 7461 12971
rect 8110 12968 8116 12980
rect 7449 12940 8116 12968
rect 7449 12937 7461 12940
rect 7403 12931 7461 12937
rect 8110 12928 8116 12940
rect 8168 12968 8174 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 8168 12940 8309 12968
rect 8168 12928 8174 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 11054 12968 11060 12980
rect 11015 12940 11060 12968
rect 8297 12931 8355 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12937 11759 12971
rect 12802 12968 12808 12980
rect 12763 12940 12808 12968
rect 11701 12931 11759 12937
rect 7193 12903 7251 12909
rect 7193 12869 7205 12903
rect 7239 12900 7251 12903
rect 8665 12903 8723 12909
rect 7239 12872 8524 12900
rect 7239 12869 7251 12872
rect 7193 12863 7251 12869
rect 5169 12841 5227 12847
rect 5077 12835 5135 12841
rect 4948 12804 4993 12832
rect 4948 12792 4954 12804
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5169 12807 5181 12841
rect 5215 12832 5227 12841
rect 5626 12832 5632 12844
rect 5215 12807 5632 12832
rect 5169 12804 5632 12807
rect 5169 12801 5227 12804
rect 5077 12795 5135 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 8018 12832 8024 12844
rect 7432 12804 8024 12832
rect 7432 12792 7438 12804
rect 8018 12792 8024 12804
rect 8076 12832 8082 12844
rect 8496 12841 8524 12872
rect 8665 12869 8677 12903
rect 8711 12900 8723 12903
rect 9030 12900 9036 12912
rect 8711 12872 9036 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 9030 12860 9036 12872
rect 9088 12900 9094 12912
rect 9309 12903 9367 12909
rect 9309 12900 9321 12903
rect 9088 12872 9321 12900
rect 9088 12860 9094 12872
rect 9309 12869 9321 12872
rect 9355 12869 9367 12903
rect 9309 12863 9367 12869
rect 10873 12903 10931 12909
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 11716 12900 11744 12931
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 43254 12968 43260 12980
rect 43215 12940 43260 12968
rect 43254 12928 43260 12940
rect 43312 12928 43318 12980
rect 43901 12971 43959 12977
rect 43901 12937 43913 12971
rect 43947 12968 43959 12971
rect 45278 12968 45284 12980
rect 43947 12940 45284 12968
rect 43947 12937 43959 12940
rect 43901 12931 43959 12937
rect 45278 12928 45284 12940
rect 45336 12928 45342 12980
rect 10919 12872 11744 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 11882 12860 11888 12912
rect 11940 12860 11946 12912
rect 39384 12903 39442 12909
rect 39384 12869 39396 12903
rect 39430 12900 39442 12903
rect 40034 12900 40040 12912
rect 39430 12872 40040 12900
rect 39430 12869 39442 12872
rect 39384 12863 39442 12869
rect 40034 12860 40040 12872
rect 40092 12860 40098 12912
rect 43349 12903 43407 12909
rect 43349 12869 43361 12903
rect 43395 12900 43407 12903
rect 43806 12900 43812 12912
rect 43395 12872 43812 12900
rect 43395 12869 43407 12872
rect 43349 12863 43407 12869
rect 43806 12860 43812 12872
rect 43864 12860 43870 12912
rect 44174 12900 44180 12912
rect 44135 12872 44180 12900
rect 44174 12860 44180 12872
rect 44232 12860 44238 12912
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8076 12804 8401 12832
rect 8076 12792 8082 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 8570 12832 8576 12844
rect 8527 12804 8576 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 10505 12835 10563 12841
rect 9171 12804 9260 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 4816 12764 4844 12792
rect 4816 12736 7512 12764
rect 7374 12628 7380 12640
rect 7335 12600 7380 12628
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 7484 12628 7512 12736
rect 7561 12699 7619 12705
rect 7561 12665 7573 12699
rect 7607 12696 7619 12699
rect 9232 12696 9260 12804
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10962 12832 10968 12844
rect 10551 12804 10968 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11900 12832 11928 12860
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11900 12804 12173 12832
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 12713 12835 12771 12841
rect 12713 12832 12725 12835
rect 12308 12804 12725 12832
rect 12308 12792 12314 12804
rect 12713 12801 12725 12804
rect 12759 12801 12771 12835
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 12713 12795 12771 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 42981 12835 43039 12841
rect 42981 12801 42993 12835
rect 43027 12832 43039 12835
rect 44192 12832 44220 12860
rect 43027 12804 44220 12832
rect 43027 12801 43039 12804
rect 42981 12795 43039 12801
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11848 12736 11897 12764
rect 11848 12724 11854 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12912 12764 12940 12792
rect 39114 12764 39120 12776
rect 12115 12736 12940 12764
rect 39075 12736 39120 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 9398 12696 9404 12708
rect 7607 12668 9404 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 11992 12696 12020 12727
rect 39114 12724 39120 12736
rect 39172 12724 39178 12776
rect 12250 12696 12256 12708
rect 11992 12668 12256 12696
rect 12250 12656 12256 12668
rect 12308 12656 12314 12708
rect 44085 12699 44143 12705
rect 44085 12696 44097 12699
rect 43088 12668 44097 12696
rect 43088 12640 43116 12668
rect 44085 12665 44097 12668
rect 44131 12665 44143 12699
rect 44085 12659 44143 12665
rect 7742 12628 7748 12640
rect 7484 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12628 7806 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7800 12600 8125 12628
rect 7800 12588 7806 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 8113 12591 8171 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 9640 12600 10885 12628
rect 9640 12588 9646 12600
rect 10873 12597 10885 12600
rect 10919 12628 10931 12631
rect 11790 12628 11796 12640
rect 10919 12600 11796 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 40497 12631 40555 12637
rect 40497 12597 40509 12631
rect 40543 12628 40555 12631
rect 40862 12628 40868 12640
rect 40543 12600 40868 12628
rect 40543 12597 40555 12600
rect 40497 12591 40555 12597
rect 40862 12588 40868 12600
rect 40920 12588 40926 12640
rect 43070 12628 43076 12640
rect 43031 12600 43076 12628
rect 43070 12588 43076 12600
rect 43128 12588 43134 12640
rect 43165 12631 43223 12637
rect 43165 12597 43177 12631
rect 43211 12628 43223 12631
rect 43993 12631 44051 12637
rect 43993 12628 44005 12631
rect 43211 12600 44005 12628
rect 43211 12597 43223 12600
rect 43165 12591 43223 12597
rect 43993 12597 44005 12600
rect 44039 12628 44051 12631
rect 44450 12628 44456 12640
rect 44039 12600 44456 12628
rect 44039 12597 44051 12600
rect 43993 12591 44051 12597
rect 44450 12588 44456 12600
rect 44508 12588 44514 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 8570 12424 8576 12436
rect 8531 12396 8576 12424
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 9582 12424 9588 12436
rect 9355 12396 9588 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 9324 12356 9352 12387
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 8260 12328 9352 12356
rect 8260 12316 8266 12328
rect 9398 12316 9404 12368
rect 9456 12356 9462 12368
rect 9677 12359 9735 12365
rect 9677 12356 9689 12359
rect 9456 12328 9689 12356
rect 9456 12316 9462 12328
rect 9677 12325 9689 12328
rect 9723 12325 9735 12359
rect 9677 12319 9735 12325
rect 3970 12220 3976 12232
rect 3931 12192 3976 12220
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 5500 12192 7205 12220
rect 5500 12180 5506 12192
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 7742 12220 7748 12232
rect 7239 12192 7748 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10778 12229 10784 12232
rect 10772 12183 10784 12229
rect 10836 12220 10842 12232
rect 38838 12220 38844 12232
rect 10836 12192 10872 12220
rect 38799 12192 38844 12220
rect 10778 12180 10784 12183
rect 10836 12180 10842 12192
rect 38838 12180 38844 12192
rect 38896 12180 38902 12232
rect 39298 12220 39304 12232
rect 39259 12192 39304 12220
rect 39298 12180 39304 12192
rect 39356 12180 39362 12232
rect 42886 12220 42892 12232
rect 42847 12192 42892 12220
rect 42886 12180 42892 12192
rect 42944 12180 42950 12232
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7438 12155 7496 12161
rect 7438 12152 7450 12155
rect 7340 12124 7450 12152
rect 7340 12112 7346 12124
rect 7438 12121 7450 12124
rect 7484 12121 7496 12155
rect 7438 12115 7496 12121
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 8444 12124 9321 12152
rect 8444 12112 8450 12124
rect 9309 12121 9321 12124
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 7156 12056 9137 12084
rect 7156 12044 7162 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 41598 12084 41604 12096
rect 41559 12056 41604 12084
rect 9125 12047 9183 12053
rect 41598 12044 41604 12056
rect 41656 12044 41662 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 9088 11852 9137 11880
rect 9088 11840 9094 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11849 9643 11883
rect 9585 11843 9643 11849
rect 41325 11883 41383 11889
rect 41325 11849 41337 11883
rect 41371 11880 41383 11883
rect 43070 11880 43076 11892
rect 41371 11852 43076 11880
rect 41371 11849 41383 11852
rect 41325 11843 41383 11849
rect 8012 11815 8070 11821
rect 8012 11781 8024 11815
rect 8058 11812 8070 11815
rect 9600 11812 9628 11843
rect 43070 11840 43076 11852
rect 43128 11840 43134 11892
rect 8058 11784 9628 11812
rect 12161 11815 12219 11821
rect 8058 11781 8070 11784
rect 8012 11775 8070 11781
rect 12161 11781 12173 11815
rect 12207 11812 12219 11815
rect 12250 11812 12256 11824
rect 12207 11784 12256 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 39298 11821 39304 11824
rect 39292 11812 39304 11821
rect 39259 11784 39304 11812
rect 39292 11775 39304 11784
rect 39298 11772 39304 11775
rect 39356 11772 39362 11824
rect 2952 11747 3010 11753
rect 2952 11713 2964 11747
rect 2998 11744 3010 11747
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 2998 11716 4629 11744
rect 2998 11713 3010 11716
rect 2952 11707 3010 11713
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 7098 11744 7104 11756
rect 7059 11716 7104 11744
rect 4617 11707 4675 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 9766 11744 9772 11756
rect 9727 11716 9772 11744
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 39025 11747 39083 11753
rect 39025 11713 39037 11747
rect 39071 11744 39083 11747
rect 39114 11744 39120 11756
rect 39071 11716 39120 11744
rect 39071 11713 39083 11716
rect 39025 11707 39083 11713
rect 39114 11704 39120 11716
rect 39172 11704 39178 11756
rect 39574 11704 39580 11756
rect 39632 11744 39638 11756
rect 40865 11747 40923 11753
rect 40865 11744 40877 11747
rect 39632 11716 40877 11744
rect 39632 11704 39638 11716
rect 40865 11713 40877 11716
rect 40911 11713 40923 11747
rect 40865 11707 40923 11713
rect 41141 11747 41199 11753
rect 41141 11713 41153 11747
rect 41187 11744 41199 11747
rect 41414 11744 41420 11756
rect 41187 11716 41420 11744
rect 41187 11713 41199 11716
rect 41141 11707 41199 11713
rect 41414 11704 41420 11716
rect 41472 11704 41478 11756
rect 2682 11676 2688 11688
rect 2643 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 40957 11679 41015 11685
rect 40957 11645 40969 11679
rect 41003 11645 41015 11679
rect 40957 11639 41015 11645
rect 4065 11611 4123 11617
rect 4065 11577 4077 11611
rect 4111 11608 4123 11611
rect 4706 11608 4712 11620
rect 4111 11580 4712 11608
rect 4111 11577 4123 11580
rect 4065 11571 4123 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 11790 11608 11796 11620
rect 11751 11580 11796 11608
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 40405 11611 40463 11617
rect 40405 11577 40417 11611
rect 40451 11608 40463 11611
rect 40972 11608 41000 11639
rect 40451 11580 41000 11608
rect 40451 11577 40463 11580
rect 40405 11571 40463 11577
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 11882 11540 11888 11552
rect 11747 11512 11888 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 38378 11540 38384 11552
rect 38339 11512 38384 11540
rect 38378 11500 38384 11512
rect 38436 11500 38442 11552
rect 40862 11540 40868 11552
rect 40823 11512 40868 11540
rect 40862 11500 40868 11512
rect 40920 11500 40926 11552
rect 42426 11500 42432 11552
rect 42484 11540 42490 11552
rect 42613 11543 42671 11549
rect 42613 11540 42625 11543
rect 42484 11512 42625 11540
rect 42484 11500 42490 11512
rect 42613 11509 42625 11512
rect 42659 11509 42671 11543
rect 42613 11503 42671 11509
rect 43441 11543 43499 11549
rect 43441 11509 43453 11543
rect 43487 11540 43499 11543
rect 44726 11540 44732 11552
rect 43487 11512 44732 11540
rect 43487 11509 43499 11512
rect 43441 11503 43499 11509
rect 44726 11500 44732 11512
rect 44784 11500 44790 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12308 11308 12725 11336
rect 12308 11296 12314 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 12713 11299 12771 11305
rect 39485 11339 39543 11345
rect 39485 11305 39497 11339
rect 39531 11336 39543 11339
rect 39574 11336 39580 11348
rect 39531 11308 39580 11336
rect 39531 11305 39543 11308
rect 39485 11299 39543 11305
rect 39574 11296 39580 11308
rect 39632 11296 39638 11348
rect 41414 11336 41420 11348
rect 41375 11308 41420 11336
rect 41414 11296 41420 11308
rect 41472 11296 41478 11348
rect 43533 11339 43591 11345
rect 43533 11305 43545 11339
rect 43579 11336 43591 11339
rect 43993 11339 44051 11345
rect 43993 11336 44005 11339
rect 43579 11308 44005 11336
rect 43579 11305 43591 11308
rect 43533 11299 43591 11305
rect 43993 11305 44005 11308
rect 44039 11305 44051 11339
rect 44450 11336 44456 11348
rect 44411 11308 44456 11336
rect 43993 11299 44051 11305
rect 44450 11296 44456 11308
rect 44508 11296 44514 11348
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 5500 11172 6561 11200
rect 5500 11160 5506 11172
rect 6549 11169 6561 11172
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 10560 11172 11345 11200
rect 10560 11160 10566 11172
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2682 11132 2688 11144
rect 1995 11104 2688 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6454 11132 6460 11144
rect 6135 11104 6460 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 20346 11132 20352 11144
rect 20307 11104 20352 11132
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 38105 11135 38163 11141
rect 38105 11101 38117 11135
rect 38151 11132 38163 11135
rect 39114 11132 39120 11144
rect 38151 11104 39120 11132
rect 38151 11101 38163 11104
rect 38105 11095 38163 11101
rect 39114 11092 39120 11104
rect 39172 11132 39178 11144
rect 40037 11135 40095 11141
rect 40037 11132 40049 11135
rect 39172 11104 40049 11132
rect 39172 11092 39178 11104
rect 40037 11101 40049 11104
rect 40083 11132 40095 11135
rect 41598 11132 41604 11144
rect 40083 11104 41604 11132
rect 40083 11101 40095 11104
rect 40037 11095 40095 11101
rect 41598 11092 41604 11104
rect 41656 11132 41662 11144
rect 42153 11135 42211 11141
rect 42153 11132 42165 11135
rect 41656 11104 42165 11132
rect 41656 11092 41662 11104
rect 42153 11101 42165 11104
rect 42199 11132 42211 11135
rect 44174 11132 44180 11144
rect 42199 11104 42564 11132
rect 44135 11104 44180 11132
rect 42199 11101 42211 11104
rect 42153 11095 42211 11101
rect 42536 11076 42564 11104
rect 44174 11092 44180 11104
rect 44232 11092 44238 11144
rect 44269 11135 44327 11141
rect 44269 11101 44281 11135
rect 44315 11132 44327 11135
rect 45830 11132 45836 11144
rect 44315 11104 45836 11132
rect 44315 11101 44327 11104
rect 44269 11095 44327 11101
rect 45830 11092 45836 11104
rect 45888 11092 45894 11144
rect 2222 11073 2228 11076
rect 2216 11064 2228 11073
rect 2183 11036 2228 11064
rect 2216 11027 2228 11036
rect 2222 11024 2228 11027
rect 2280 11024 2286 11076
rect 4338 11064 4344 11076
rect 4299 11036 4344 11064
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 6794 11067 6852 11073
rect 6794 11064 6806 11067
rect 5868 11036 6806 11064
rect 5868 11024 5874 11036
rect 6794 11033 6806 11036
rect 6840 11033 6852 11067
rect 6794 11027 6852 11033
rect 11600 11067 11658 11073
rect 11600 11033 11612 11067
rect 11646 11064 11658 11067
rect 11698 11064 11704 11076
rect 11646 11036 11704 11064
rect 11646 11033 11658 11036
rect 11600 11027 11658 11033
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 38378 11073 38384 11076
rect 38372 11064 38384 11073
rect 38339 11036 38384 11064
rect 38372 11027 38384 11036
rect 38378 11024 38384 11027
rect 38436 11024 38442 11076
rect 38838 11024 38844 11076
rect 38896 11064 38902 11076
rect 42426 11073 42432 11076
rect 40282 11067 40340 11073
rect 40282 11064 40294 11067
rect 38896 11036 40294 11064
rect 38896 11024 38902 11036
rect 40282 11033 40294 11036
rect 40328 11033 40340 11067
rect 42420 11064 42432 11073
rect 42387 11036 42432 11064
rect 40282 11027 40340 11033
rect 42420 11027 42432 11036
rect 42426 11024 42432 11027
rect 42484 11024 42490 11076
rect 42518 11024 42524 11076
rect 42576 11024 42582 11076
rect 43990 11064 43996 11076
rect 43951 11036 43996 11064
rect 43990 11024 43996 11036
rect 44048 11024 44054 11076
rect 3326 10996 3332 11008
rect 3287 10968 3332 10996
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7929 10999 7987 11005
rect 7929 10996 7941 10999
rect 6972 10968 7941 10996
rect 6972 10956 6978 10968
rect 7929 10965 7941 10968
rect 7975 10965 7987 10999
rect 7929 10959 7987 10965
rect 20165 10999 20223 11005
rect 20165 10965 20177 10999
rect 20211 10996 20223 10999
rect 20254 10996 20260 11008
rect 20211 10968 20260 10996
rect 20211 10965 20223 10968
rect 20165 10959 20223 10965
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 9766 10792 9772 10804
rect 8343 10764 9772 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 11698 10792 11704 10804
rect 11659 10764 11704 10792
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 43990 10792 43996 10804
rect 43951 10764 43996 10792
rect 43990 10752 43996 10764
rect 44048 10752 44054 10804
rect 45830 10792 45836 10804
rect 45791 10764 45836 10792
rect 45830 10752 45836 10764
rect 45888 10752 45894 10804
rect 4338 10724 4344 10736
rect 1596 10696 2728 10724
rect 1596 10665 1624 10696
rect 2700 10668 2728 10696
rect 3436 10696 4344 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 1848 10659 1906 10665
rect 1848 10625 1860 10659
rect 1894 10656 1906 10659
rect 1894 10628 2636 10656
rect 1894 10625 1906 10628
rect 1848 10619 1906 10625
rect 2608 10588 2636 10628
rect 2682 10616 2688 10668
rect 2740 10656 2746 10668
rect 3436 10665 3464 10696
rect 4338 10684 4344 10696
rect 4396 10724 4402 10736
rect 5442 10724 5448 10736
rect 4396 10696 5448 10724
rect 4396 10684 4402 10696
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 9490 10724 9496 10736
rect 8159 10696 9496 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 44726 10733 44732 10736
rect 44720 10724 44732 10733
rect 42628 10696 44496 10724
rect 44687 10696 44732 10724
rect 3421 10659 3479 10665
rect 3421 10656 3433 10659
rect 2740 10628 3433 10656
rect 2740 10616 2746 10628
rect 3421 10625 3433 10628
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 3688 10659 3746 10665
rect 3688 10625 3700 10659
rect 3734 10656 3746 10659
rect 3970 10656 3976 10668
rect 3734 10628 3976 10656
rect 3734 10625 3746 10628
rect 3688 10619 3746 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 2774 10588 2780 10600
rect 2608 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 7024 10588 7052 10619
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7708 10628 7757 10656
rect 7708 10616 7714 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 11882 10656 11888 10668
rect 11843 10628 11888 10656
rect 7745 10619 7803 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 40126 10656 40132 10668
rect 40087 10628 40132 10656
rect 40126 10616 40132 10628
rect 40184 10616 40190 10668
rect 42518 10616 42524 10668
rect 42576 10656 42582 10668
rect 42628 10665 42656 10696
rect 42613 10659 42671 10665
rect 42613 10656 42625 10659
rect 42576 10628 42625 10656
rect 42576 10616 42582 10628
rect 42613 10625 42625 10628
rect 42659 10625 42671 10659
rect 42869 10659 42927 10665
rect 42869 10656 42881 10659
rect 42613 10619 42671 10625
rect 42720 10628 42881 10656
rect 4672 10560 7052 10588
rect 42061 10591 42119 10597
rect 4672 10548 4678 10560
rect 42061 10557 42073 10591
rect 42107 10588 42119 10591
rect 42720 10588 42748 10628
rect 42869 10625 42881 10628
rect 42915 10625 42927 10659
rect 42869 10619 42927 10625
rect 44468 10600 44496 10696
rect 44720 10687 44732 10696
rect 44726 10684 44732 10687
rect 44784 10684 44790 10736
rect 44450 10588 44456 10600
rect 42107 10560 42748 10588
rect 44411 10560 44456 10588
rect 42107 10557 42119 10560
rect 42061 10551 42119 10557
rect 44450 10548 44456 10560
rect 44508 10548 44514 10600
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 4062 10452 4068 10464
rect 3007 10424 4068 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 8113 10455 8171 10461
rect 8113 10421 8125 10455
rect 8159 10452 8171 10455
rect 8202 10452 8208 10464
rect 8159 10424 8208 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 40313 10455 40371 10461
rect 40313 10421 40325 10455
rect 40359 10452 40371 10455
rect 40586 10452 40592 10464
rect 40359 10424 40592 10452
rect 40359 10421 40371 10424
rect 40313 10415 40371 10421
rect 40586 10412 40592 10424
rect 40644 10412 40650 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 4062 10248 4068 10260
rect 2740 10220 3004 10248
rect 4023 10220 4068 10248
rect 2740 10208 2746 10220
rect 2976 10121 3004 10220
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 4614 10248 4620 10260
rect 4571 10220 4620 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 43901 10251 43959 10257
rect 43901 10217 43913 10251
rect 43947 10248 43959 10251
rect 44174 10248 44180 10260
rect 43947 10220 44180 10248
rect 43947 10217 43959 10220
rect 43901 10211 43959 10217
rect 44174 10208 44180 10220
rect 44232 10208 44238 10260
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10081 3019 10115
rect 2961 10075 3019 10081
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 4706 10112 4712 10124
rect 4295 10084 4712 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 42518 10112 42524 10124
rect 42479 10084 42524 10112
rect 42518 10072 42524 10084
rect 42576 10072 42582 10124
rect 44450 10072 44456 10124
rect 44508 10112 44514 10124
rect 45189 10115 45247 10121
rect 45189 10112 45201 10115
rect 44508 10084 45201 10112
rect 44508 10072 44514 10084
rect 45189 10081 45201 10084
rect 45235 10081 45247 10115
rect 45189 10075 45247 10081
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3384 10016 4077 10044
rect 3384 10004 3390 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4798 10044 4804 10056
rect 4387 10016 4804 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 5718 10053 5724 10056
rect 5712 10044 5724 10053
rect 5679 10016 5724 10044
rect 5712 10007 5724 10016
rect 5718 10004 5724 10007
rect 5776 10004 5782 10056
rect 20254 10053 20260 10056
rect 20248 10044 20260 10053
rect 20215 10016 20260 10044
rect 20248 10007 20260 10016
rect 20254 10004 20260 10007
rect 20312 10004 20318 10056
rect 45278 10004 45284 10056
rect 45336 10044 45342 10056
rect 45445 10047 45503 10053
rect 45445 10044 45457 10047
rect 45336 10016 45457 10044
rect 45336 10004 45342 10016
rect 45445 10013 45457 10016
rect 45491 10013 45503 10047
rect 45445 10007 45503 10013
rect 2716 9979 2774 9985
rect 2716 9945 2728 9979
rect 2762 9976 2774 9979
rect 4982 9976 4988 9988
rect 2762 9948 4988 9976
rect 2762 9945 2774 9948
rect 2716 9939 2774 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 42794 9985 42800 9988
rect 42788 9939 42800 9985
rect 42852 9976 42858 9988
rect 42852 9948 42888 9976
rect 42794 9936 42800 9939
rect 42852 9936 42858 9948
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1854 9908 1860 9920
rect 1627 9880 1860 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 21361 9911 21419 9917
rect 21361 9877 21373 9911
rect 21407 9908 21419 9911
rect 22002 9908 22008 9920
rect 21407 9880 22008 9908
rect 21407 9877 21419 9880
rect 21361 9871 21419 9877
rect 22002 9868 22008 9880
rect 22060 9868 22066 9920
rect 46569 9911 46627 9917
rect 46569 9877 46581 9911
rect 46615 9908 46627 9911
rect 57514 9908 57520 9920
rect 46615 9880 57520 9908
rect 46615 9877 46627 9880
rect 46569 9871 46627 9877
rect 57514 9868 57520 9880
rect 57572 9868 57578 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 42518 9636 42524 9648
rect 40512 9608 42524 9636
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 5721 9571 5779 9577
rect 2832 9540 2877 9568
rect 2832 9528 2838 9540
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 5810 9568 5816 9580
rect 5767 9540 5816 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 40512 9577 40540 9608
rect 42518 9596 42524 9608
rect 42576 9596 42582 9648
rect 40497 9571 40555 9577
rect 40497 9537 40509 9571
rect 40543 9537 40555 9571
rect 40497 9531 40555 9537
rect 40586 9528 40592 9580
rect 40644 9568 40650 9580
rect 40753 9571 40811 9577
rect 40753 9568 40765 9571
rect 40644 9540 40765 9568
rect 40644 9528 40650 9540
rect 40753 9537 40765 9540
rect 40799 9537 40811 9571
rect 42794 9568 42800 9580
rect 42755 9540 42800 9568
rect 40753 9531 40811 9537
rect 42794 9528 42800 9540
rect 42852 9528 42858 9580
rect 41877 9367 41935 9373
rect 41877 9333 41889 9367
rect 41923 9364 41935 9367
rect 42610 9364 42616 9376
rect 41923 9336 42616 9364
rect 41923 9333 41935 9336
rect 41877 9327 41935 9333
rect 42610 9324 42616 9336
rect 42668 9324 42674 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 57514 3720 57520 3732
rect 57475 3692 57520 3720
rect 57514 3680 57520 3692
rect 57572 3680 57578 3732
rect 57514 3476 57520 3528
rect 57572 3516 57578 3528
rect 58069 3519 58127 3525
rect 58069 3516 58081 3519
rect 57572 3488 58081 3516
rect 57572 3476 57578 3488
rect 58069 3485 58081 3488
rect 58115 3485 58127 3519
rect 58069 3479 58127 3485
rect 58250 3380 58256 3392
rect 58211 3352 58256 3380
rect 58250 3340 58256 3352
rect 58308 3340 58314 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1854 2428 1860 2440
rect 1815 2400 1860 2428
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 42610 2428 42616 2440
rect 42571 2400 42616 2428
rect 42610 2388 42616 2400
rect 42668 2388 42674 2440
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21324 2264 22201 2292
rect 21324 2252 21330 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 42518 2252 42524 2304
rect 42576 2292 42582 2304
rect 42797 2295 42855 2301
rect 42797 2292 42809 2295
rect 42576 2264 42809 2292
rect 42576 2252 42582 2264
rect 42797 2261 42809 2264
rect 42843 2261 42855 2295
rect 42797 2255 42855 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 6460 57536 6512 57588
rect 28356 57536 28408 57588
rect 49700 57536 49752 57588
rect 6644 57400 6696 57452
rect 28540 57400 28592 57452
rect 46572 57400 46624 57452
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 45560 49172 45612 49224
rect 58256 49079 58308 49088
rect 58256 49045 58265 49079
rect 58265 49045 58299 49079
rect 58299 49045 58308 49079
rect 58256 49036 58308 49045
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 6644 46155 6696 46164
rect 6644 46121 6653 46155
rect 6653 46121 6687 46155
rect 6687 46121 6696 46155
rect 6644 46112 6696 46121
rect 46572 46155 46624 46164
rect 46572 46121 46581 46155
rect 46581 46121 46615 46155
rect 46615 46121 46624 46155
rect 46572 46112 46624 46121
rect 6736 45908 6788 45960
rect 40500 45951 40552 45960
rect 40500 45917 40509 45951
rect 40509 45917 40543 45951
rect 40543 45917 40552 45951
rect 40500 45908 40552 45917
rect 44272 45908 44324 45960
rect 5816 45840 5868 45892
rect 45836 45840 45888 45892
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 5816 45611 5868 45620
rect 5816 45577 5825 45611
rect 5825 45577 5859 45611
rect 5859 45577 5868 45611
rect 5816 45568 5868 45577
rect 9128 45500 9180 45552
rect 7104 45432 7156 45484
rect 8300 45432 8352 45484
rect 9680 45475 9732 45484
rect 9680 45441 9689 45475
rect 9689 45441 9723 45475
rect 9723 45441 9732 45475
rect 9680 45432 9732 45441
rect 29000 45500 29052 45552
rect 40500 45500 40552 45552
rect 27252 45432 27304 45484
rect 44272 45432 44324 45484
rect 44456 45475 44508 45484
rect 44456 45441 44490 45475
rect 44490 45441 44508 45475
rect 44456 45432 44508 45441
rect 7380 45364 7432 45416
rect 40132 45407 40184 45416
rect 6736 45296 6788 45348
rect 6920 45296 6972 45348
rect 40132 45373 40141 45407
rect 40141 45373 40175 45407
rect 40175 45373 40184 45407
rect 40132 45364 40184 45373
rect 28540 45339 28592 45348
rect 28540 45305 28549 45339
rect 28549 45305 28583 45339
rect 28583 45305 28592 45339
rect 28540 45296 28592 45305
rect 45560 45339 45612 45348
rect 45560 45305 45569 45339
rect 45569 45305 45603 45339
rect 45603 45305 45612 45339
rect 45560 45296 45612 45305
rect 6460 45228 6512 45280
rect 7656 45228 7708 45280
rect 37740 45228 37792 45280
rect 41512 45271 41564 45280
rect 41512 45237 41521 45271
rect 41521 45237 41555 45271
rect 41555 45237 41564 45271
rect 41512 45228 41564 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 7656 45067 7708 45076
rect 7656 45033 7665 45067
rect 7665 45033 7699 45067
rect 7699 45033 7708 45067
rect 7656 45024 7708 45033
rect 8300 45067 8352 45076
rect 8300 45033 8309 45067
rect 8309 45033 8343 45067
rect 8343 45033 8352 45067
rect 8300 45024 8352 45033
rect 9036 45024 9088 45076
rect 45836 45067 45888 45076
rect 6736 44931 6788 44940
rect 6736 44897 6745 44931
rect 6745 44897 6779 44931
rect 6779 44897 6788 44931
rect 6736 44888 6788 44897
rect 45836 45033 45845 45067
rect 45845 45033 45879 45067
rect 45879 45033 45888 45067
rect 45836 45024 45888 45033
rect 10784 44999 10836 45008
rect 10784 44965 10793 44999
rect 10793 44965 10827 44999
rect 10827 44965 10836 44999
rect 10784 44956 10836 44965
rect 44364 44956 44416 45008
rect 6460 44863 6512 44872
rect 6460 44829 6478 44863
rect 6478 44829 6512 44863
rect 6460 44820 6512 44829
rect 6828 44820 6880 44872
rect 7288 44863 7340 44872
rect 7288 44829 7297 44863
rect 7297 44829 7331 44863
rect 7331 44829 7340 44863
rect 7288 44820 7340 44829
rect 5908 44684 5960 44736
rect 7012 44684 7064 44736
rect 9680 44727 9732 44736
rect 9680 44693 9689 44727
rect 9689 44693 9723 44727
rect 9723 44693 9732 44727
rect 9680 44684 9732 44693
rect 11152 44820 11204 44872
rect 40132 44820 40184 44872
rect 41052 44820 41104 44872
rect 10048 44795 10100 44804
rect 10048 44761 10057 44795
rect 10057 44761 10091 44795
rect 10091 44761 10100 44795
rect 10048 44752 10100 44761
rect 36268 44752 36320 44804
rect 37280 44752 37332 44804
rect 43996 44752 44048 44804
rect 45468 44820 45520 44872
rect 45560 44752 45612 44804
rect 9956 44684 10008 44736
rect 38476 44684 38528 44736
rect 42156 44684 42208 44736
rect 43168 44727 43220 44736
rect 43168 44693 43177 44727
rect 43177 44693 43211 44727
rect 43211 44693 43220 44727
rect 43168 44684 43220 44693
rect 45192 44727 45244 44736
rect 45192 44693 45201 44727
rect 45201 44693 45235 44727
rect 45235 44693 45244 44727
rect 45192 44684 45244 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 7104 44523 7156 44532
rect 7104 44489 7113 44523
rect 7113 44489 7147 44523
rect 7147 44489 7156 44523
rect 7104 44480 7156 44489
rect 9128 44523 9180 44532
rect 9128 44489 9137 44523
rect 9137 44489 9171 44523
rect 9171 44489 9180 44523
rect 9128 44480 9180 44489
rect 9956 44480 10008 44532
rect 11152 44523 11204 44532
rect 11152 44489 11161 44523
rect 11161 44489 11195 44523
rect 11195 44489 11204 44523
rect 11152 44480 11204 44489
rect 45468 44523 45520 44532
rect 45468 44489 45477 44523
rect 45477 44489 45511 44523
rect 45511 44489 45520 44523
rect 45468 44480 45520 44489
rect 7012 44412 7064 44464
rect 7288 44412 7340 44464
rect 9036 44455 9088 44464
rect 9036 44421 9045 44455
rect 9045 44421 9079 44455
rect 9079 44421 9088 44455
rect 9036 44412 9088 44421
rect 5908 44387 5960 44396
rect 5908 44353 5917 44387
rect 5917 44353 5951 44387
rect 5951 44353 5960 44387
rect 5908 44344 5960 44353
rect 9680 44344 9732 44396
rect 36268 44387 36320 44396
rect 36268 44353 36277 44387
rect 36277 44353 36311 44387
rect 36311 44353 36320 44387
rect 36268 44344 36320 44353
rect 37740 44387 37792 44396
rect 37740 44353 37774 44387
rect 37774 44353 37792 44387
rect 37740 44344 37792 44353
rect 40132 44344 40184 44396
rect 44548 44387 44600 44396
rect 44548 44353 44557 44387
rect 44557 44353 44591 44387
rect 44591 44353 44600 44387
rect 44548 44344 44600 44353
rect 6828 44276 6880 44328
rect 9772 44319 9824 44328
rect 9772 44285 9781 44319
rect 9781 44285 9815 44319
rect 9815 44285 9824 44319
rect 9772 44276 9824 44285
rect 37280 44276 37332 44328
rect 44180 44276 44232 44328
rect 5632 44251 5684 44260
rect 5632 44217 5641 44251
rect 5641 44217 5675 44251
rect 5675 44217 5684 44251
rect 5632 44208 5684 44217
rect 41052 44208 41104 44260
rect 44364 44208 44416 44260
rect 45376 44208 45428 44260
rect 10048 44140 10100 44192
rect 10508 44140 10560 44192
rect 24860 44140 24912 44192
rect 37740 44140 37792 44192
rect 38752 44140 38804 44192
rect 40316 44140 40368 44192
rect 41972 44140 42024 44192
rect 43260 44183 43312 44192
rect 43260 44149 43269 44183
rect 43269 44149 43303 44183
rect 43303 44149 43312 44183
rect 43260 44140 43312 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 5908 43936 5960 43988
rect 9680 43936 9732 43988
rect 38476 43979 38528 43988
rect 38476 43945 38485 43979
rect 38485 43945 38519 43979
rect 38519 43945 38528 43979
rect 38476 43936 38528 43945
rect 41512 43936 41564 43988
rect 43996 43936 44048 43988
rect 45376 43979 45428 43988
rect 45376 43945 45385 43979
rect 45385 43945 45419 43979
rect 45419 43945 45428 43979
rect 45376 43936 45428 43945
rect 45560 43979 45612 43988
rect 45560 43945 45569 43979
rect 45569 43945 45603 43979
rect 45603 43945 45612 43979
rect 45560 43936 45612 43945
rect 9864 43800 9916 43852
rect 38660 43843 38712 43852
rect 38660 43809 38669 43843
rect 38669 43809 38703 43843
rect 38703 43809 38712 43843
rect 38660 43800 38712 43809
rect 41972 43843 42024 43852
rect 41972 43809 41981 43843
rect 41981 43809 42015 43843
rect 42015 43809 42024 43843
rect 41972 43800 42024 43809
rect 6276 43707 6328 43716
rect 6276 43673 6285 43707
rect 6285 43673 6319 43707
rect 6319 43673 6328 43707
rect 6276 43664 6328 43673
rect 6828 43664 6880 43716
rect 9128 43664 9180 43716
rect 9772 43732 9824 43784
rect 24584 43775 24636 43784
rect 24584 43741 24593 43775
rect 24593 43741 24627 43775
rect 24627 43741 24636 43775
rect 24584 43732 24636 43741
rect 24860 43775 24912 43784
rect 24860 43741 24894 43775
rect 24894 43741 24912 43775
rect 24860 43732 24912 43741
rect 10784 43664 10836 43716
rect 10968 43707 11020 43716
rect 10968 43673 10986 43707
rect 10986 43673 11020 43707
rect 10968 43664 11020 43673
rect 12348 43707 12400 43716
rect 12348 43673 12382 43707
rect 12382 43673 12400 43707
rect 37280 43732 37332 43784
rect 38752 43775 38804 43784
rect 38752 43741 38761 43775
rect 38761 43741 38795 43775
rect 38795 43741 38804 43775
rect 38752 43732 38804 43741
rect 40132 43732 40184 43784
rect 40316 43775 40368 43784
rect 40316 43741 40350 43775
rect 40350 43741 40368 43775
rect 40316 43732 40368 43741
rect 42156 43775 42208 43784
rect 42156 43741 42165 43775
rect 42165 43741 42199 43775
rect 42199 43741 42208 43775
rect 42156 43732 42208 43741
rect 43260 43775 43312 43784
rect 43260 43741 43269 43775
rect 43269 43741 43303 43775
rect 43303 43741 43312 43775
rect 43260 43732 43312 43741
rect 44272 43732 44324 43784
rect 45008 43732 45060 43784
rect 12348 43664 12400 43673
rect 7104 43596 7156 43648
rect 9864 43639 9916 43648
rect 9864 43605 9873 43639
rect 9873 43605 9907 43639
rect 9907 43605 9916 43639
rect 9864 43596 9916 43605
rect 13268 43596 13320 43648
rect 25504 43596 25556 43648
rect 40960 43596 41012 43648
rect 43168 43664 43220 43716
rect 43628 43664 43680 43716
rect 42340 43639 42392 43648
rect 42340 43605 42349 43639
rect 42349 43605 42383 43639
rect 42383 43605 42392 43639
rect 42340 43596 42392 43605
rect 44824 43596 44876 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 10968 43392 11020 43444
rect 38660 43392 38712 43444
rect 43628 43392 43680 43444
rect 5632 43367 5684 43376
rect 5632 43333 5641 43367
rect 5641 43333 5675 43367
rect 5675 43333 5684 43367
rect 5632 43324 5684 43333
rect 7012 43324 7064 43376
rect 7656 43324 7708 43376
rect 9128 43324 9180 43376
rect 37740 43367 37792 43376
rect 6276 43256 6328 43308
rect 7104 43299 7156 43308
rect 7104 43265 7113 43299
rect 7113 43265 7147 43299
rect 7147 43265 7156 43299
rect 7104 43256 7156 43265
rect 8760 43299 8812 43308
rect 8760 43265 8769 43299
rect 8769 43265 8803 43299
rect 8803 43265 8812 43299
rect 8760 43256 8812 43265
rect 10968 43299 11020 43308
rect 10968 43265 10977 43299
rect 10977 43265 11011 43299
rect 11011 43265 11020 43299
rect 10968 43256 11020 43265
rect 37740 43333 37774 43367
rect 37774 43333 37792 43367
rect 37740 43324 37792 43333
rect 40960 43367 41012 43376
rect 40960 43333 40969 43367
rect 40969 43333 41003 43367
rect 41003 43333 41012 43367
rect 40960 43324 41012 43333
rect 12348 43299 12400 43308
rect 12348 43265 12357 43299
rect 12357 43265 12391 43299
rect 12391 43265 12400 43299
rect 12348 43256 12400 43265
rect 42340 43324 42392 43376
rect 41328 43299 41380 43308
rect 41328 43265 41337 43299
rect 41337 43265 41371 43299
rect 41371 43265 41380 43299
rect 41328 43256 41380 43265
rect 44180 43392 44232 43444
rect 45192 43324 45244 43376
rect 37280 43188 37332 43240
rect 45008 43256 45060 43308
rect 43996 43188 44048 43240
rect 5908 43052 5960 43104
rect 42616 43120 42668 43172
rect 9772 43052 9824 43104
rect 44364 43052 44416 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 6276 42848 6328 42900
rect 6736 42848 6788 42900
rect 9128 42848 9180 42900
rect 44824 42848 44876 42900
rect 7656 42780 7708 42832
rect 6920 42644 6972 42696
rect 7104 42687 7156 42696
rect 7104 42653 7113 42687
rect 7113 42653 7147 42687
rect 7147 42653 7156 42687
rect 7288 42687 7340 42696
rect 7104 42644 7156 42653
rect 7288 42653 7297 42687
rect 7297 42653 7331 42687
rect 7331 42653 7340 42687
rect 7288 42644 7340 42653
rect 5724 42576 5776 42628
rect 7012 42576 7064 42628
rect 9772 42644 9824 42696
rect 24216 42644 24268 42696
rect 33876 42687 33928 42696
rect 33876 42653 33885 42687
rect 33885 42653 33919 42687
rect 33919 42653 33928 42687
rect 33876 42644 33928 42653
rect 35072 42687 35124 42696
rect 35072 42653 35081 42687
rect 35081 42653 35115 42687
rect 35115 42653 35124 42687
rect 35072 42644 35124 42653
rect 37372 42644 37424 42696
rect 43996 42644 44048 42696
rect 44180 42644 44232 42696
rect 44364 42644 44416 42696
rect 8300 42619 8352 42628
rect 8300 42585 8309 42619
rect 8309 42585 8343 42619
rect 8343 42585 8352 42619
rect 8300 42576 8352 42585
rect 9036 42576 9088 42628
rect 7196 42508 7248 42560
rect 7380 42508 7432 42560
rect 10508 42551 10560 42560
rect 10508 42517 10517 42551
rect 10517 42517 10551 42551
rect 10551 42517 10560 42551
rect 10508 42508 10560 42517
rect 38108 42551 38160 42560
rect 38108 42517 38117 42551
rect 38117 42517 38151 42551
rect 38151 42517 38160 42551
rect 38108 42508 38160 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 5724 42347 5776 42356
rect 5724 42313 5733 42347
rect 5733 42313 5767 42347
rect 5767 42313 5776 42347
rect 5724 42304 5776 42313
rect 9036 42347 9088 42356
rect 9036 42313 9045 42347
rect 9045 42313 9079 42347
rect 9079 42313 9088 42347
rect 9036 42304 9088 42313
rect 10968 42304 11020 42356
rect 5908 42211 5960 42220
rect 5908 42177 5917 42211
rect 5917 42177 5951 42211
rect 5951 42177 5960 42211
rect 5908 42168 5960 42177
rect 6736 42211 6788 42220
rect 6736 42177 6745 42211
rect 6745 42177 6779 42211
rect 6779 42177 6788 42211
rect 6736 42168 6788 42177
rect 7012 42211 7064 42220
rect 7012 42177 7021 42211
rect 7021 42177 7055 42211
rect 7055 42177 7064 42211
rect 7012 42168 7064 42177
rect 7104 42168 7156 42220
rect 8300 42168 8352 42220
rect 9128 42211 9180 42220
rect 9128 42177 9137 42211
rect 9137 42177 9171 42211
rect 9171 42177 9180 42211
rect 9128 42168 9180 42177
rect 10508 42236 10560 42288
rect 24216 42279 24268 42288
rect 9864 42143 9916 42152
rect 9864 42109 9873 42143
rect 9873 42109 9907 42143
rect 9907 42109 9916 42143
rect 9864 42100 9916 42109
rect 24216 42245 24250 42279
rect 24250 42245 24268 42279
rect 24216 42236 24268 42245
rect 24768 42168 24820 42220
rect 32404 42236 32456 42288
rect 38108 42236 38160 42288
rect 39212 42236 39264 42288
rect 44180 42236 44232 42288
rect 33876 42211 33928 42220
rect 33876 42177 33910 42211
rect 33910 42177 33928 42211
rect 33876 42168 33928 42177
rect 35072 42168 35124 42220
rect 43996 42168 44048 42220
rect 44364 42211 44416 42220
rect 44364 42177 44373 42211
rect 44373 42177 44407 42211
rect 44407 42177 44416 42211
rect 44364 42168 44416 42177
rect 23388 42100 23440 42152
rect 33324 42100 33376 42152
rect 37280 42100 37332 42152
rect 38568 42100 38620 42152
rect 29000 42032 29052 42084
rect 39304 42032 39356 42084
rect 44640 42032 44692 42084
rect 5908 41964 5960 42016
rect 12072 42007 12124 42016
rect 12072 41973 12081 42007
rect 12081 41973 12115 42007
rect 12115 41973 12124 42007
rect 12072 41964 12124 41973
rect 15292 42007 15344 42016
rect 15292 41973 15301 42007
rect 15301 41973 15335 42007
rect 15335 41973 15344 42007
rect 15292 41964 15344 41973
rect 23020 41964 23072 42016
rect 25596 41964 25648 42016
rect 34796 41964 34848 42016
rect 35348 41964 35400 42016
rect 40684 42007 40736 42016
rect 40684 41973 40693 42007
rect 40693 41973 40727 42007
rect 40727 41973 40736 42007
rect 40684 41964 40736 41973
rect 43444 42007 43496 42016
rect 43444 41973 43453 42007
rect 43453 41973 43487 42007
rect 43487 41973 43496 42007
rect 43444 41964 43496 41973
rect 45100 42007 45152 42016
rect 45100 41973 45109 42007
rect 45109 41973 45143 42007
rect 45143 41973 45152 42007
rect 45100 41964 45152 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 7104 41760 7156 41812
rect 7656 41803 7708 41812
rect 7656 41769 7665 41803
rect 7665 41769 7699 41803
rect 7699 41769 7708 41803
rect 7656 41760 7708 41769
rect 13268 41803 13320 41812
rect 13268 41769 13277 41803
rect 13277 41769 13311 41803
rect 13311 41769 13320 41803
rect 13268 41760 13320 41769
rect 27252 41803 27304 41812
rect 27252 41769 27261 41803
rect 27261 41769 27295 41803
rect 27295 41769 27304 41803
rect 27252 41760 27304 41769
rect 35348 41803 35400 41812
rect 35348 41769 35357 41803
rect 35357 41769 35391 41803
rect 35391 41769 35400 41803
rect 35348 41760 35400 41769
rect 41328 41760 41380 41812
rect 44640 41803 44692 41812
rect 44640 41769 44649 41803
rect 44649 41769 44683 41803
rect 44683 41769 44692 41803
rect 44640 41760 44692 41769
rect 7288 41624 7340 41676
rect 5264 41556 5316 41608
rect 5908 41599 5960 41608
rect 5908 41565 5942 41599
rect 5942 41565 5960 41599
rect 5908 41556 5960 41565
rect 7196 41556 7248 41608
rect 9128 41624 9180 41676
rect 9772 41624 9824 41676
rect 24584 41667 24636 41676
rect 24584 41633 24593 41667
rect 24593 41633 24627 41667
rect 24627 41633 24636 41667
rect 24584 41624 24636 41633
rect 9404 41556 9456 41608
rect 13176 41599 13228 41608
rect 13176 41565 13185 41599
rect 13185 41565 13219 41599
rect 13219 41565 13228 41599
rect 13176 41556 13228 41565
rect 13268 41599 13320 41608
rect 13268 41565 13277 41599
rect 13277 41565 13311 41599
rect 13311 41565 13320 41599
rect 14924 41599 14976 41608
rect 13268 41556 13320 41565
rect 14924 41565 14933 41599
rect 14933 41565 14967 41599
rect 14967 41565 14976 41599
rect 14924 41556 14976 41565
rect 22100 41556 22152 41608
rect 11152 41488 11204 41540
rect 12440 41420 12492 41472
rect 21088 41488 21140 41540
rect 25228 41556 25280 41608
rect 29000 41624 29052 41676
rect 27068 41599 27120 41608
rect 27068 41565 27077 41599
rect 27077 41565 27111 41599
rect 27111 41565 27120 41599
rect 27068 41556 27120 41565
rect 27436 41556 27488 41608
rect 38568 41692 38620 41744
rect 34796 41624 34848 41676
rect 38660 41624 38712 41676
rect 37188 41556 37240 41608
rect 37372 41599 37424 41608
rect 37372 41565 37406 41599
rect 37406 41565 37424 41599
rect 37372 41556 37424 41565
rect 39304 41599 39356 41608
rect 39304 41565 39313 41599
rect 39313 41565 39347 41599
rect 39347 41565 39356 41599
rect 39304 41556 39356 41565
rect 40684 41599 40736 41608
rect 40684 41565 40718 41599
rect 40718 41565 40736 41599
rect 40684 41556 40736 41565
rect 27344 41531 27396 41540
rect 27344 41497 27353 41531
rect 27353 41497 27387 41531
rect 27387 41497 27396 41531
rect 27344 41488 27396 41497
rect 13452 41463 13504 41472
rect 13452 41429 13461 41463
rect 13461 41429 13495 41463
rect 13495 41429 13504 41463
rect 13452 41420 13504 41429
rect 16764 41420 16816 41472
rect 22744 41420 22796 41472
rect 25780 41420 25832 41472
rect 33324 41488 33376 41540
rect 35072 41531 35124 41540
rect 35072 41497 35081 41531
rect 35081 41497 35115 41531
rect 35115 41497 35124 41531
rect 35072 41488 35124 41497
rect 39120 41488 39172 41540
rect 34980 41420 35032 41472
rect 38752 41420 38804 41472
rect 42156 41420 42208 41472
rect 43444 41488 43496 41540
rect 45008 41420 45060 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 13268 41216 13320 41268
rect 22100 41216 22152 41268
rect 23388 41216 23440 41268
rect 22744 41191 22796 41200
rect 22744 41157 22753 41191
rect 22753 41157 22787 41191
rect 22787 41157 22796 41191
rect 22744 41148 22796 41157
rect 9128 41123 9180 41132
rect 9128 41089 9137 41123
rect 9137 41089 9171 41123
rect 9171 41089 9180 41123
rect 9128 41080 9180 41089
rect 8576 41012 8628 41064
rect 11152 41123 11204 41132
rect 11152 41089 11161 41123
rect 11161 41089 11195 41123
rect 11195 41089 11204 41123
rect 11152 41080 11204 41089
rect 15200 41123 15252 41132
rect 15200 41089 15234 41123
rect 15234 41089 15252 41123
rect 21088 41123 21140 41132
rect 15200 41080 15252 41089
rect 21088 41089 21097 41123
rect 21097 41089 21131 41123
rect 21131 41089 21140 41123
rect 21088 41080 21140 41089
rect 27344 41216 27396 41268
rect 27988 41216 28040 41268
rect 35072 41216 35124 41268
rect 44180 41216 44232 41268
rect 45100 41148 45152 41200
rect 13820 41012 13872 41064
rect 14924 41055 14976 41064
rect 14924 41021 14933 41055
rect 14933 41021 14967 41055
rect 14967 41021 14976 41055
rect 14924 41012 14976 41021
rect 22928 41055 22980 41064
rect 22928 41021 22937 41055
rect 22937 41021 22971 41055
rect 22971 41021 22980 41055
rect 22928 41012 22980 41021
rect 24492 41080 24544 41132
rect 25780 41123 25832 41132
rect 25780 41089 25789 41123
rect 25789 41089 25823 41123
rect 25823 41089 25832 41123
rect 25780 41080 25832 41089
rect 28264 41080 28316 41132
rect 29000 41080 29052 41132
rect 30380 41080 30432 41132
rect 33324 41080 33376 41132
rect 33508 41123 33560 41132
rect 33508 41089 33542 41123
rect 33542 41089 33560 41123
rect 33508 41080 33560 41089
rect 34980 41080 35032 41132
rect 37740 41123 37792 41132
rect 37740 41089 37774 41123
rect 37774 41089 37792 41123
rect 37740 41080 37792 41089
rect 41328 41080 41380 41132
rect 45008 41123 45060 41132
rect 45008 41089 45017 41123
rect 45017 41089 45051 41123
rect 45051 41089 45060 41123
rect 45008 41080 45060 41089
rect 23572 41012 23624 41064
rect 25596 41055 25648 41064
rect 25596 41021 25605 41055
rect 25605 41021 25639 41055
rect 25639 41021 25648 41055
rect 25596 41012 25648 41021
rect 37280 41012 37332 41064
rect 40316 41012 40368 41064
rect 5540 40919 5592 40928
rect 5540 40885 5549 40919
rect 5549 40885 5583 40919
rect 5583 40885 5592 40919
rect 5540 40876 5592 40885
rect 11152 40876 11204 40928
rect 16856 40876 16908 40928
rect 22284 40876 22336 40928
rect 23020 40919 23072 40928
rect 23020 40885 23029 40919
rect 23029 40885 23063 40919
rect 23063 40885 23072 40919
rect 23020 40876 23072 40885
rect 23204 40919 23256 40928
rect 23204 40885 23213 40919
rect 23213 40885 23247 40919
rect 23247 40885 23256 40919
rect 23204 40876 23256 40885
rect 25504 40919 25556 40928
rect 25504 40885 25513 40919
rect 25513 40885 25547 40919
rect 25547 40885 25556 40919
rect 25504 40876 25556 40885
rect 25688 40876 25740 40928
rect 30104 40919 30156 40928
rect 30104 40885 30113 40919
rect 30113 40885 30147 40919
rect 30147 40885 30156 40919
rect 30104 40876 30156 40885
rect 39028 40876 39080 40928
rect 40132 40919 40184 40928
rect 40132 40885 40141 40919
rect 40141 40885 40175 40919
rect 40175 40885 40184 40919
rect 40132 40876 40184 40885
rect 42432 40876 42484 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 8576 40715 8628 40724
rect 8576 40681 8585 40715
rect 8585 40681 8619 40715
rect 8619 40681 8628 40715
rect 8576 40672 8628 40681
rect 13176 40715 13228 40724
rect 13176 40681 13185 40715
rect 13185 40681 13219 40715
rect 13219 40681 13228 40715
rect 13176 40672 13228 40681
rect 16764 40715 16816 40724
rect 16764 40681 16773 40715
rect 16773 40681 16807 40715
rect 16807 40681 16816 40715
rect 16764 40672 16816 40681
rect 24492 40672 24544 40724
rect 26332 40715 26384 40724
rect 26332 40681 26341 40715
rect 26341 40681 26375 40715
rect 26375 40681 26384 40715
rect 26332 40672 26384 40681
rect 27068 40672 27120 40724
rect 33508 40715 33560 40724
rect 5264 40579 5316 40588
rect 5264 40545 5273 40579
rect 5273 40545 5307 40579
rect 5307 40545 5316 40579
rect 5264 40536 5316 40545
rect 9128 40579 9180 40588
rect 9128 40545 9137 40579
rect 9137 40545 9171 40579
rect 9171 40545 9180 40579
rect 9128 40536 9180 40545
rect 13820 40536 13872 40588
rect 14924 40579 14976 40588
rect 14924 40545 14933 40579
rect 14933 40545 14967 40579
rect 14967 40545 14976 40579
rect 14924 40536 14976 40545
rect 5540 40511 5592 40520
rect 5540 40477 5574 40511
rect 5574 40477 5592 40511
rect 5540 40468 5592 40477
rect 9404 40511 9456 40520
rect 9404 40477 9438 40511
rect 9438 40477 9456 40511
rect 9404 40468 9456 40477
rect 11796 40511 11848 40520
rect 11796 40477 11805 40511
rect 11805 40477 11839 40511
rect 11839 40477 11848 40511
rect 11796 40468 11848 40477
rect 12072 40511 12124 40520
rect 12072 40477 12106 40511
rect 12106 40477 12124 40511
rect 12072 40468 12124 40477
rect 16856 40579 16908 40588
rect 16856 40545 16865 40579
rect 16865 40545 16899 40579
rect 16899 40545 16908 40579
rect 16856 40536 16908 40545
rect 22100 40536 22152 40588
rect 33508 40681 33517 40715
rect 33517 40681 33551 40715
rect 33551 40681 33560 40715
rect 33508 40672 33560 40681
rect 38752 40715 38804 40724
rect 38752 40681 38761 40715
rect 38761 40681 38795 40715
rect 38795 40681 38804 40715
rect 38752 40672 38804 40681
rect 39120 40672 39172 40724
rect 42156 40715 42208 40724
rect 42156 40681 42165 40715
rect 42165 40681 42199 40715
rect 42199 40681 42208 40715
rect 42156 40672 42208 40681
rect 42616 40715 42668 40724
rect 42616 40681 42625 40715
rect 42625 40681 42659 40715
rect 42659 40681 42668 40715
rect 42616 40672 42668 40681
rect 22468 40468 22520 40520
rect 23204 40468 23256 40520
rect 25688 40511 25740 40520
rect 25688 40477 25697 40511
rect 25697 40477 25731 40511
rect 25731 40477 25740 40511
rect 25688 40468 25740 40477
rect 27436 40511 27488 40520
rect 13820 40400 13872 40452
rect 16764 40443 16816 40452
rect 16764 40409 16773 40443
rect 16773 40409 16807 40443
rect 16807 40409 16816 40443
rect 16764 40400 16816 40409
rect 24216 40400 24268 40452
rect 24768 40400 24820 40452
rect 27436 40477 27445 40511
rect 27445 40477 27479 40511
rect 27479 40477 27488 40511
rect 27436 40468 27488 40477
rect 27528 40400 27580 40452
rect 27988 40511 28040 40520
rect 27988 40477 27997 40511
rect 27997 40477 28031 40511
rect 28031 40477 28040 40511
rect 27988 40468 28040 40477
rect 29736 40468 29788 40520
rect 30104 40511 30156 40520
rect 30104 40477 30138 40511
rect 30138 40477 30156 40511
rect 30104 40468 30156 40477
rect 39028 40511 39080 40520
rect 39028 40477 39037 40511
rect 39037 40477 39071 40511
rect 39071 40477 39080 40511
rect 39028 40468 39080 40477
rect 40316 40511 40368 40520
rect 40316 40477 40325 40511
rect 40325 40477 40359 40511
rect 40359 40477 40368 40511
rect 40316 40468 40368 40477
rect 41788 40468 41840 40520
rect 42432 40511 42484 40520
rect 42432 40477 42441 40511
rect 42441 40477 42475 40511
rect 42475 40477 42484 40511
rect 42432 40468 42484 40477
rect 37280 40400 37332 40452
rect 38844 40400 38896 40452
rect 40592 40443 40644 40452
rect 40592 40409 40626 40443
rect 40626 40409 40644 40443
rect 40592 40400 40644 40409
rect 6920 40332 6972 40384
rect 11244 40332 11296 40384
rect 17224 40375 17276 40384
rect 17224 40341 17233 40375
rect 17233 40341 17267 40375
rect 17267 40341 17276 40375
rect 17224 40332 17276 40341
rect 26700 40375 26752 40384
rect 26700 40341 26709 40375
rect 26709 40341 26743 40375
rect 26743 40341 26752 40375
rect 26700 40332 26752 40341
rect 28448 40332 28500 40384
rect 31208 40375 31260 40384
rect 31208 40341 31217 40375
rect 31217 40341 31251 40375
rect 31251 40341 31260 40375
rect 31208 40332 31260 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 7196 40171 7248 40180
rect 7196 40137 7205 40171
rect 7205 40137 7239 40171
rect 7239 40137 7248 40171
rect 7196 40128 7248 40137
rect 12440 40128 12492 40180
rect 7656 39992 7708 40044
rect 8760 40035 8812 40044
rect 8760 40001 8769 40035
rect 8769 40001 8803 40035
rect 8803 40001 8812 40035
rect 8760 39992 8812 40001
rect 6644 39924 6696 39976
rect 13820 40103 13872 40112
rect 13820 40069 13829 40103
rect 13829 40069 13863 40103
rect 13863 40069 13872 40103
rect 13820 40060 13872 40069
rect 22928 40128 22980 40180
rect 28264 40171 28316 40180
rect 17224 40060 17276 40112
rect 26700 40060 26752 40112
rect 13176 40035 13228 40044
rect 13176 40001 13185 40035
rect 13185 40001 13219 40035
rect 13219 40001 13228 40035
rect 13176 39992 13228 40001
rect 13544 39924 13596 39976
rect 11060 39899 11112 39908
rect 11060 39865 11069 39899
rect 11069 39865 11103 39899
rect 11103 39865 11112 39899
rect 22100 39992 22152 40044
rect 22284 40035 22336 40044
rect 22284 40001 22318 40035
rect 22318 40001 22336 40035
rect 22284 39992 22336 40001
rect 25228 40035 25280 40044
rect 25228 40001 25237 40035
rect 25237 40001 25271 40035
rect 25271 40001 25280 40035
rect 25228 39992 25280 40001
rect 27620 40035 27672 40044
rect 27620 40001 27629 40035
rect 27629 40001 27663 40035
rect 27663 40001 27672 40035
rect 27620 39992 27672 40001
rect 27712 39992 27764 40044
rect 28264 40137 28273 40171
rect 28273 40137 28307 40171
rect 28307 40137 28316 40171
rect 28264 40128 28316 40137
rect 30380 40171 30432 40180
rect 30380 40137 30389 40171
rect 30389 40137 30423 40171
rect 30423 40137 30432 40171
rect 30380 40128 30432 40137
rect 38844 40171 38896 40180
rect 38844 40137 38853 40171
rect 38853 40137 38887 40171
rect 38887 40137 38896 40171
rect 38844 40128 38896 40137
rect 41788 40171 41840 40180
rect 41788 40137 41797 40171
rect 41797 40137 41831 40171
rect 41831 40137 41840 40171
rect 41788 40128 41840 40137
rect 40132 40060 40184 40112
rect 28448 40035 28500 40044
rect 28448 40001 28457 40035
rect 28457 40001 28491 40035
rect 28491 40001 28500 40035
rect 28448 39992 28500 40001
rect 27988 39924 28040 39976
rect 11060 39856 11112 39865
rect 27528 39856 27580 39908
rect 30564 39992 30616 40044
rect 31208 39992 31260 40044
rect 37280 39924 37332 39976
rect 40316 39924 40368 39976
rect 5540 39788 5592 39840
rect 6920 39831 6972 39840
rect 6920 39797 6929 39831
rect 6929 39797 6963 39831
rect 6963 39797 6972 39831
rect 6920 39788 6972 39797
rect 9220 39788 9272 39840
rect 13452 39788 13504 39840
rect 24216 39831 24268 39840
rect 24216 39797 24225 39831
rect 24225 39797 24259 39831
rect 24259 39797 24268 39831
rect 24216 39788 24268 39797
rect 40684 39788 40736 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 6644 39627 6696 39636
rect 6644 39593 6653 39627
rect 6653 39593 6687 39627
rect 6687 39593 6696 39627
rect 6644 39584 6696 39593
rect 7288 39627 7340 39636
rect 7288 39593 7297 39627
rect 7297 39593 7331 39627
rect 7331 39593 7340 39627
rect 7288 39584 7340 39593
rect 7656 39627 7708 39636
rect 7656 39593 7665 39627
rect 7665 39593 7699 39627
rect 7699 39593 7708 39627
rect 7656 39584 7708 39593
rect 11152 39627 11204 39636
rect 11152 39593 11161 39627
rect 11161 39593 11195 39627
rect 11195 39593 11204 39627
rect 11152 39584 11204 39593
rect 13176 39584 13228 39636
rect 15200 39584 15252 39636
rect 16764 39584 16816 39636
rect 23572 39627 23624 39636
rect 23572 39593 23581 39627
rect 23581 39593 23615 39627
rect 23615 39593 23624 39627
rect 23572 39584 23624 39593
rect 37740 39584 37792 39636
rect 40592 39584 40644 39636
rect 41328 39627 41380 39636
rect 41328 39593 41337 39627
rect 41337 39593 41371 39627
rect 41371 39593 41380 39627
rect 41328 39584 41380 39593
rect 5264 39491 5316 39500
rect 5264 39457 5273 39491
rect 5273 39457 5307 39491
rect 5307 39457 5316 39491
rect 5264 39448 5316 39457
rect 7380 39491 7432 39500
rect 7380 39457 7389 39491
rect 7389 39457 7423 39491
rect 7423 39457 7432 39491
rect 7380 39448 7432 39457
rect 14924 39448 14976 39500
rect 22100 39448 22152 39500
rect 5540 39423 5592 39432
rect 5540 39389 5574 39423
rect 5574 39389 5592 39423
rect 5540 39380 5592 39389
rect 7472 39423 7524 39432
rect 7472 39389 7481 39423
rect 7481 39389 7515 39423
rect 7515 39389 7524 39423
rect 7472 39380 7524 39389
rect 8392 39380 8444 39432
rect 8760 39380 8812 39432
rect 9220 39380 9272 39432
rect 7196 39355 7248 39364
rect 7196 39321 7205 39355
rect 7205 39321 7239 39355
rect 7239 39321 7248 39355
rect 7196 39312 7248 39321
rect 11244 39380 11296 39432
rect 15292 39423 15344 39432
rect 15292 39389 15326 39423
rect 15326 39389 15344 39423
rect 15292 39380 15344 39389
rect 22468 39423 22520 39432
rect 22468 39389 22502 39423
rect 22502 39389 22520 39423
rect 22468 39380 22520 39389
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 11060 39040 11112 39092
rect 27528 39040 27580 39092
rect 22100 38904 22152 38956
rect 23296 38904 23348 38956
rect 23480 38947 23532 38956
rect 23480 38913 23514 38947
rect 23514 38913 23532 38947
rect 23480 38904 23532 38913
rect 27712 39015 27764 39024
rect 27712 38981 27721 39015
rect 27721 38981 27755 39015
rect 27755 38981 27764 39015
rect 27712 38972 27764 38981
rect 27436 38947 27488 38956
rect 27436 38913 27445 38947
rect 27445 38913 27479 38947
rect 27479 38913 27488 38947
rect 27436 38904 27488 38913
rect 28172 38904 28224 38956
rect 30564 38947 30616 38956
rect 30564 38913 30573 38947
rect 30573 38913 30607 38947
rect 30607 38913 30616 38947
rect 30564 38904 30616 38913
rect 30840 38904 30892 38956
rect 40776 38947 40828 38956
rect 40776 38913 40785 38947
rect 40785 38913 40819 38947
rect 40819 38913 40828 38947
rect 40776 38904 40828 38913
rect 41604 38904 41656 38956
rect 28356 38836 28408 38888
rect 5264 38768 5316 38820
rect 6920 38768 6972 38820
rect 5540 38700 5592 38752
rect 7012 38700 7064 38752
rect 8760 38743 8812 38752
rect 8760 38709 8769 38743
rect 8769 38709 8803 38743
rect 8803 38709 8812 38743
rect 8760 38700 8812 38709
rect 11704 38743 11756 38752
rect 11704 38709 11713 38743
rect 11713 38709 11747 38743
rect 11747 38709 11756 38743
rect 11704 38700 11756 38709
rect 24584 38743 24636 38752
rect 24584 38709 24593 38743
rect 24593 38709 24627 38743
rect 24627 38709 24636 38743
rect 24584 38700 24636 38709
rect 30748 38700 30800 38752
rect 36636 38700 36688 38752
rect 41972 38700 42024 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 7472 38496 7524 38548
rect 13544 38539 13596 38548
rect 13544 38505 13553 38539
rect 13553 38505 13587 38539
rect 13587 38505 13596 38539
rect 13544 38496 13596 38505
rect 23480 38496 23532 38548
rect 27712 38496 27764 38548
rect 28448 38496 28500 38548
rect 7288 38428 7340 38480
rect 5264 38403 5316 38412
rect 5264 38369 5273 38403
rect 5273 38369 5307 38403
rect 5307 38369 5316 38403
rect 5264 38360 5316 38369
rect 13176 38403 13228 38412
rect 13176 38369 13185 38403
rect 13185 38369 13219 38403
rect 13219 38369 13228 38403
rect 13176 38360 13228 38369
rect 5540 38335 5592 38344
rect 5540 38301 5574 38335
rect 5574 38301 5592 38335
rect 5540 38292 5592 38301
rect 8392 38292 8444 38344
rect 8760 38292 8812 38344
rect 9772 38292 9824 38344
rect 10600 38335 10652 38344
rect 10600 38301 10609 38335
rect 10609 38301 10643 38335
rect 10643 38301 10652 38335
rect 10600 38292 10652 38301
rect 11796 38292 11848 38344
rect 12532 38292 12584 38344
rect 13912 38292 13964 38344
rect 23572 38335 23624 38344
rect 23572 38301 23581 38335
rect 23581 38301 23615 38335
rect 23615 38301 23624 38335
rect 23572 38292 23624 38301
rect 27620 38428 27672 38480
rect 28908 38496 28960 38548
rect 39212 38539 39264 38548
rect 39212 38505 39221 38539
rect 39221 38505 39255 38539
rect 39255 38505 39264 38539
rect 39212 38496 39264 38505
rect 42800 38496 42852 38548
rect 44456 38496 44508 38548
rect 31760 38428 31812 38480
rect 27436 38292 27488 38344
rect 28356 38292 28408 38344
rect 11704 38224 11756 38276
rect 13084 38267 13136 38276
rect 13084 38233 13093 38267
rect 13093 38233 13127 38267
rect 13127 38233 13136 38267
rect 13084 38224 13136 38233
rect 29644 38224 29696 38276
rect 30748 38267 30800 38276
rect 30748 38233 30757 38267
rect 30757 38233 30791 38267
rect 30791 38233 30800 38267
rect 30748 38224 30800 38233
rect 26240 38199 26292 38208
rect 26240 38165 26249 38199
rect 26249 38165 26283 38199
rect 26283 38165 26292 38199
rect 26240 38156 26292 38165
rect 28172 38156 28224 38208
rect 28356 38156 28408 38208
rect 30012 38199 30064 38208
rect 30012 38165 30037 38199
rect 30037 38165 30064 38199
rect 30012 38156 30064 38165
rect 30932 38199 30984 38208
rect 37280 38292 37332 38344
rect 40132 38292 40184 38344
rect 40684 38335 40736 38344
rect 40684 38301 40693 38335
rect 40693 38301 40727 38335
rect 40727 38301 40736 38335
rect 40684 38292 40736 38301
rect 42064 38292 42116 38344
rect 42708 38224 42760 38276
rect 30932 38165 30957 38199
rect 30957 38165 30984 38199
rect 30932 38156 30984 38165
rect 31852 38199 31904 38208
rect 31852 38165 31861 38199
rect 31861 38165 31895 38199
rect 31895 38165 31904 38199
rect 31852 38156 31904 38165
rect 38292 38156 38344 38208
rect 40316 38156 40368 38208
rect 41604 38156 41656 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 6920 37952 6972 38004
rect 7380 37952 7432 38004
rect 13084 37952 13136 38004
rect 13912 37995 13964 38004
rect 13912 37961 13921 37995
rect 13921 37961 13955 37995
rect 13955 37961 13964 37995
rect 13912 37952 13964 37961
rect 8760 37884 8812 37936
rect 10600 37884 10652 37936
rect 7012 37859 7064 37868
rect 7012 37825 7046 37859
rect 7046 37825 7064 37859
rect 23572 37927 23624 37936
rect 23572 37893 23606 37927
rect 23606 37893 23624 37927
rect 23572 37884 23624 37893
rect 27528 37927 27580 37936
rect 27528 37893 27537 37927
rect 27537 37893 27571 37927
rect 27571 37893 27580 37927
rect 27528 37884 27580 37893
rect 30564 37952 30616 38004
rect 30932 37952 30984 38004
rect 42064 37995 42116 38004
rect 42064 37961 42073 37995
rect 42073 37961 42107 37995
rect 42107 37961 42116 37995
rect 42064 37952 42116 37961
rect 7012 37816 7064 37825
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 23296 37859 23348 37868
rect 23296 37825 23305 37859
rect 23305 37825 23339 37859
rect 23339 37825 23348 37859
rect 23296 37816 23348 37825
rect 28172 37859 28224 37868
rect 28172 37825 28181 37859
rect 28181 37825 28215 37859
rect 28215 37825 28224 37859
rect 28172 37816 28224 37825
rect 28356 37859 28408 37868
rect 28356 37825 28365 37859
rect 28365 37825 28399 37859
rect 28399 37825 28408 37859
rect 28356 37816 28408 37825
rect 30840 37884 30892 37936
rect 30380 37859 30432 37868
rect 9772 37791 9824 37800
rect 9772 37757 9781 37791
rect 9781 37757 9815 37791
rect 9815 37757 9824 37791
rect 9772 37748 9824 37757
rect 30380 37825 30389 37859
rect 30389 37825 30423 37859
rect 30423 37825 30432 37859
rect 30380 37816 30432 37825
rect 31116 37816 31168 37868
rect 31484 37859 31536 37868
rect 31484 37825 31493 37859
rect 31493 37825 31527 37859
rect 31527 37825 31536 37859
rect 31484 37816 31536 37825
rect 28356 37680 28408 37732
rect 30288 37680 30340 37732
rect 5816 37655 5868 37664
rect 5816 37621 5825 37655
rect 5825 37621 5859 37655
rect 5859 37621 5868 37655
rect 5816 37612 5868 37621
rect 24676 37655 24728 37664
rect 24676 37621 24685 37655
rect 24685 37621 24719 37655
rect 24719 37621 24728 37655
rect 24676 37612 24728 37621
rect 27068 37612 27120 37664
rect 27712 37612 27764 37664
rect 28816 37612 28868 37664
rect 29644 37655 29696 37664
rect 29644 37621 29653 37655
rect 29653 37621 29687 37655
rect 29687 37621 29696 37655
rect 29644 37612 29696 37621
rect 31852 37884 31904 37936
rect 39212 37884 39264 37936
rect 39396 37927 39448 37936
rect 39396 37893 39405 37927
rect 39405 37893 39439 37927
rect 39439 37893 39448 37927
rect 39396 37884 39448 37893
rect 42800 37927 42852 37936
rect 42800 37893 42809 37927
rect 42809 37893 42843 37927
rect 42843 37893 42852 37927
rect 42800 37884 42852 37893
rect 44548 37927 44600 37936
rect 44548 37893 44557 37927
rect 44557 37893 44591 37927
rect 44591 37893 44600 37927
rect 44548 37884 44600 37893
rect 36636 37859 36688 37868
rect 36636 37825 36654 37859
rect 36654 37825 36688 37859
rect 36636 37816 36688 37825
rect 37280 37816 37332 37868
rect 37740 37859 37792 37868
rect 37740 37825 37774 37859
rect 37774 37825 37792 37859
rect 37740 37816 37792 37825
rect 32312 37791 32364 37800
rect 32312 37757 32321 37791
rect 32321 37757 32355 37791
rect 32355 37757 32364 37791
rect 32312 37748 32364 37757
rect 37464 37791 37516 37800
rect 37464 37757 37473 37791
rect 37473 37757 37507 37791
rect 37507 37757 37516 37791
rect 37464 37748 37516 37757
rect 41604 37791 41656 37800
rect 41604 37757 41613 37791
rect 41613 37757 41647 37791
rect 41647 37757 41656 37791
rect 41604 37748 41656 37757
rect 41880 37723 41932 37732
rect 41880 37689 41889 37723
rect 41889 37689 41923 37723
rect 41923 37689 41932 37723
rect 41880 37680 41932 37689
rect 31852 37612 31904 37664
rect 38200 37612 38252 37664
rect 38844 37655 38896 37664
rect 38844 37621 38853 37655
rect 38853 37621 38887 37655
rect 38887 37621 38896 37655
rect 38844 37612 38896 37621
rect 40040 37612 40092 37664
rect 40684 37655 40736 37664
rect 40684 37621 40693 37655
rect 40693 37621 40727 37655
rect 40727 37621 40736 37655
rect 40684 37612 40736 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 13176 37408 13228 37460
rect 24584 37451 24636 37460
rect 24584 37417 24593 37451
rect 24593 37417 24627 37451
rect 24627 37417 24636 37451
rect 24584 37408 24636 37417
rect 27436 37451 27488 37460
rect 27436 37417 27445 37451
rect 27445 37417 27479 37451
rect 27479 37417 27488 37451
rect 27436 37408 27488 37417
rect 28356 37408 28408 37460
rect 28816 37451 28868 37460
rect 28816 37417 28825 37451
rect 28825 37417 28859 37451
rect 28859 37417 28868 37451
rect 28816 37408 28868 37417
rect 30656 37408 30708 37460
rect 31116 37451 31168 37460
rect 31116 37417 31125 37451
rect 31125 37417 31159 37451
rect 31159 37417 31168 37451
rect 38200 37451 38252 37460
rect 31116 37408 31168 37417
rect 5264 37272 5316 37324
rect 24676 37315 24728 37324
rect 24676 37281 24685 37315
rect 24685 37281 24719 37315
rect 24719 37281 24728 37315
rect 24676 37272 24728 37281
rect 5816 37247 5868 37256
rect 5816 37213 5850 37247
rect 5850 37213 5868 37247
rect 5816 37204 5868 37213
rect 9772 37204 9824 37256
rect 23296 37204 23348 37256
rect 24860 37247 24912 37256
rect 24860 37213 24869 37247
rect 24869 37213 24903 37247
rect 24903 37213 24912 37247
rect 24860 37204 24912 37213
rect 31484 37340 31536 37392
rect 29736 37247 29788 37256
rect 11888 37179 11940 37188
rect 11888 37145 11922 37179
rect 11922 37145 11940 37179
rect 11888 37136 11940 37145
rect 22928 37179 22980 37188
rect 22928 37145 22962 37179
rect 22962 37145 22980 37179
rect 22928 37136 22980 37145
rect 7196 37068 7248 37120
rect 25596 37068 25648 37120
rect 26240 37136 26292 37188
rect 27804 37136 27856 37188
rect 28632 37136 28684 37188
rect 27160 37068 27212 37120
rect 28908 37136 28960 37188
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 30288 37204 30340 37256
rect 31852 37315 31904 37324
rect 31852 37281 31861 37315
rect 31861 37281 31895 37315
rect 31895 37281 31904 37315
rect 31852 37272 31904 37281
rect 38200 37417 38209 37451
rect 38209 37417 38243 37451
rect 38243 37417 38252 37451
rect 38200 37408 38252 37417
rect 40224 37408 40276 37460
rect 42708 37451 42760 37460
rect 42708 37417 42717 37451
rect 42717 37417 42751 37451
rect 42751 37417 42760 37451
rect 42708 37408 42760 37417
rect 38292 37315 38344 37324
rect 38292 37281 38301 37315
rect 38301 37281 38335 37315
rect 38335 37281 38344 37315
rect 38292 37272 38344 37281
rect 40040 37315 40092 37324
rect 36176 37204 36228 37256
rect 37464 37204 37516 37256
rect 40040 37281 40049 37315
rect 40049 37281 40083 37315
rect 40083 37281 40092 37315
rect 40040 37272 40092 37281
rect 38844 37204 38896 37256
rect 39304 37247 39356 37256
rect 39304 37213 39313 37247
rect 39313 37213 39347 37247
rect 39347 37213 39356 37247
rect 39304 37204 39356 37213
rect 40316 37247 40368 37256
rect 40316 37213 40350 37247
rect 40350 37213 40368 37247
rect 36636 37179 36688 37188
rect 36636 37145 36670 37179
rect 36670 37145 36688 37179
rect 36636 37136 36688 37145
rect 40316 37204 40368 37213
rect 41604 37136 41656 37188
rect 41880 37179 41932 37188
rect 41880 37145 41889 37179
rect 41889 37145 41923 37179
rect 41923 37145 41932 37179
rect 41880 37136 41932 37145
rect 41972 37136 42024 37188
rect 38660 37111 38712 37120
rect 38660 37077 38669 37111
rect 38669 37077 38703 37111
rect 38703 37077 38712 37111
rect 38660 37068 38712 37077
rect 41420 37111 41472 37120
rect 41420 37077 41429 37111
rect 41429 37077 41463 37111
rect 41463 37077 41472 37111
rect 41420 37068 41472 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 24860 36907 24912 36916
rect 24860 36873 24869 36907
rect 24869 36873 24903 36907
rect 24903 36873 24912 36907
rect 24860 36864 24912 36873
rect 27528 36864 27580 36916
rect 11888 36771 11940 36780
rect 11888 36737 11897 36771
rect 11897 36737 11931 36771
rect 11931 36737 11940 36771
rect 11888 36728 11940 36737
rect 22928 36728 22980 36780
rect 23756 36771 23808 36780
rect 23756 36737 23790 36771
rect 23790 36737 23808 36771
rect 28172 36796 28224 36848
rect 29736 36864 29788 36916
rect 31116 36864 31168 36916
rect 32312 36864 32364 36916
rect 32404 36907 32456 36916
rect 32404 36873 32413 36907
rect 32413 36873 32447 36907
rect 32447 36873 32456 36907
rect 40132 36907 40184 36916
rect 32404 36864 32456 36873
rect 40132 36873 40141 36907
rect 40141 36873 40175 36907
rect 40175 36873 40184 36907
rect 40132 36864 40184 36873
rect 40316 36907 40368 36916
rect 40316 36873 40325 36907
rect 40325 36873 40359 36907
rect 40359 36873 40368 36907
rect 40316 36864 40368 36873
rect 41880 36864 41932 36916
rect 23756 36728 23808 36737
rect 27160 36771 27212 36780
rect 23480 36703 23532 36712
rect 23480 36669 23489 36703
rect 23489 36669 23523 36703
rect 23523 36669 23532 36703
rect 23480 36660 23532 36669
rect 27160 36737 27169 36771
rect 27169 36737 27203 36771
rect 27203 36737 27212 36771
rect 27160 36728 27212 36737
rect 27252 36728 27304 36780
rect 36636 36771 36688 36780
rect 36636 36737 36645 36771
rect 36645 36737 36679 36771
rect 36679 36737 36688 36771
rect 36636 36728 36688 36737
rect 37740 36728 37792 36780
rect 39488 36771 39540 36780
rect 39488 36737 39497 36771
rect 39497 36737 39531 36771
rect 39531 36737 39540 36771
rect 39488 36728 39540 36737
rect 41420 36728 41472 36780
rect 39304 36635 39356 36644
rect 39304 36601 39313 36635
rect 39313 36601 39347 36635
rect 39347 36601 39356 36635
rect 39304 36592 39356 36601
rect 40776 36592 40828 36644
rect 28356 36524 28408 36576
rect 33232 36524 33284 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 23756 36363 23808 36372
rect 23756 36329 23765 36363
rect 23765 36329 23799 36363
rect 23799 36329 23808 36363
rect 23756 36320 23808 36329
rect 27252 36363 27304 36372
rect 27252 36329 27261 36363
rect 27261 36329 27295 36363
rect 27295 36329 27304 36363
rect 27252 36320 27304 36329
rect 30196 36320 30248 36372
rect 40316 36363 40368 36372
rect 40316 36329 40325 36363
rect 40325 36329 40359 36363
rect 40359 36329 40368 36363
rect 40316 36320 40368 36329
rect 31116 36227 31168 36236
rect 31116 36193 31125 36227
rect 31125 36193 31159 36227
rect 31159 36193 31168 36227
rect 31116 36184 31168 36193
rect 32312 36184 32364 36236
rect 32956 36227 33008 36236
rect 32956 36193 32965 36227
rect 32965 36193 32999 36227
rect 32999 36193 33008 36227
rect 32956 36184 33008 36193
rect 36176 36227 36228 36236
rect 36176 36193 36185 36227
rect 36185 36193 36219 36227
rect 36219 36193 36228 36227
rect 36176 36184 36228 36193
rect 27068 36159 27120 36168
rect 27068 36125 27077 36159
rect 27077 36125 27111 36159
rect 27111 36125 27120 36159
rect 27068 36116 27120 36125
rect 31760 36159 31812 36168
rect 31760 36125 31769 36159
rect 31769 36125 31803 36159
rect 31803 36125 31812 36159
rect 31760 36116 31812 36125
rect 33232 36159 33284 36168
rect 33232 36125 33266 36159
rect 33266 36125 33284 36159
rect 33232 36116 33284 36125
rect 41144 36116 41196 36168
rect 38108 36048 38160 36100
rect 40224 36048 40276 36100
rect 34796 35980 34848 36032
rect 37648 35980 37700 36032
rect 40132 36023 40184 36032
rect 40132 35989 40141 36023
rect 40141 35989 40175 36023
rect 40175 35989 40184 36023
rect 40132 35980 40184 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 26332 35776 26384 35828
rect 30012 35819 30064 35828
rect 30012 35785 30021 35819
rect 30021 35785 30055 35819
rect 30055 35785 30064 35819
rect 30012 35776 30064 35785
rect 30380 35819 30432 35828
rect 30380 35785 30389 35819
rect 30389 35785 30423 35819
rect 30423 35785 30432 35819
rect 30380 35776 30432 35785
rect 41144 35819 41196 35828
rect 41144 35785 41153 35819
rect 41153 35785 41187 35819
rect 41187 35785 41196 35819
rect 41144 35776 41196 35785
rect 23572 35640 23624 35692
rect 27068 35640 27120 35692
rect 30196 35683 30248 35692
rect 30196 35649 30205 35683
rect 30205 35649 30239 35683
rect 30239 35649 30248 35683
rect 30196 35640 30248 35649
rect 30564 35640 30616 35692
rect 40224 35708 40276 35760
rect 32956 35640 33008 35692
rect 22008 35479 22060 35488
rect 22008 35445 22017 35479
rect 22017 35445 22051 35479
rect 22051 35445 22060 35479
rect 22008 35436 22060 35445
rect 25596 35479 25648 35488
rect 25596 35445 25605 35479
rect 25605 35445 25639 35479
rect 25639 35445 25648 35479
rect 25596 35436 25648 35445
rect 34428 35479 34480 35488
rect 34428 35445 34437 35479
rect 34437 35445 34471 35479
rect 34471 35445 34480 35479
rect 34428 35436 34480 35445
rect 34520 35436 34572 35488
rect 36544 35479 36596 35488
rect 36544 35445 36553 35479
rect 36553 35445 36587 35479
rect 36587 35445 36596 35479
rect 36544 35436 36596 35445
rect 40040 35436 40092 35488
rect 40500 35436 40552 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 20076 35232 20128 35284
rect 23572 35275 23624 35284
rect 23572 35241 23581 35275
rect 23581 35241 23615 35275
rect 23615 35241 23624 35275
rect 23572 35232 23624 35241
rect 34796 35232 34848 35284
rect 38108 35275 38160 35284
rect 38108 35241 38117 35275
rect 38117 35241 38151 35275
rect 38151 35241 38160 35275
rect 38108 35232 38160 35241
rect 40224 35275 40276 35284
rect 40224 35241 40233 35275
rect 40233 35241 40267 35275
rect 40267 35241 40276 35275
rect 40224 35232 40276 35241
rect 23480 35096 23532 35148
rect 24584 35096 24636 35148
rect 32956 35139 33008 35148
rect 32956 35105 32965 35139
rect 32965 35105 32999 35139
rect 32999 35105 33008 35139
rect 32956 35096 33008 35105
rect 21364 35028 21416 35080
rect 23296 35071 23348 35080
rect 23296 35037 23305 35071
rect 23305 35037 23339 35071
rect 23339 35037 23348 35071
rect 23296 35028 23348 35037
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 34520 35096 34572 35148
rect 34428 35028 34480 35080
rect 35164 35071 35216 35080
rect 35164 35037 35173 35071
rect 35173 35037 35207 35071
rect 35207 35037 35216 35071
rect 35164 35028 35216 35037
rect 36268 35071 36320 35080
rect 36268 35037 36277 35071
rect 36277 35037 36311 35071
rect 36311 35037 36320 35071
rect 36268 35028 36320 35037
rect 36544 35071 36596 35080
rect 36544 35037 36578 35071
rect 36578 35037 36596 35071
rect 36544 35028 36596 35037
rect 40132 35028 40184 35080
rect 26608 34892 26660 34944
rect 37464 34892 37516 34944
rect 37740 34892 37792 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 20076 34731 20128 34740
rect 20076 34697 20085 34731
rect 20085 34697 20119 34731
rect 20119 34697 20128 34731
rect 20076 34688 20128 34697
rect 23296 34688 23348 34740
rect 26700 34688 26752 34740
rect 35164 34688 35216 34740
rect 22008 34620 22060 34672
rect 37464 34663 37516 34672
rect 37464 34629 37473 34663
rect 37473 34629 37507 34663
rect 37507 34629 37516 34663
rect 37464 34620 37516 34629
rect 22284 34595 22336 34604
rect 22284 34561 22318 34595
rect 22318 34561 22336 34595
rect 24584 34595 24636 34604
rect 22284 34552 22336 34561
rect 24584 34561 24593 34595
rect 24593 34561 24627 34595
rect 24627 34561 24636 34595
rect 24584 34552 24636 34561
rect 24860 34595 24912 34604
rect 24860 34561 24894 34595
rect 24894 34561 24912 34595
rect 24860 34552 24912 34561
rect 33876 34595 33928 34604
rect 33876 34561 33910 34595
rect 33910 34561 33928 34595
rect 37740 34595 37792 34604
rect 33876 34552 33928 34561
rect 37740 34561 37749 34595
rect 37749 34561 37783 34595
rect 37783 34561 37792 34595
rect 37740 34552 37792 34561
rect 21548 34484 21600 34536
rect 23480 34416 23532 34468
rect 32312 34416 32364 34468
rect 37556 34527 37608 34536
rect 37556 34493 37565 34527
rect 37565 34493 37599 34527
rect 37599 34493 37608 34527
rect 37556 34484 37608 34493
rect 39304 34484 39356 34536
rect 39764 34595 39816 34604
rect 39764 34561 39773 34595
rect 39773 34561 39807 34595
rect 39807 34561 39816 34595
rect 39948 34595 40000 34604
rect 39764 34552 39816 34561
rect 39948 34561 39957 34595
rect 39957 34561 39991 34595
rect 39991 34561 40000 34595
rect 39948 34552 40000 34561
rect 39856 34484 39908 34536
rect 41052 34484 41104 34536
rect 28172 34391 28224 34400
rect 28172 34357 28181 34391
rect 28181 34357 28215 34391
rect 28215 34357 28224 34391
rect 28172 34348 28224 34357
rect 28816 34391 28868 34400
rect 28816 34357 28825 34391
rect 28825 34357 28859 34391
rect 28859 34357 28868 34391
rect 28816 34348 28868 34357
rect 31208 34348 31260 34400
rect 36452 34391 36504 34400
rect 36452 34357 36461 34391
rect 36461 34357 36495 34391
rect 36495 34357 36504 34391
rect 36452 34348 36504 34357
rect 37648 34391 37700 34400
rect 37648 34357 37657 34391
rect 37657 34357 37691 34391
rect 37691 34357 37700 34391
rect 37648 34348 37700 34357
rect 38016 34348 38068 34400
rect 40224 34348 40276 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 22284 34144 22336 34196
rect 23388 34144 23440 34196
rect 26608 34187 26660 34196
rect 26608 34153 26617 34187
rect 26617 34153 26651 34187
rect 26651 34153 26660 34187
rect 26608 34144 26660 34153
rect 27068 34187 27120 34196
rect 27068 34153 27077 34187
rect 27077 34153 27111 34187
rect 27111 34153 27120 34187
rect 27068 34144 27120 34153
rect 33048 34187 33100 34196
rect 33048 34153 33057 34187
rect 33057 34153 33091 34187
rect 33091 34153 33100 34187
rect 33048 34144 33100 34153
rect 33876 34144 33928 34196
rect 37556 34187 37608 34196
rect 37556 34153 37565 34187
rect 37565 34153 37599 34187
rect 37599 34153 37608 34187
rect 37556 34144 37608 34153
rect 39304 34187 39356 34196
rect 39304 34153 39313 34187
rect 39313 34153 39347 34187
rect 39347 34153 39356 34187
rect 39304 34144 39356 34153
rect 39488 34187 39540 34196
rect 39488 34153 39497 34187
rect 39497 34153 39531 34187
rect 39531 34153 39540 34187
rect 39488 34144 39540 34153
rect 40224 34187 40276 34196
rect 40224 34153 40233 34187
rect 40233 34153 40267 34187
rect 40267 34153 40276 34187
rect 40224 34144 40276 34153
rect 21548 34051 21600 34060
rect 21548 34017 21557 34051
rect 21557 34017 21591 34051
rect 21591 34017 21600 34051
rect 21548 34008 21600 34017
rect 24584 34008 24636 34060
rect 24860 33940 24912 33992
rect 26700 34051 26752 34060
rect 26700 34017 26709 34051
rect 26709 34017 26743 34051
rect 26743 34017 26752 34051
rect 26700 34008 26752 34017
rect 27804 34051 27856 34060
rect 27804 34017 27813 34051
rect 27813 34017 27847 34051
rect 27847 34017 27856 34051
rect 27804 34008 27856 34017
rect 28816 33940 28868 33992
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 31024 33940 31076 33992
rect 31208 33983 31260 33992
rect 31208 33949 31242 33983
rect 31242 33949 31260 33983
rect 31208 33940 31260 33949
rect 32496 33940 32548 33992
rect 36268 33940 36320 33992
rect 38016 33983 38068 33992
rect 22008 33872 22060 33924
rect 26148 33872 26200 33924
rect 26240 33872 26292 33924
rect 31760 33872 31812 33924
rect 36452 33915 36504 33924
rect 36452 33881 36486 33915
rect 36486 33881 36504 33915
rect 36452 33872 36504 33881
rect 38016 33949 38025 33983
rect 38025 33949 38059 33983
rect 38059 33949 38068 33983
rect 38016 33940 38068 33949
rect 38200 33983 38252 33992
rect 38200 33949 38209 33983
rect 38209 33949 38243 33983
rect 38243 33949 38252 33983
rect 38200 33940 38252 33949
rect 38384 33872 38436 33924
rect 39764 34008 39816 34060
rect 29736 33804 29788 33856
rect 33232 33847 33284 33856
rect 33232 33813 33241 33847
rect 33241 33813 33275 33847
rect 33275 33813 33284 33847
rect 33232 33804 33284 33813
rect 40132 33872 40184 33924
rect 40316 33940 40368 33992
rect 41052 33983 41104 33992
rect 41052 33949 41061 33983
rect 41061 33949 41095 33983
rect 41095 33949 41104 33983
rect 41052 33940 41104 33949
rect 41236 33983 41288 33992
rect 41236 33949 41245 33983
rect 41245 33949 41279 33983
rect 41279 33949 41288 33983
rect 41236 33940 41288 33949
rect 43444 33983 43496 33992
rect 43444 33949 43453 33983
rect 43453 33949 43487 33983
rect 43487 33949 43496 33983
rect 43444 33940 43496 33949
rect 39304 33847 39356 33856
rect 39304 33813 39329 33847
rect 39329 33813 39356 33847
rect 40040 33847 40092 33856
rect 39304 33804 39356 33813
rect 40040 33813 40049 33847
rect 40049 33813 40083 33847
rect 40083 33813 40092 33847
rect 40040 33804 40092 33813
rect 40316 33804 40368 33856
rect 43260 33847 43312 33856
rect 43260 33813 43269 33847
rect 43269 33813 43303 33847
rect 43303 33813 43312 33847
rect 43260 33804 43312 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 24584 33600 24636 33652
rect 30472 33600 30524 33652
rect 31760 33643 31812 33652
rect 28172 33575 28224 33584
rect 28172 33541 28206 33575
rect 28206 33541 28224 33575
rect 28172 33532 28224 33541
rect 22008 33507 22060 33516
rect 22008 33473 22017 33507
rect 22017 33473 22051 33507
rect 22051 33473 22060 33507
rect 22008 33464 22060 33473
rect 24216 33464 24268 33516
rect 26424 33464 26476 33516
rect 31024 33532 31076 33584
rect 31760 33609 31769 33643
rect 31769 33609 31803 33643
rect 31803 33609 31812 33643
rect 31760 33600 31812 33609
rect 33048 33600 33100 33652
rect 39304 33600 39356 33652
rect 39948 33600 40000 33652
rect 41236 33600 41288 33652
rect 43260 33575 43312 33584
rect 43260 33541 43294 33575
rect 43294 33541 43312 33575
rect 43260 33532 43312 33541
rect 30932 33464 30984 33516
rect 39212 33464 39264 33516
rect 40500 33507 40552 33516
rect 40500 33473 40509 33507
rect 40509 33473 40543 33507
rect 40543 33473 40552 33507
rect 40500 33464 40552 33473
rect 40776 33507 40828 33516
rect 40776 33473 40810 33507
rect 40810 33473 40828 33507
rect 40776 33464 40828 33473
rect 26148 33439 26200 33448
rect 26148 33405 26157 33439
rect 26157 33405 26191 33439
rect 26191 33405 26200 33439
rect 26148 33396 26200 33405
rect 27804 33396 27856 33448
rect 32312 33439 32364 33448
rect 32312 33405 32321 33439
rect 32321 33405 32355 33439
rect 32355 33405 32364 33439
rect 32312 33396 32364 33405
rect 38384 33396 38436 33448
rect 42800 33396 42852 33448
rect 27896 33260 27948 33312
rect 29276 33303 29328 33312
rect 29276 33269 29285 33303
rect 29285 33269 29319 33303
rect 29319 33269 29328 33303
rect 29276 33260 29328 33269
rect 31392 33260 31444 33312
rect 44364 33303 44416 33312
rect 44364 33269 44373 33303
rect 44373 33269 44407 33303
rect 44407 33269 44416 33303
rect 44364 33260 44416 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 26240 33056 26292 33108
rect 26424 33099 26476 33108
rect 26424 33065 26433 33099
rect 26433 33065 26467 33099
rect 26467 33065 26476 33099
rect 26424 33056 26476 33065
rect 29736 33099 29788 33108
rect 29736 33065 29745 33099
rect 29745 33065 29779 33099
rect 29779 33065 29788 33099
rect 29736 33056 29788 33065
rect 32496 33099 32548 33108
rect 32496 33065 32505 33099
rect 32505 33065 32539 33099
rect 32539 33065 32548 33099
rect 32496 33056 32548 33065
rect 33232 33056 33284 33108
rect 38200 33056 38252 33108
rect 39212 33099 39264 33108
rect 39212 33065 39221 33099
rect 39221 33065 39255 33099
rect 39255 33065 39264 33099
rect 39212 33056 39264 33065
rect 40316 33056 40368 33108
rect 40776 33056 40828 33108
rect 43444 33056 43496 33108
rect 23296 32920 23348 32972
rect 24584 32963 24636 32972
rect 24584 32929 24593 32963
rect 24593 32929 24627 32963
rect 24627 32929 24636 32963
rect 24584 32920 24636 32929
rect 43352 33031 43404 33040
rect 27804 32895 27856 32904
rect 27804 32861 27813 32895
rect 27813 32861 27847 32895
rect 27847 32861 27856 32895
rect 27804 32852 27856 32861
rect 27896 32852 27948 32904
rect 29276 32852 29328 32904
rect 31116 32895 31168 32904
rect 31116 32861 31125 32895
rect 31125 32861 31159 32895
rect 31159 32861 31168 32895
rect 31116 32852 31168 32861
rect 32312 32852 32364 32904
rect 33140 32895 33192 32904
rect 33140 32861 33149 32895
rect 33149 32861 33183 32895
rect 33183 32861 33192 32895
rect 33140 32852 33192 32861
rect 33232 32895 33284 32904
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 35440 32852 35492 32904
rect 40040 32920 40092 32972
rect 43352 32997 43361 33031
rect 43361 32997 43395 33031
rect 43395 32997 43404 33031
rect 43352 32988 43404 32997
rect 24860 32827 24912 32836
rect 24860 32793 24894 32827
rect 24894 32793 24912 32827
rect 24860 32784 24912 32793
rect 28908 32784 28960 32836
rect 31392 32827 31444 32836
rect 31392 32793 31426 32827
rect 31426 32793 31444 32827
rect 31392 32784 31444 32793
rect 40132 32784 40184 32836
rect 42064 32784 42116 32836
rect 43628 32784 43680 32836
rect 44364 32784 44416 32836
rect 44548 32784 44600 32836
rect 40224 32759 40276 32768
rect 40224 32725 40249 32759
rect 40249 32725 40276 32759
rect 40224 32716 40276 32725
rect 41144 32716 41196 32768
rect 42524 32716 42576 32768
rect 45376 32759 45428 32768
rect 45376 32725 45401 32759
rect 45401 32725 45428 32759
rect 45376 32716 45428 32725
rect 46020 32716 46072 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 33232 32512 33284 32564
rect 40224 32512 40276 32564
rect 42064 32555 42116 32564
rect 42064 32521 42073 32555
rect 42073 32521 42107 32555
rect 42107 32521 42116 32555
rect 42064 32512 42116 32521
rect 42524 32512 42576 32564
rect 42708 32512 42760 32564
rect 43720 32512 43772 32564
rect 36912 32487 36964 32496
rect 36912 32453 36921 32487
rect 36921 32453 36955 32487
rect 36955 32453 36964 32487
rect 36912 32444 36964 32453
rect 39396 32444 39448 32496
rect 44456 32444 44508 32496
rect 24860 32376 24912 32428
rect 30932 32376 30984 32428
rect 35808 32419 35860 32428
rect 35808 32385 35817 32419
rect 35817 32385 35851 32419
rect 35851 32385 35860 32419
rect 35808 32376 35860 32385
rect 36452 32376 36504 32428
rect 39856 32376 39908 32428
rect 41144 32419 41196 32428
rect 35992 32351 36044 32360
rect 35992 32317 36001 32351
rect 36001 32317 36035 32351
rect 36035 32317 36044 32351
rect 35992 32308 36044 32317
rect 41144 32385 41153 32419
rect 41153 32385 41187 32419
rect 41187 32385 41196 32419
rect 41144 32376 41196 32385
rect 42800 32419 42852 32428
rect 41236 32308 41288 32360
rect 42800 32385 42809 32419
rect 42809 32385 42843 32419
rect 42843 32385 42852 32419
rect 42800 32376 42852 32385
rect 43628 32376 43680 32428
rect 46204 32419 46256 32428
rect 42708 32308 42760 32360
rect 46204 32385 46222 32419
rect 46222 32385 46256 32419
rect 46204 32376 46256 32385
rect 46480 32351 46532 32360
rect 46480 32317 46489 32351
rect 46489 32317 46523 32351
rect 46523 32317 46532 32351
rect 46480 32308 46532 32317
rect 43628 32240 43680 32292
rect 44088 32283 44140 32292
rect 44088 32249 44097 32283
rect 44097 32249 44131 32283
rect 44131 32249 44140 32283
rect 44088 32240 44140 32249
rect 27620 32172 27672 32224
rect 35348 32172 35400 32224
rect 36084 32215 36136 32224
rect 36084 32181 36093 32215
rect 36093 32181 36127 32215
rect 36127 32181 36136 32215
rect 36084 32172 36136 32181
rect 38384 32172 38436 32224
rect 41788 32172 41840 32224
rect 43536 32215 43588 32224
rect 43536 32181 43545 32215
rect 43545 32181 43579 32215
rect 43579 32181 43588 32215
rect 43536 32172 43588 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 24584 31832 24636 31884
rect 27804 31968 27856 32020
rect 28908 32011 28960 32020
rect 28908 31977 28917 32011
rect 28917 31977 28951 32011
rect 28951 31977 28960 32011
rect 28908 31968 28960 31977
rect 36084 31968 36136 32020
rect 42800 31968 42852 32020
rect 44548 32011 44600 32020
rect 44548 31977 44557 32011
rect 44557 31977 44591 32011
rect 44591 31977 44600 32011
rect 44548 31968 44600 31977
rect 45376 31968 45428 32020
rect 46204 32011 46256 32020
rect 46204 31977 46213 32011
rect 46213 31977 46247 32011
rect 46247 31977 46256 32011
rect 46204 31968 46256 31977
rect 42892 31832 42944 31884
rect 43720 31875 43772 31884
rect 43720 31841 43729 31875
rect 43729 31841 43763 31875
rect 43763 31841 43772 31875
rect 43720 31832 43772 31841
rect 44088 31832 44140 31884
rect 27620 31764 27672 31816
rect 34704 31764 34756 31816
rect 34796 31764 34848 31816
rect 35440 31764 35492 31816
rect 36728 31807 36780 31816
rect 36728 31773 36737 31807
rect 36737 31773 36771 31807
rect 36771 31773 36780 31807
rect 36728 31764 36780 31773
rect 43628 31807 43680 31816
rect 41788 31696 41840 31748
rect 43628 31773 43637 31807
rect 43637 31773 43671 31807
rect 43671 31773 43680 31807
rect 43628 31764 43680 31773
rect 46020 31807 46072 31816
rect 46020 31773 46029 31807
rect 46029 31773 46063 31807
rect 46063 31773 46072 31807
rect 46020 31764 46072 31773
rect 42616 31628 42668 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 36452 31467 36504 31476
rect 36452 31433 36461 31467
rect 36461 31433 36495 31467
rect 36495 31433 36504 31467
rect 36452 31424 36504 31433
rect 32496 31356 32548 31408
rect 36912 31356 36964 31408
rect 43536 31356 43588 31408
rect 44456 31356 44508 31408
rect 23296 31288 23348 31340
rect 25136 31288 25188 31340
rect 34704 31288 34756 31340
rect 41880 31331 41932 31340
rect 41880 31297 41889 31331
rect 41889 31297 41923 31331
rect 41923 31297 41932 31331
rect 41880 31288 41932 31297
rect 34796 31220 34848 31272
rect 42616 31152 42668 31204
rect 46480 31152 46532 31204
rect 24584 31127 24636 31136
rect 24584 31093 24593 31127
rect 24593 31093 24627 31127
rect 24627 31093 24636 31127
rect 24584 31084 24636 31093
rect 30840 31127 30892 31136
rect 30840 31093 30849 31127
rect 30849 31093 30883 31127
rect 30883 31093 30892 31127
rect 30840 31084 30892 31093
rect 31484 31127 31536 31136
rect 31484 31093 31493 31127
rect 31493 31093 31527 31127
rect 31527 31093 31536 31127
rect 31484 31084 31536 31093
rect 42708 31084 42760 31136
rect 43628 31127 43680 31136
rect 43628 31093 43637 31127
rect 43637 31093 43671 31127
rect 43671 31093 43680 31127
rect 43628 31084 43680 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 33140 30880 33192 30932
rect 35992 30880 36044 30932
rect 44088 30880 44140 30932
rect 44456 30923 44508 30932
rect 44456 30889 44465 30923
rect 44465 30889 44499 30923
rect 44499 30889 44508 30923
rect 44456 30880 44508 30889
rect 31760 30744 31812 30796
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 30380 30676 30432 30728
rect 31116 30676 31168 30728
rect 31392 30676 31444 30728
rect 32680 30719 32732 30728
rect 32680 30685 32689 30719
rect 32689 30685 32723 30719
rect 32723 30685 32732 30719
rect 32680 30676 32732 30685
rect 34796 30676 34848 30728
rect 42616 30719 42668 30728
rect 42616 30685 42625 30719
rect 42625 30685 42659 30719
rect 42659 30685 42668 30719
rect 42616 30676 42668 30685
rect 42708 30676 42760 30728
rect 30840 30651 30892 30660
rect 30840 30617 30874 30651
rect 30874 30617 30892 30651
rect 30840 30608 30892 30617
rect 32404 30651 32456 30660
rect 32404 30617 32413 30651
rect 32413 30617 32447 30651
rect 32447 30617 32456 30651
rect 32404 30608 32456 30617
rect 35348 30608 35400 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 31392 30336 31444 30388
rect 34796 30336 34848 30388
rect 41880 30336 41932 30388
rect 23572 30311 23624 30320
rect 23572 30277 23606 30311
rect 23606 30277 23624 30311
rect 23572 30268 23624 30277
rect 31484 30268 31536 30320
rect 36728 30268 36780 30320
rect 42892 30311 42944 30320
rect 42892 30277 42901 30311
rect 42901 30277 42935 30311
rect 42935 30277 42944 30311
rect 42892 30268 42944 30277
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 30380 30243 30432 30252
rect 30380 30209 30389 30243
rect 30389 30209 30423 30243
rect 30423 30209 30432 30243
rect 30380 30200 30432 30209
rect 43076 30200 43128 30252
rect 43628 30200 43680 30252
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 38384 30132 38436 30184
rect 31760 30107 31812 30116
rect 31760 30073 31769 30107
rect 31769 30073 31803 30107
rect 31803 30073 31812 30107
rect 31760 30064 31812 30073
rect 22836 30039 22888 30048
rect 22836 30005 22845 30039
rect 22845 30005 22879 30039
rect 22879 30005 22888 30039
rect 22836 29996 22888 30005
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 31944 29996 31996 30048
rect 35808 29996 35860 30048
rect 43352 29996 43404 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 24676 29835 24728 29844
rect 24676 29801 24685 29835
rect 24685 29801 24719 29835
rect 24719 29801 24728 29835
rect 24676 29792 24728 29801
rect 32680 29792 32732 29844
rect 24584 29656 24636 29708
rect 31392 29699 31444 29708
rect 31392 29665 31401 29699
rect 31401 29665 31435 29699
rect 31435 29665 31444 29699
rect 31392 29656 31444 29665
rect 23296 29588 23348 29640
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 30288 29588 30340 29640
rect 31944 29588 31996 29640
rect 43904 29588 43956 29640
rect 46480 29588 46532 29640
rect 25136 29452 25188 29504
rect 44640 29452 44692 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 24860 29248 24912 29300
rect 32404 29248 32456 29300
rect 43904 29291 43956 29300
rect 43904 29257 43913 29291
rect 43913 29257 43947 29291
rect 43947 29257 43956 29291
rect 43904 29248 43956 29257
rect 22836 29180 22888 29232
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 30380 29180 30432 29232
rect 45284 29223 45336 29232
rect 30288 29155 30340 29164
rect 30288 29121 30322 29155
rect 30322 29121 30340 29155
rect 30288 29112 30340 29121
rect 43076 29155 43128 29164
rect 43076 29121 43085 29155
rect 43085 29121 43119 29155
rect 43119 29121 43128 29155
rect 43076 29112 43128 29121
rect 44548 29155 44600 29164
rect 44548 29121 44557 29155
rect 44557 29121 44591 29155
rect 44591 29121 44600 29155
rect 44732 29155 44784 29164
rect 44548 29112 44600 29121
rect 44732 29121 44741 29155
rect 44741 29121 44775 29155
rect 44775 29121 44784 29155
rect 44732 29112 44784 29121
rect 45284 29189 45293 29223
rect 45293 29189 45327 29223
rect 45327 29189 45336 29223
rect 45284 29180 45336 29189
rect 45376 29180 45428 29232
rect 43260 29044 43312 29096
rect 35440 28976 35492 29028
rect 38660 29019 38712 29028
rect 38660 28985 38669 29019
rect 38669 28985 38703 29019
rect 38703 28985 38712 29019
rect 38660 28976 38712 28985
rect 17316 28951 17368 28960
rect 17316 28917 17325 28951
rect 17325 28917 17359 28951
rect 17359 28917 17368 28951
rect 17316 28908 17368 28917
rect 18328 28951 18380 28960
rect 18328 28917 18337 28951
rect 18337 28917 18371 28951
rect 18371 28917 18380 28951
rect 18328 28908 18380 28917
rect 36176 28951 36228 28960
rect 36176 28917 36185 28951
rect 36185 28917 36219 28951
rect 36219 28917 36228 28951
rect 36176 28908 36228 28917
rect 42892 28908 42944 28960
rect 43352 28908 43404 28960
rect 46296 28951 46348 28960
rect 46296 28917 46305 28951
rect 46305 28917 46339 28951
rect 46339 28917 46348 28951
rect 46296 28908 46348 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 31760 28704 31812 28756
rect 32496 28747 32548 28756
rect 32496 28713 32505 28747
rect 32505 28713 32539 28747
rect 32539 28713 32548 28747
rect 32496 28704 32548 28713
rect 44640 28611 44692 28620
rect 44640 28577 44649 28611
rect 44649 28577 44683 28611
rect 44683 28577 44692 28611
rect 44640 28568 44692 28577
rect 16948 28500 17000 28552
rect 17316 28543 17368 28552
rect 17316 28509 17350 28543
rect 17350 28509 17368 28543
rect 17316 28500 17368 28509
rect 24860 28500 24912 28552
rect 34796 28500 34848 28552
rect 35072 28500 35124 28552
rect 38752 28543 38804 28552
rect 38752 28509 38761 28543
rect 38761 28509 38795 28543
rect 38795 28509 38804 28543
rect 38752 28500 38804 28509
rect 42984 28543 43036 28552
rect 42984 28509 42993 28543
rect 42993 28509 43027 28543
rect 43027 28509 43036 28543
rect 42984 28500 43036 28509
rect 43260 28543 43312 28552
rect 43260 28509 43269 28543
rect 43269 28509 43303 28543
rect 43303 28509 43312 28543
rect 43260 28500 43312 28509
rect 43720 28500 43772 28552
rect 44732 28500 44784 28552
rect 20076 28364 20128 28416
rect 30656 28407 30708 28416
rect 30656 28373 30665 28407
rect 30665 28373 30699 28407
rect 30699 28373 30708 28407
rect 36176 28432 36228 28484
rect 43076 28432 43128 28484
rect 46296 28543 46348 28552
rect 46296 28509 46314 28543
rect 46314 28509 46348 28543
rect 46296 28500 46348 28509
rect 46480 28500 46532 28552
rect 30656 28364 30708 28373
rect 37648 28364 37700 28416
rect 42800 28407 42852 28416
rect 42800 28373 42809 28407
rect 42809 28373 42843 28407
rect 42843 28373 42852 28407
rect 42800 28364 42852 28373
rect 45192 28407 45244 28416
rect 45192 28373 45201 28407
rect 45201 28373 45235 28407
rect 45235 28373 45244 28407
rect 45192 28364 45244 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 18328 28135 18380 28144
rect 18328 28101 18362 28135
rect 18362 28101 18380 28135
rect 18328 28092 18380 28101
rect 19340 28024 19392 28076
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 38752 28092 38804 28144
rect 42984 28160 43036 28212
rect 43904 28160 43956 28212
rect 45376 28160 45428 28212
rect 43076 28092 43128 28144
rect 44916 28135 44968 28144
rect 44916 28101 44925 28135
rect 44925 28101 44959 28135
rect 44959 28101 44968 28135
rect 44916 28092 44968 28101
rect 16948 27956 17000 28008
rect 35072 28067 35124 28076
rect 35072 28033 35081 28067
rect 35081 28033 35115 28067
rect 35115 28033 35124 28067
rect 35072 28024 35124 28033
rect 37648 28067 37700 28076
rect 37648 28033 37657 28067
rect 37657 28033 37691 28067
rect 37691 28033 37700 28067
rect 37648 28024 37700 28033
rect 37740 28067 37792 28076
rect 37740 28033 37749 28067
rect 37749 28033 37783 28067
rect 37783 28033 37792 28067
rect 38384 28067 38436 28076
rect 37740 28024 37792 28033
rect 38384 28033 38393 28067
rect 38393 28033 38427 28067
rect 38427 28033 38436 28067
rect 38384 28024 38436 28033
rect 41880 28067 41932 28076
rect 41880 28033 41889 28067
rect 41889 28033 41923 28067
rect 41923 28033 41932 28067
rect 41880 28024 41932 28033
rect 42616 28067 42668 28076
rect 42616 28033 42625 28067
rect 42625 28033 42659 28067
rect 42659 28033 42668 28067
rect 42616 28024 42668 28033
rect 45192 28024 45244 28076
rect 45376 28024 45428 28076
rect 3424 27820 3476 27872
rect 16764 27820 16816 27872
rect 17316 27863 17368 27872
rect 17316 27829 17325 27863
rect 17325 27829 17359 27863
rect 17359 27829 17368 27863
rect 17316 27820 17368 27829
rect 30656 27888 30708 27940
rect 19892 27863 19944 27872
rect 19892 27829 19901 27863
rect 19901 27829 19935 27863
rect 19935 27829 19944 27863
rect 19892 27820 19944 27829
rect 20352 27863 20404 27872
rect 20352 27829 20361 27863
rect 20361 27829 20395 27863
rect 20395 27829 20404 27863
rect 20352 27820 20404 27829
rect 20996 27820 21048 27872
rect 24676 27863 24728 27872
rect 24676 27829 24685 27863
rect 24685 27829 24719 27863
rect 24719 27829 24728 27863
rect 24676 27820 24728 27829
rect 25596 27863 25648 27872
rect 25596 27829 25605 27863
rect 25605 27829 25639 27863
rect 25639 27829 25648 27863
rect 25596 27820 25648 27829
rect 28632 27863 28684 27872
rect 28632 27829 28641 27863
rect 28641 27829 28675 27863
rect 28675 27829 28684 27863
rect 28632 27820 28684 27829
rect 31944 27820 31996 27872
rect 32956 27863 33008 27872
rect 32956 27829 32965 27863
rect 32965 27829 32999 27863
rect 32999 27829 33008 27863
rect 32956 27820 33008 27829
rect 37464 27863 37516 27872
rect 37464 27829 37473 27863
rect 37473 27829 37507 27863
rect 37507 27829 37516 27863
rect 37464 27820 37516 27829
rect 37924 27863 37976 27872
rect 37924 27829 37933 27863
rect 37933 27829 37967 27863
rect 37967 27829 37976 27863
rect 37924 27820 37976 27829
rect 40040 27820 40092 27872
rect 40132 27820 40184 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 41880 27616 41932 27668
rect 42892 27616 42944 27668
rect 43168 27616 43220 27668
rect 19892 27548 19944 27600
rect 37464 27548 37516 27600
rect 45284 27591 45336 27600
rect 45284 27557 45293 27591
rect 45293 27557 45327 27591
rect 45327 27557 45336 27591
rect 45284 27548 45336 27557
rect 16948 27412 17000 27464
rect 17316 27455 17368 27464
rect 17316 27421 17350 27455
rect 17350 27421 17368 27455
rect 17316 27412 17368 27421
rect 20628 27412 20680 27464
rect 20996 27455 21048 27464
rect 20996 27421 21030 27455
rect 21030 27421 21048 27455
rect 20996 27412 21048 27421
rect 23204 27455 23256 27464
rect 23204 27421 23213 27455
rect 23213 27421 23247 27455
rect 23247 27421 23256 27455
rect 23204 27412 23256 27421
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 31208 27455 31260 27464
rect 31208 27421 31217 27455
rect 31217 27421 31251 27455
rect 31251 27421 31260 27455
rect 31208 27412 31260 27421
rect 32312 27412 32364 27464
rect 34520 27412 34572 27464
rect 35440 27455 35492 27464
rect 35440 27421 35474 27455
rect 35474 27421 35492 27455
rect 35440 27412 35492 27421
rect 37004 27455 37056 27464
rect 37004 27421 37013 27455
rect 37013 27421 37047 27455
rect 37047 27421 37056 27455
rect 37004 27412 37056 27421
rect 38108 27455 38160 27464
rect 38108 27421 38117 27455
rect 38117 27421 38151 27455
rect 38151 27421 38160 27455
rect 38108 27412 38160 27421
rect 42064 27412 42116 27464
rect 44916 27412 44968 27464
rect 45376 27455 45428 27464
rect 45376 27421 45385 27455
rect 45385 27421 45419 27455
rect 45419 27421 45428 27455
rect 45376 27412 45428 27421
rect 27344 27344 27396 27396
rect 31944 27387 31996 27396
rect 31944 27353 31978 27387
rect 31978 27353 31996 27387
rect 31944 27344 31996 27353
rect 40132 27344 40184 27396
rect 40316 27387 40368 27396
rect 40316 27353 40350 27387
rect 40350 27353 40368 27387
rect 40316 27344 40368 27353
rect 42800 27344 42852 27396
rect 43720 27387 43772 27396
rect 43720 27353 43747 27387
rect 43747 27353 43772 27387
rect 43720 27344 43772 27353
rect 43904 27387 43956 27396
rect 43904 27353 43913 27387
rect 43913 27353 43947 27387
rect 43947 27353 43956 27387
rect 43904 27344 43956 27353
rect 22284 27276 22336 27328
rect 25044 27276 25096 27328
rect 29092 27319 29144 27328
rect 29092 27285 29101 27319
rect 29101 27285 29135 27319
rect 29135 27285 29144 27319
rect 29092 27276 29144 27285
rect 33416 27276 33468 27328
rect 39488 27319 39540 27328
rect 39488 27285 39497 27319
rect 39497 27285 39531 27319
rect 39531 27285 39540 27319
rect 39488 27276 39540 27285
rect 40500 27276 40552 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 19340 27072 19392 27124
rect 31208 27072 31260 27124
rect 16764 27004 16816 27056
rect 23204 27004 23256 27056
rect 25596 27004 25648 27056
rect 16948 26936 17000 26988
rect 27712 26936 27764 26988
rect 32312 27004 32364 27056
rect 37740 27072 37792 27124
rect 43904 27072 43956 27124
rect 32956 26936 33008 26988
rect 38108 27004 38160 27056
rect 38660 27047 38712 27056
rect 37004 26936 37056 26988
rect 38660 27013 38694 27047
rect 38694 27013 38712 27047
rect 38660 27004 38712 27013
rect 39488 27004 39540 27056
rect 40316 27004 40368 27056
rect 43720 27004 43772 27056
rect 40500 26979 40552 26988
rect 20628 26868 20680 26920
rect 24584 26911 24636 26920
rect 24584 26877 24593 26911
rect 24593 26877 24627 26911
rect 24627 26877 24636 26911
rect 24584 26868 24636 26877
rect 32312 26911 32364 26920
rect 32312 26877 32321 26911
rect 32321 26877 32355 26911
rect 32355 26877 32364 26911
rect 32312 26868 32364 26877
rect 40500 26945 40509 26979
rect 40509 26945 40543 26979
rect 40543 26945 40552 26979
rect 40500 26936 40552 26945
rect 43076 26979 43128 26988
rect 43076 26945 43085 26979
rect 43085 26945 43119 26979
rect 43119 26945 43128 26979
rect 43076 26936 43128 26945
rect 58072 26979 58124 26988
rect 58072 26945 58081 26979
rect 58081 26945 58115 26979
rect 58115 26945 58124 26979
rect 58072 26936 58124 26945
rect 42984 26911 43036 26920
rect 42984 26877 42993 26911
rect 42993 26877 43027 26911
rect 43027 26877 43036 26911
rect 42984 26868 43036 26877
rect 43720 26868 43772 26920
rect 43444 26800 43496 26852
rect 24952 26732 25004 26784
rect 25320 26732 25372 26784
rect 27896 26732 27948 26784
rect 29828 26732 29880 26784
rect 33324 26732 33376 26784
rect 33600 26732 33652 26784
rect 40040 26732 40092 26784
rect 40684 26775 40736 26784
rect 40684 26741 40693 26775
rect 40693 26741 40727 26775
rect 40727 26741 40736 26775
rect 40684 26732 40736 26741
rect 43352 26775 43404 26784
rect 43352 26741 43361 26775
rect 43361 26741 43395 26775
rect 43395 26741 43404 26775
rect 43352 26732 43404 26741
rect 44364 26775 44416 26784
rect 44364 26741 44373 26775
rect 44373 26741 44407 26775
rect 44407 26741 44416 26775
rect 44364 26732 44416 26741
rect 58256 26775 58308 26784
rect 58256 26741 58265 26775
rect 58265 26741 58299 26775
rect 58299 26741 58308 26775
rect 58256 26732 58308 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 20628 26528 20680 26580
rect 27344 26571 27396 26580
rect 27344 26537 27353 26571
rect 27353 26537 27387 26571
rect 27387 26537 27396 26571
rect 27344 26528 27396 26537
rect 40684 26528 40736 26580
rect 43168 26528 43220 26580
rect 43444 26571 43496 26580
rect 43444 26537 43453 26571
rect 43453 26537 43487 26571
rect 43487 26537 43496 26571
rect 43444 26528 43496 26537
rect 45560 26528 45612 26580
rect 24584 26435 24636 26444
rect 24584 26401 24593 26435
rect 24593 26401 24627 26435
rect 24627 26401 24636 26435
rect 24584 26392 24636 26401
rect 27712 26392 27764 26444
rect 37832 26392 37884 26444
rect 13544 26367 13596 26376
rect 13544 26333 13553 26367
rect 13553 26333 13587 26367
rect 13587 26333 13596 26367
rect 13544 26324 13596 26333
rect 24860 26367 24912 26376
rect 24860 26333 24894 26367
rect 24894 26333 24912 26367
rect 24860 26324 24912 26333
rect 28632 26324 28684 26376
rect 31760 26324 31812 26376
rect 32312 26367 32364 26376
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 34520 26324 34572 26376
rect 37924 26324 37976 26376
rect 17960 26256 18012 26308
rect 23112 26256 23164 26308
rect 32588 26299 32640 26308
rect 32588 26265 32622 26299
rect 32622 26265 32640 26299
rect 32588 26256 32640 26265
rect 13360 26231 13412 26240
rect 13360 26197 13369 26231
rect 13369 26197 13403 26231
rect 13403 26197 13412 26231
rect 13360 26188 13412 26197
rect 25228 26188 25280 26240
rect 30012 26188 30064 26240
rect 33692 26231 33744 26240
rect 33692 26197 33701 26231
rect 33701 26197 33735 26231
rect 33735 26197 33744 26231
rect 33692 26188 33744 26197
rect 42064 26367 42116 26376
rect 42064 26333 42073 26367
rect 42073 26333 42107 26367
rect 42107 26333 42116 26367
rect 42064 26324 42116 26333
rect 42708 26324 42760 26376
rect 43168 26324 43220 26376
rect 43996 26367 44048 26376
rect 43996 26333 44005 26367
rect 44005 26333 44039 26367
rect 44039 26333 44048 26367
rect 43996 26324 44048 26333
rect 41880 26256 41932 26308
rect 44180 26299 44232 26308
rect 44180 26265 44189 26299
rect 44189 26265 44223 26299
rect 44223 26265 44232 26299
rect 44180 26256 44232 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 41880 26027 41932 26036
rect 13360 25916 13412 25968
rect 41880 25993 41889 26027
rect 41889 25993 41923 26027
rect 41923 25993 41932 26027
rect 41880 25984 41932 25993
rect 24952 25916 25004 25968
rect 27712 25916 27764 25968
rect 15844 25780 15896 25832
rect 20352 25848 20404 25900
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 22192 25848 22244 25900
rect 19340 25780 19392 25832
rect 22100 25823 22152 25832
rect 22100 25789 22109 25823
rect 22109 25789 22143 25823
rect 22143 25789 22152 25823
rect 22100 25780 22152 25789
rect 24860 25848 24912 25900
rect 25136 25848 25188 25900
rect 25320 25891 25372 25900
rect 25320 25857 25329 25891
rect 25329 25857 25363 25891
rect 25363 25857 25372 25891
rect 25320 25848 25372 25857
rect 29920 25916 29972 25968
rect 33692 25959 33744 25968
rect 33692 25925 33701 25959
rect 33701 25925 33735 25959
rect 33735 25925 33744 25959
rect 33692 25916 33744 25925
rect 42708 25916 42760 25968
rect 45560 25959 45612 25968
rect 27896 25848 27948 25900
rect 29092 25848 29144 25900
rect 30012 25891 30064 25900
rect 30012 25857 30021 25891
rect 30021 25857 30055 25891
rect 30055 25857 30064 25891
rect 30012 25848 30064 25857
rect 32588 25848 32640 25900
rect 33324 25848 33376 25900
rect 42064 25891 42116 25900
rect 42064 25857 42073 25891
rect 42073 25857 42107 25891
rect 42107 25857 42116 25891
rect 42064 25848 42116 25857
rect 43444 25891 43496 25900
rect 43444 25857 43453 25891
rect 43453 25857 43487 25891
rect 43487 25857 43496 25891
rect 43444 25848 43496 25857
rect 43996 25848 44048 25900
rect 44180 25848 44232 25900
rect 44364 25891 44416 25900
rect 44364 25857 44373 25891
rect 44373 25857 44407 25891
rect 44407 25857 44416 25891
rect 44364 25848 44416 25857
rect 45560 25925 45594 25959
rect 45594 25925 45612 25959
rect 45560 25916 45612 25925
rect 24952 25780 25004 25832
rect 25228 25823 25280 25832
rect 25228 25789 25237 25823
rect 25237 25789 25271 25823
rect 25271 25789 25280 25823
rect 25228 25780 25280 25789
rect 29828 25823 29880 25832
rect 29828 25789 29837 25823
rect 29837 25789 29871 25823
rect 29871 25789 29880 25823
rect 29828 25780 29880 25789
rect 33600 25823 33652 25832
rect 33600 25789 33609 25823
rect 33609 25789 33643 25823
rect 33643 25789 33652 25823
rect 33600 25780 33652 25789
rect 43168 25780 43220 25832
rect 42892 25712 42944 25764
rect 13820 25644 13872 25696
rect 14004 25644 14056 25696
rect 17316 25687 17368 25696
rect 17316 25653 17325 25687
rect 17325 25653 17359 25687
rect 17359 25653 17368 25687
rect 17316 25644 17368 25653
rect 20996 25644 21048 25696
rect 21088 25644 21140 25696
rect 22284 25687 22336 25696
rect 22284 25653 22293 25687
rect 22293 25653 22327 25687
rect 22327 25653 22336 25687
rect 22284 25644 22336 25653
rect 24860 25644 24912 25696
rect 25044 25687 25096 25696
rect 25044 25653 25053 25687
rect 25053 25653 25087 25687
rect 25087 25653 25096 25687
rect 25044 25644 25096 25653
rect 31576 25644 31628 25696
rect 31760 25687 31812 25696
rect 31760 25653 31769 25687
rect 31769 25653 31803 25687
rect 31803 25653 31812 25687
rect 31760 25644 31812 25653
rect 33232 25687 33284 25696
rect 33232 25653 33241 25687
rect 33241 25653 33275 25687
rect 33275 25653 33284 25687
rect 33232 25644 33284 25653
rect 33416 25687 33468 25696
rect 33416 25653 33425 25687
rect 33425 25653 33459 25687
rect 33459 25653 33468 25687
rect 33416 25644 33468 25653
rect 40316 25687 40368 25696
rect 40316 25653 40325 25687
rect 40325 25653 40359 25687
rect 40359 25653 40368 25687
rect 40316 25644 40368 25653
rect 58072 25644 58124 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 13544 25440 13596 25492
rect 22192 25483 22244 25492
rect 22192 25449 22201 25483
rect 22201 25449 22235 25483
rect 22235 25449 22244 25483
rect 22192 25440 22244 25449
rect 33232 25483 33284 25492
rect 33232 25449 33241 25483
rect 33241 25449 33275 25483
rect 33275 25449 33284 25483
rect 33232 25440 33284 25449
rect 44180 25440 44232 25492
rect 13452 25415 13504 25424
rect 13452 25381 13461 25415
rect 13461 25381 13495 25415
rect 13495 25381 13504 25415
rect 13452 25372 13504 25381
rect 20628 25304 20680 25356
rect 33140 25347 33192 25356
rect 33140 25313 33149 25347
rect 33149 25313 33183 25347
rect 33183 25313 33192 25347
rect 33140 25304 33192 25313
rect 14004 25236 14056 25288
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17316 25279 17368 25288
rect 17316 25245 17350 25279
rect 17350 25245 17368 25279
rect 17316 25236 17368 25245
rect 20352 25279 20404 25288
rect 20352 25245 20361 25279
rect 20361 25245 20395 25279
rect 20395 25245 20404 25279
rect 20352 25236 20404 25245
rect 21088 25279 21140 25288
rect 21088 25245 21122 25279
rect 21122 25245 21140 25279
rect 21088 25236 21140 25245
rect 24860 25236 24912 25288
rect 30656 25279 30708 25288
rect 30656 25245 30665 25279
rect 30665 25245 30699 25279
rect 30699 25245 30708 25279
rect 30656 25236 30708 25245
rect 31576 25236 31628 25288
rect 33968 25279 34020 25288
rect 13912 25168 13964 25220
rect 33968 25245 33977 25279
rect 33977 25245 34011 25279
rect 34011 25245 34020 25279
rect 33968 25236 34020 25245
rect 36268 25279 36320 25288
rect 36268 25245 36277 25279
rect 36277 25245 36311 25279
rect 36311 25245 36320 25279
rect 36268 25236 36320 25245
rect 36360 25236 36412 25288
rect 38568 25279 38620 25288
rect 38568 25245 38577 25279
rect 38577 25245 38611 25279
rect 38611 25245 38620 25279
rect 38568 25236 38620 25245
rect 40040 25279 40092 25288
rect 34704 25168 34756 25220
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 40316 25279 40368 25288
rect 40316 25245 40350 25279
rect 40350 25245 40368 25279
rect 40316 25236 40368 25245
rect 42708 25279 42760 25288
rect 42708 25245 42717 25279
rect 42717 25245 42751 25279
rect 42751 25245 42760 25279
rect 42708 25236 42760 25245
rect 40224 25168 40276 25220
rect 43812 25168 43864 25220
rect 14556 25100 14608 25152
rect 18880 25100 18932 25152
rect 33876 25100 33928 25152
rect 41696 25100 41748 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 13452 24896 13504 24948
rect 14004 24828 14056 24880
rect 14556 24939 14608 24948
rect 14556 24905 14581 24939
rect 14581 24905 14608 24939
rect 14556 24896 14608 24905
rect 22008 24896 22060 24948
rect 42064 24896 42116 24948
rect 42892 24896 42944 24948
rect 43812 24939 43864 24948
rect 13176 24760 13228 24812
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 13912 24760 13964 24812
rect 15844 24828 15896 24880
rect 17040 24828 17092 24880
rect 20628 24828 20680 24880
rect 31760 24828 31812 24880
rect 36084 24828 36136 24880
rect 38568 24871 38620 24880
rect 38568 24837 38602 24871
rect 38602 24837 38620 24871
rect 38568 24828 38620 24837
rect 40040 24828 40092 24880
rect 20352 24803 20404 24812
rect 20352 24769 20386 24803
rect 20386 24769 20404 24803
rect 20352 24760 20404 24769
rect 23112 24803 23164 24812
rect 23112 24769 23121 24803
rect 23121 24769 23155 24803
rect 23155 24769 23164 24803
rect 23112 24760 23164 24769
rect 29828 24760 29880 24812
rect 36268 24760 36320 24812
rect 36912 24760 36964 24812
rect 38108 24760 38160 24812
rect 41420 24828 41472 24880
rect 40224 24760 40276 24812
rect 42984 24828 43036 24880
rect 43444 24828 43496 24880
rect 43352 24803 43404 24812
rect 43352 24769 43361 24803
rect 43361 24769 43395 24803
rect 43395 24769 43404 24803
rect 43352 24760 43404 24769
rect 43812 24905 43821 24939
rect 43821 24905 43855 24939
rect 43855 24905 43864 24939
rect 43812 24896 43864 24905
rect 44180 24760 44232 24812
rect 24584 24624 24636 24676
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13360 24556 13412 24608
rect 15200 24556 15252 24608
rect 15384 24599 15436 24608
rect 15384 24565 15393 24599
rect 15393 24565 15427 24599
rect 15427 24565 15436 24599
rect 15384 24556 15436 24565
rect 17132 24599 17184 24608
rect 17132 24565 17141 24599
rect 17141 24565 17175 24599
rect 17175 24565 17184 24599
rect 17132 24556 17184 24565
rect 19156 24556 19208 24608
rect 29644 24599 29696 24608
rect 29644 24565 29653 24599
rect 29653 24565 29687 24599
rect 29687 24565 29696 24599
rect 29644 24556 29696 24565
rect 29920 24556 29972 24608
rect 31852 24556 31904 24608
rect 34520 24556 34572 24608
rect 34796 24599 34848 24608
rect 34796 24565 34805 24599
rect 34805 24565 34839 24599
rect 34839 24565 34848 24599
rect 34796 24556 34848 24565
rect 38200 24692 38252 24744
rect 37832 24667 37884 24676
rect 37832 24633 37841 24667
rect 37841 24633 37875 24667
rect 37875 24633 37884 24667
rect 37832 24624 37884 24633
rect 44364 24624 44416 24676
rect 35900 24556 35952 24608
rect 40868 24556 40920 24608
rect 41604 24556 41656 24608
rect 43168 24599 43220 24608
rect 43168 24565 43177 24599
rect 43177 24565 43211 24599
rect 43211 24565 43220 24599
rect 43168 24556 43220 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 22100 24352 22152 24361
rect 33140 24352 33192 24404
rect 41420 24352 41472 24404
rect 42708 24352 42760 24404
rect 13452 24284 13504 24336
rect 34704 24284 34756 24336
rect 17040 24216 17092 24268
rect 24584 24259 24636 24268
rect 12072 24148 12124 24200
rect 13544 24148 13596 24200
rect 12256 24080 12308 24132
rect 13820 24148 13872 24200
rect 16028 24191 16080 24200
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 17132 24148 17184 24200
rect 24584 24225 24593 24259
rect 24593 24225 24627 24259
rect 24627 24225 24636 24259
rect 24584 24216 24636 24225
rect 29920 24259 29972 24268
rect 29920 24225 29929 24259
rect 29929 24225 29963 24259
rect 29963 24225 29972 24259
rect 29920 24216 29972 24225
rect 31852 24259 31904 24268
rect 31852 24225 31861 24259
rect 31861 24225 31895 24259
rect 31895 24225 31904 24259
rect 31852 24216 31904 24225
rect 34796 24216 34848 24268
rect 38108 24216 38160 24268
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 24032 24191 24084 24200
rect 23020 24148 23072 24157
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29644 24148 29696 24200
rect 31668 24148 31720 24200
rect 32956 24191 33008 24200
rect 32956 24157 32965 24191
rect 32965 24157 32999 24191
rect 32999 24157 33008 24191
rect 32956 24148 33008 24157
rect 33968 24148 34020 24200
rect 34612 24148 34664 24200
rect 13912 24080 13964 24132
rect 15384 24080 15436 24132
rect 16212 24080 16264 24132
rect 20996 24123 21048 24132
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 13268 24055 13320 24064
rect 13268 24021 13277 24055
rect 13277 24021 13311 24055
rect 13311 24021 13320 24055
rect 13268 24012 13320 24021
rect 14004 24012 14056 24064
rect 14464 24012 14516 24064
rect 14648 24055 14700 24064
rect 14648 24021 14657 24055
rect 14657 24021 14691 24055
rect 14691 24021 14700 24055
rect 14648 24012 14700 24021
rect 18696 24055 18748 24064
rect 18696 24021 18705 24055
rect 18705 24021 18739 24055
rect 18739 24021 18748 24055
rect 20996 24089 21030 24123
rect 21030 24089 21048 24123
rect 20996 24080 21048 24089
rect 24676 24080 24728 24132
rect 18696 24012 18748 24021
rect 23296 24012 23348 24064
rect 31852 24080 31904 24132
rect 36084 24123 36136 24132
rect 36084 24089 36093 24123
rect 36093 24089 36127 24123
rect 36127 24089 36136 24123
rect 36084 24080 36136 24089
rect 25780 24012 25832 24064
rect 41144 24012 41196 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 19340 23851 19392 23860
rect 12256 23740 12308 23792
rect 16212 23740 16264 23792
rect 16856 23740 16908 23792
rect 19340 23817 19349 23851
rect 19349 23817 19383 23851
rect 19383 23817 19392 23851
rect 19340 23808 19392 23817
rect 24952 23808 25004 23860
rect 31668 23851 31720 23860
rect 31668 23817 31677 23851
rect 31677 23817 31711 23851
rect 31711 23817 31720 23851
rect 31668 23808 31720 23817
rect 34612 23851 34664 23860
rect 34612 23817 34621 23851
rect 34621 23817 34655 23851
rect 34655 23817 34664 23851
rect 34612 23808 34664 23817
rect 36912 23851 36964 23860
rect 36912 23817 36921 23851
rect 36921 23817 36955 23851
rect 36955 23817 36964 23851
rect 36912 23808 36964 23817
rect 38108 23808 38160 23860
rect 38200 23808 38252 23860
rect 42984 23851 43036 23860
rect 42984 23817 42993 23851
rect 42993 23817 43027 23851
rect 43027 23817 43036 23851
rect 42984 23808 43036 23817
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 15200 23672 15252 23724
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 16028 23672 16080 23724
rect 19156 23715 19208 23724
rect 19156 23681 19165 23715
rect 19165 23681 19199 23715
rect 19199 23681 19208 23715
rect 19156 23672 19208 23681
rect 23296 23715 23348 23724
rect 23296 23681 23305 23715
rect 23305 23681 23339 23715
rect 23339 23681 23348 23715
rect 23296 23672 23348 23681
rect 24584 23740 24636 23792
rect 30656 23740 30708 23792
rect 24032 23715 24084 23724
rect 24032 23681 24066 23715
rect 24066 23681 24084 23715
rect 24032 23672 24084 23681
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 25872 23715 25924 23724
rect 25872 23681 25881 23715
rect 25881 23681 25915 23715
rect 25915 23681 25924 23715
rect 25872 23672 25924 23681
rect 29828 23715 29880 23724
rect 29828 23681 29837 23715
rect 29837 23681 29871 23715
rect 29871 23681 29880 23715
rect 29828 23672 29880 23681
rect 29920 23672 29972 23724
rect 32956 23672 33008 23724
rect 33508 23715 33560 23724
rect 33508 23681 33542 23715
rect 33542 23681 33560 23715
rect 35900 23740 35952 23792
rect 33508 23672 33560 23681
rect 36360 23672 36412 23724
rect 37924 23672 37976 23724
rect 40040 23715 40092 23724
rect 40040 23681 40049 23715
rect 40049 23681 40083 23715
rect 40083 23681 40092 23715
rect 40040 23672 40092 23681
rect 40316 23715 40368 23724
rect 40316 23681 40350 23715
rect 40350 23681 40368 23715
rect 42616 23715 42668 23724
rect 40316 23672 40368 23681
rect 42616 23681 42625 23715
rect 42625 23681 42659 23715
rect 42659 23681 42668 23715
rect 42616 23672 42668 23681
rect 43628 23672 43680 23724
rect 18696 23604 18748 23656
rect 25780 23647 25832 23656
rect 25780 23613 25789 23647
rect 25789 23613 25823 23647
rect 25823 23613 25832 23647
rect 25780 23604 25832 23613
rect 11060 23536 11112 23588
rect 14004 23468 14056 23520
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 18880 23511 18932 23520
rect 18880 23477 18889 23511
rect 18889 23477 18923 23511
rect 18923 23477 18932 23511
rect 18880 23468 18932 23477
rect 41512 23468 41564 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12256 23264 12308 23316
rect 13820 23128 13872 23180
rect 15660 23264 15712 23316
rect 16212 23307 16264 23316
rect 16212 23273 16221 23307
rect 16221 23273 16255 23307
rect 16255 23273 16264 23307
rect 16212 23264 16264 23273
rect 25596 23264 25648 23316
rect 25872 23264 25924 23316
rect 31852 23264 31904 23316
rect 33508 23264 33560 23316
rect 37924 23264 37976 23316
rect 40316 23264 40368 23316
rect 41512 23264 41564 23316
rect 15476 23196 15528 23248
rect 42616 23196 42668 23248
rect 14648 23171 14700 23180
rect 14648 23137 14657 23171
rect 14657 23137 14691 23171
rect 14691 23137 14700 23171
rect 24584 23171 24636 23180
rect 14648 23128 14700 23137
rect 12348 23060 12400 23112
rect 12072 22992 12124 23044
rect 14556 23103 14608 23112
rect 14556 23069 14565 23103
rect 14565 23069 14599 23103
rect 14599 23069 14608 23103
rect 24584 23137 24593 23171
rect 24593 23137 24627 23171
rect 24627 23137 24636 23171
rect 24584 23128 24636 23137
rect 41604 23128 41656 23180
rect 14556 23060 14608 23069
rect 24860 23103 24912 23112
rect 24860 23069 24894 23103
rect 24894 23069 24912 23103
rect 24860 23060 24912 23069
rect 28908 23060 28960 23112
rect 40868 23103 40920 23112
rect 40868 23069 40877 23103
rect 40877 23069 40911 23103
rect 40911 23069 40920 23103
rect 40868 23060 40920 23069
rect 41696 23060 41748 23112
rect 15200 22992 15252 23044
rect 23020 22992 23072 23044
rect 29184 22992 29236 23044
rect 2872 22967 2924 22976
rect 2872 22933 2881 22967
rect 2881 22933 2915 22967
rect 2915 22933 2924 22967
rect 2872 22924 2924 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 12072 22720 12124 22772
rect 13820 22720 13872 22772
rect 2872 22652 2924 22704
rect 12992 22652 13044 22704
rect 13820 22584 13872 22636
rect 14004 22627 14056 22636
rect 14004 22593 14013 22627
rect 14013 22593 14047 22627
rect 14047 22593 14056 22627
rect 14004 22584 14056 22593
rect 37556 22584 37608 22636
rect 38200 22584 38252 22636
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 16672 22380 16724 22432
rect 37924 22423 37976 22432
rect 37924 22389 37933 22423
rect 37933 22389 37967 22423
rect 37967 22389 37976 22423
rect 37924 22380 37976 22389
rect 41604 22423 41656 22432
rect 41604 22389 41613 22423
rect 41613 22389 41647 22423
rect 41647 22389 41656 22423
rect 41604 22380 41656 22389
rect 42616 22423 42668 22432
rect 42616 22389 42625 22423
rect 42625 22389 42659 22423
rect 42659 22389 42668 22423
rect 42616 22380 42668 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1768 22219 1820 22228
rect 1768 22185 1777 22219
rect 1777 22185 1811 22219
rect 1811 22185 1820 22219
rect 1768 22176 1820 22185
rect 13360 22219 13412 22228
rect 13360 22185 13369 22219
rect 13369 22185 13403 22219
rect 13403 22185 13412 22219
rect 13360 22176 13412 22185
rect 2872 22151 2924 22160
rect 2872 22117 2881 22151
rect 2881 22117 2915 22151
rect 2915 22117 2924 22151
rect 2872 22108 2924 22117
rect 32864 22151 32916 22160
rect 32864 22117 32873 22151
rect 32873 22117 32907 22151
rect 32907 22117 32916 22151
rect 32864 22108 32916 22117
rect 42892 22108 42944 22160
rect 35900 22040 35952 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 13268 21972 13320 22024
rect 17040 21972 17092 22024
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 33876 22015 33928 22024
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 34060 22015 34112 22024
rect 34060 21981 34069 22015
rect 34069 21981 34103 22015
rect 34103 21981 34112 22015
rect 34060 21972 34112 21981
rect 38844 22015 38896 22024
rect 38844 21981 38853 22015
rect 38853 21981 38887 22015
rect 38887 21981 38896 22015
rect 38844 21972 38896 21981
rect 39028 22015 39080 22024
rect 39028 21981 39037 22015
rect 39037 21981 39071 22015
rect 39071 21981 39080 22015
rect 39028 21972 39080 21981
rect 41420 21972 41472 22024
rect 41604 22015 41656 22024
rect 41604 21981 41638 22015
rect 41638 21981 41656 22015
rect 41604 21972 41656 21981
rect 43352 22015 43404 22024
rect 43352 21981 43361 22015
rect 43361 21981 43395 22015
rect 43395 21981 43404 22015
rect 43352 21972 43404 21981
rect 43720 21972 43772 22024
rect 13452 21904 13504 21956
rect 36636 21904 36688 21956
rect 38200 21947 38252 21956
rect 4620 21836 4672 21888
rect 13176 21879 13228 21888
rect 13176 21845 13185 21879
rect 13185 21845 13219 21879
rect 13219 21845 13228 21879
rect 13176 21836 13228 21845
rect 14372 21879 14424 21888
rect 14372 21845 14381 21879
rect 14381 21845 14415 21879
rect 14415 21845 14424 21879
rect 14372 21836 14424 21845
rect 37372 21836 37424 21888
rect 37556 21879 37608 21888
rect 37556 21845 37565 21879
rect 37565 21845 37599 21879
rect 37599 21845 37608 21879
rect 38200 21913 38209 21947
rect 38209 21913 38243 21947
rect 38243 21913 38252 21947
rect 38200 21904 38252 21913
rect 41880 21904 41932 21956
rect 38384 21879 38436 21888
rect 37556 21836 37608 21845
rect 38384 21845 38393 21879
rect 38393 21845 38427 21879
rect 38427 21845 38436 21879
rect 38384 21836 38436 21845
rect 39212 21879 39264 21888
rect 39212 21845 39221 21879
rect 39221 21845 39255 21879
rect 39255 21845 39264 21879
rect 39212 21836 39264 21845
rect 43628 21879 43680 21888
rect 43628 21845 43637 21879
rect 43637 21845 43671 21879
rect 43671 21845 43680 21879
rect 43628 21836 43680 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2596 21632 2648 21684
rect 2964 21632 3016 21684
rect 38200 21632 38252 21684
rect 43352 21632 43404 21684
rect 17592 21564 17644 21616
rect 20352 21607 20404 21616
rect 20352 21573 20386 21607
rect 20386 21573 20404 21607
rect 20352 21564 20404 21573
rect 4620 21496 4672 21548
rect 14004 21496 14056 21548
rect 14372 21496 14424 21548
rect 14832 21496 14884 21548
rect 16948 21496 17000 21548
rect 18052 21496 18104 21548
rect 30748 21539 30800 21548
rect 18788 21471 18840 21480
rect 18788 21437 18797 21471
rect 18797 21437 18831 21471
rect 18831 21437 18840 21471
rect 18788 21428 18840 21437
rect 30748 21505 30757 21539
rect 30757 21505 30791 21539
rect 30791 21505 30800 21539
rect 30748 21496 30800 21505
rect 31024 21539 31076 21548
rect 31024 21505 31033 21539
rect 31033 21505 31067 21539
rect 31067 21505 31076 21539
rect 31024 21496 31076 21505
rect 35900 21564 35952 21616
rect 37556 21564 37608 21616
rect 34152 21496 34204 21548
rect 35440 21539 35492 21548
rect 35440 21505 35449 21539
rect 35449 21505 35483 21539
rect 35483 21505 35492 21539
rect 35440 21496 35492 21505
rect 35532 21496 35584 21548
rect 37740 21539 37792 21548
rect 37740 21505 37774 21539
rect 37774 21505 37792 21539
rect 37740 21496 37792 21505
rect 39396 21496 39448 21548
rect 41420 21496 41472 21548
rect 42340 21496 42392 21548
rect 42892 21539 42944 21548
rect 42892 21505 42926 21539
rect 42926 21505 42944 21539
rect 42892 21496 42944 21505
rect 20076 21471 20128 21480
rect 20076 21437 20085 21471
rect 20085 21437 20119 21471
rect 20119 21437 20128 21471
rect 20076 21428 20128 21437
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 30840 21471 30892 21480
rect 30840 21437 30849 21471
rect 30849 21437 30883 21471
rect 30883 21437 30892 21471
rect 30840 21428 30892 21437
rect 36268 21428 36320 21480
rect 33232 21360 33284 21412
rect 2320 21292 2372 21344
rect 5540 21292 5592 21344
rect 16580 21292 16632 21344
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 19064 21292 19116 21344
rect 21456 21335 21508 21344
rect 21456 21301 21465 21335
rect 21465 21301 21499 21335
rect 21499 21301 21508 21335
rect 21456 21292 21508 21301
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 31760 21335 31812 21344
rect 31760 21301 31769 21335
rect 31769 21301 31803 21335
rect 31803 21301 31812 21335
rect 31760 21292 31812 21301
rect 32588 21292 32640 21344
rect 34520 21292 34572 21344
rect 37372 21360 37424 21412
rect 36820 21292 36872 21344
rect 39120 21292 39172 21344
rect 40776 21292 40828 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3976 21131 4028 21140
rect 3976 21097 3985 21131
rect 3985 21097 4019 21131
rect 4019 21097 4028 21131
rect 3976 21088 4028 21097
rect 18696 21088 18748 21140
rect 21456 21088 21508 21140
rect 30840 21088 30892 21140
rect 34152 21131 34204 21140
rect 34152 21097 34161 21131
rect 34161 21097 34195 21131
rect 34195 21097 34204 21131
rect 34152 21088 34204 21097
rect 36268 21131 36320 21140
rect 36268 21097 36277 21131
rect 36277 21097 36311 21131
rect 36311 21097 36320 21131
rect 36268 21088 36320 21097
rect 38384 21088 38436 21140
rect 39028 21088 39080 21140
rect 39396 21131 39448 21140
rect 39396 21097 39405 21131
rect 39405 21097 39439 21131
rect 39439 21097 39448 21131
rect 39396 21088 39448 21097
rect 37372 21020 37424 21072
rect 38844 21020 38896 21072
rect 2596 20884 2648 20936
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 13636 20884 13688 20936
rect 13912 20884 13964 20936
rect 16764 20884 16816 20936
rect 19984 20884 20036 20936
rect 20076 20884 20128 20936
rect 20996 20884 21048 20936
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 27896 20884 27948 20936
rect 28908 20884 28960 20936
rect 29920 20884 29972 20936
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 32588 20927 32640 20936
rect 32588 20893 32622 20927
rect 32622 20893 32640 20927
rect 32588 20884 32640 20893
rect 35900 20884 35952 20936
rect 36728 20927 36780 20936
rect 36728 20893 36737 20927
rect 36737 20893 36771 20927
rect 36771 20893 36780 20927
rect 36728 20884 36780 20893
rect 2136 20816 2188 20868
rect 3424 20816 3476 20868
rect 17040 20816 17092 20868
rect 22100 20859 22152 20868
rect 22100 20825 22109 20859
rect 22109 20825 22143 20859
rect 22143 20825 22152 20859
rect 22100 20816 22152 20825
rect 4712 20748 4764 20800
rect 22560 20791 22612 20800
rect 22560 20757 22569 20791
rect 22569 20757 22603 20791
rect 22603 20757 22612 20791
rect 22560 20748 22612 20757
rect 31760 20816 31812 20868
rect 35348 20816 35400 20868
rect 37924 20952 37976 21004
rect 39120 20952 39172 21004
rect 41420 21088 41472 21140
rect 41880 21131 41932 21140
rect 41880 21097 41889 21131
rect 41889 21097 41923 21131
rect 41923 21097 41932 21131
rect 41880 21088 41932 21097
rect 43720 21131 43772 21140
rect 43720 21097 43729 21131
rect 43729 21097 43763 21131
rect 43763 21097 43772 21131
rect 43720 21088 43772 21097
rect 42340 20995 42392 21004
rect 42340 20961 42349 20995
rect 42349 20961 42383 20995
rect 42383 20961 42392 20995
rect 42340 20952 42392 20961
rect 39212 20927 39264 20936
rect 39212 20893 39221 20927
rect 39221 20893 39255 20927
rect 39255 20893 39264 20927
rect 39212 20884 39264 20893
rect 40776 20927 40828 20936
rect 40776 20893 40810 20927
rect 40810 20893 40828 20927
rect 40776 20884 40828 20893
rect 42616 20927 42668 20936
rect 42616 20893 42650 20927
rect 42650 20893 42668 20927
rect 42616 20884 42668 20893
rect 30472 20748 30524 20800
rect 33508 20748 33560 20800
rect 37924 20748 37976 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 3976 20587 4028 20596
rect 3976 20553 3985 20587
rect 3985 20553 4019 20587
rect 4019 20553 4028 20587
rect 3976 20544 4028 20553
rect 4252 20544 4304 20596
rect 2872 20519 2924 20528
rect 2872 20485 2906 20519
rect 2906 20485 2924 20519
rect 2872 20476 2924 20485
rect 5540 20519 5592 20528
rect 5540 20485 5558 20519
rect 5558 20485 5592 20519
rect 5540 20476 5592 20485
rect 2136 20451 2188 20460
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 2136 20408 2188 20417
rect 2596 20451 2648 20460
rect 2596 20417 2605 20451
rect 2605 20417 2639 20451
rect 2639 20417 2648 20451
rect 2596 20408 2648 20417
rect 13820 20476 13872 20528
rect 16580 20476 16632 20528
rect 22376 20544 22428 20596
rect 30748 20544 30800 20596
rect 31024 20544 31076 20596
rect 32864 20519 32916 20528
rect 13912 20408 13964 20460
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15660 20408 15712 20460
rect 16948 20408 17000 20460
rect 19984 20408 20036 20460
rect 32864 20485 32898 20519
rect 32898 20485 32916 20519
rect 32864 20476 32916 20485
rect 35440 20544 35492 20596
rect 36636 20587 36688 20596
rect 36636 20553 36645 20587
rect 36645 20553 36679 20587
rect 36679 20553 36688 20587
rect 36636 20544 36688 20553
rect 37740 20587 37792 20596
rect 37740 20553 37749 20587
rect 37749 20553 37783 20587
rect 37783 20553 37792 20587
rect 37740 20544 37792 20553
rect 35532 20476 35584 20528
rect 36728 20476 36780 20528
rect 39120 20519 39172 20528
rect 39120 20485 39129 20519
rect 39129 20485 39163 20519
rect 39163 20485 39172 20519
rect 39120 20476 39172 20485
rect 22560 20408 22612 20460
rect 27896 20408 27948 20460
rect 28264 20451 28316 20460
rect 28264 20417 28298 20451
rect 28298 20417 28316 20451
rect 29920 20451 29972 20460
rect 28264 20408 28316 20417
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 30012 20408 30064 20460
rect 35900 20408 35952 20460
rect 36820 20451 36872 20460
rect 36820 20417 36829 20451
rect 36829 20417 36863 20451
rect 36863 20417 36872 20451
rect 36820 20408 36872 20417
rect 37924 20451 37976 20460
rect 37924 20417 37933 20451
rect 37933 20417 37967 20451
rect 37967 20417 37976 20451
rect 37924 20408 37976 20417
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 14740 20340 14792 20392
rect 18972 20383 19024 20392
rect 18972 20349 18981 20383
rect 18981 20349 19015 20383
rect 19015 20349 19024 20383
rect 18972 20340 19024 20349
rect 20076 20383 20128 20392
rect 20076 20349 20085 20383
rect 20085 20349 20119 20383
rect 20119 20349 20128 20383
rect 20076 20340 20128 20349
rect 32312 20340 32364 20392
rect 18788 20272 18840 20324
rect 38844 20272 38896 20324
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19340 20204 19392 20256
rect 40132 20204 40184 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3424 20043 3476 20052
rect 3424 20009 3433 20043
rect 3433 20009 3467 20043
rect 3467 20009 3476 20043
rect 3424 20000 3476 20009
rect 15200 20000 15252 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 18052 20000 18104 20052
rect 22100 20000 22152 20052
rect 28264 20043 28316 20052
rect 28264 20009 28273 20043
rect 28273 20009 28307 20043
rect 28307 20009 28316 20043
rect 28264 20000 28316 20009
rect 30012 20043 30064 20052
rect 30012 20009 30021 20043
rect 30021 20009 30055 20043
rect 30055 20009 30064 20043
rect 30012 20000 30064 20009
rect 30472 20043 30524 20052
rect 30472 20009 30481 20043
rect 30481 20009 30515 20043
rect 30515 20009 30524 20043
rect 30472 20000 30524 20009
rect 33508 20043 33560 20052
rect 33508 20009 33517 20043
rect 33517 20009 33551 20043
rect 33551 20009 33560 20043
rect 33508 20000 33560 20009
rect 34060 20000 34112 20052
rect 35348 20000 35400 20052
rect 13820 19864 13872 19916
rect 34520 19864 34572 19916
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 2320 19839 2372 19848
rect 2320 19805 2354 19839
rect 2354 19805 2372 19839
rect 2320 19796 2372 19805
rect 20076 19796 20128 19848
rect 22008 19796 22060 19848
rect 32128 19839 32180 19848
rect 32128 19805 32137 19839
rect 32137 19805 32171 19839
rect 32171 19805 32180 19839
rect 32128 19796 32180 19805
rect 33232 19839 33284 19848
rect 33232 19805 33241 19839
rect 33241 19805 33275 19839
rect 33275 19805 33284 19839
rect 33232 19796 33284 19805
rect 33692 19796 33744 19848
rect 12716 19728 12768 19780
rect 14556 19771 14608 19780
rect 14556 19737 14590 19771
rect 14590 19737 14608 19771
rect 14556 19728 14608 19737
rect 16672 19728 16724 19780
rect 16948 19728 17000 19780
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 14740 19499 14792 19508
rect 14740 19465 14749 19499
rect 14749 19465 14783 19499
rect 14783 19465 14792 19499
rect 14740 19456 14792 19465
rect 33692 19499 33744 19508
rect 33692 19465 33701 19499
rect 33701 19465 33735 19499
rect 33735 19465 33744 19499
rect 33692 19456 33744 19465
rect 5816 19320 5868 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 13820 19388 13872 19440
rect 32128 19388 32180 19440
rect 13636 19363 13688 19372
rect 13636 19329 13670 19363
rect 13670 19329 13688 19363
rect 13636 19320 13688 19329
rect 14832 19320 14884 19372
rect 17960 19320 18012 19372
rect 18420 19320 18472 19372
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 2320 19116 2372 19168
rect 7932 19159 7984 19168
rect 7932 19125 7941 19159
rect 7941 19125 7975 19159
rect 7975 19125 7984 19159
rect 7932 19116 7984 19125
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 20076 19116 20128 19168
rect 37832 19159 37884 19168
rect 37832 19125 37841 19159
rect 37841 19125 37875 19159
rect 37875 19125 37884 19159
rect 37832 19116 37884 19125
rect 40960 19159 41012 19168
rect 40960 19125 40969 19159
rect 40969 19125 41003 19159
rect 41003 19125 41012 19159
rect 40960 19116 41012 19125
rect 42800 19116 42852 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7932 18912 7984 18964
rect 14556 18912 14608 18964
rect 2044 18819 2096 18828
rect 2044 18785 2053 18819
rect 2053 18785 2087 18819
rect 2087 18785 2096 18819
rect 2044 18776 2096 18785
rect 3884 18776 3936 18828
rect 2320 18751 2372 18760
rect 2320 18717 2354 18751
rect 2354 18717 2372 18751
rect 2320 18708 2372 18717
rect 4160 18708 4212 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 7012 18708 7064 18760
rect 7932 18708 7984 18760
rect 16856 18708 16908 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 20812 18708 20864 18760
rect 21088 18751 21140 18760
rect 21088 18717 21097 18751
rect 21097 18717 21131 18751
rect 21131 18717 21140 18751
rect 21088 18708 21140 18717
rect 37372 18708 37424 18760
rect 37464 18708 37516 18760
rect 40776 18708 40828 18760
rect 40960 18751 41012 18760
rect 40960 18717 40994 18751
rect 40994 18717 41012 18751
rect 40960 18708 41012 18717
rect 44456 18751 44508 18760
rect 44456 18717 44465 18751
rect 44465 18717 44499 18751
rect 44499 18717 44508 18751
rect 44456 18708 44508 18717
rect 3516 18640 3568 18692
rect 7380 18683 7432 18692
rect 7380 18649 7389 18683
rect 7389 18649 7423 18683
rect 7423 18649 7432 18683
rect 7380 18640 7432 18649
rect 16304 18640 16356 18692
rect 37832 18683 37884 18692
rect 37832 18649 37866 18683
rect 37866 18649 37884 18683
rect 37832 18640 37884 18649
rect 4436 18615 4488 18624
rect 4436 18581 4445 18615
rect 4445 18581 4479 18615
rect 4479 18581 4488 18615
rect 4436 18572 4488 18581
rect 4804 18572 4856 18624
rect 18788 18572 18840 18624
rect 20996 18615 21048 18624
rect 20996 18581 21005 18615
rect 21005 18581 21039 18615
rect 21039 18581 21048 18615
rect 20996 18572 21048 18581
rect 38936 18615 38988 18624
rect 38936 18581 38945 18615
rect 38945 18581 38979 18615
rect 38979 18581 38988 18615
rect 38936 18572 38988 18581
rect 42616 18572 42668 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 7932 18411 7984 18420
rect 7932 18377 7941 18411
rect 7941 18377 7975 18411
rect 7975 18377 7984 18411
rect 7932 18368 7984 18377
rect 18972 18368 19024 18420
rect 2044 18232 2096 18284
rect 2228 18232 2280 18284
rect 4712 18300 4764 18352
rect 7104 18300 7156 18352
rect 18788 18343 18840 18352
rect 18788 18309 18797 18343
rect 18797 18309 18831 18343
rect 18831 18309 18840 18343
rect 18788 18300 18840 18309
rect 44456 18343 44508 18352
rect 44456 18309 44490 18343
rect 44490 18309 44508 18343
rect 44456 18300 44508 18309
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 17040 18232 17092 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 20720 18232 20772 18284
rect 21456 18232 21508 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 22928 18232 22980 18284
rect 40776 18232 40828 18284
rect 40960 18275 41012 18284
rect 40960 18241 40994 18275
rect 40994 18241 41012 18275
rect 40960 18232 41012 18241
rect 41972 18232 42024 18284
rect 43996 18232 44048 18284
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 37464 18207 37516 18216
rect 37464 18173 37473 18207
rect 37473 18173 37507 18207
rect 37507 18173 37516 18207
rect 37464 18164 37516 18173
rect 3976 18071 4028 18080
rect 3976 18037 3985 18071
rect 3985 18037 4019 18071
rect 4019 18037 4028 18071
rect 3976 18028 4028 18037
rect 4436 18028 4488 18080
rect 5080 18028 5132 18080
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 22192 18028 22244 18080
rect 36912 18071 36964 18080
rect 36912 18037 36921 18071
rect 36921 18037 36955 18071
rect 36955 18037 36964 18071
rect 36912 18028 36964 18037
rect 38844 18071 38896 18080
rect 38844 18037 38853 18071
rect 38853 18037 38887 18071
rect 38887 18037 38896 18071
rect 38844 18028 38896 18037
rect 40316 18028 40368 18080
rect 42616 18071 42668 18080
rect 42616 18037 42625 18071
rect 42625 18037 42659 18071
rect 42659 18037 42668 18071
rect 42616 18028 42668 18037
rect 43352 18028 43404 18080
rect 44548 18028 44600 18080
rect 46296 18028 46348 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3884 17824 3936 17876
rect 7012 17824 7064 17876
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 19064 17824 19116 17876
rect 38752 17867 38804 17876
rect 38752 17833 38761 17867
rect 38761 17833 38795 17867
rect 38795 17833 38804 17867
rect 38752 17824 38804 17833
rect 43352 17867 43404 17876
rect 43352 17833 43361 17867
rect 43361 17833 43395 17867
rect 43395 17833 43404 17867
rect 43352 17824 43404 17833
rect 22928 17799 22980 17808
rect 22928 17765 22937 17799
rect 22937 17765 22971 17799
rect 22971 17765 22980 17799
rect 22928 17756 22980 17765
rect 2044 17731 2096 17740
rect 2044 17697 2053 17731
rect 2053 17697 2087 17731
rect 2087 17697 2096 17731
rect 2044 17688 2096 17697
rect 16948 17688 17000 17740
rect 38844 17731 38896 17740
rect 3976 17620 4028 17672
rect 4620 17620 4672 17672
rect 6552 17620 6604 17672
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 38844 17697 38853 17731
rect 38853 17697 38887 17731
rect 38887 17697 38896 17731
rect 38844 17688 38896 17697
rect 43444 17731 43496 17740
rect 43444 17697 43453 17731
rect 43453 17697 43487 17731
rect 43487 17697 43496 17731
rect 43444 17688 43496 17697
rect 37464 17620 37516 17672
rect 38936 17663 38988 17672
rect 38936 17629 38945 17663
rect 38945 17629 38979 17663
rect 38979 17629 38988 17663
rect 38936 17620 38988 17629
rect 43628 17663 43680 17672
rect 43628 17629 43637 17663
rect 43637 17629 43671 17663
rect 43671 17629 43680 17663
rect 43628 17620 43680 17629
rect 44640 17663 44692 17672
rect 44640 17629 44649 17663
rect 44649 17629 44683 17663
rect 44683 17629 44692 17663
rect 44640 17620 44692 17629
rect 45192 17663 45244 17672
rect 45192 17629 45201 17663
rect 45201 17629 45235 17663
rect 45235 17629 45244 17663
rect 45192 17620 45244 17629
rect 4620 17484 4672 17536
rect 7104 17552 7156 17604
rect 8392 17552 8444 17604
rect 18604 17552 18656 17604
rect 20076 17552 20128 17604
rect 21640 17552 21692 17604
rect 36912 17595 36964 17604
rect 36912 17561 36946 17595
rect 36946 17561 36964 17595
rect 36912 17552 36964 17561
rect 41144 17595 41196 17604
rect 20996 17484 21048 17536
rect 22100 17484 22152 17536
rect 41144 17561 41153 17595
rect 41153 17561 41187 17595
rect 41187 17561 41196 17595
rect 41144 17552 41196 17561
rect 42892 17595 42944 17604
rect 42892 17561 42901 17595
rect 42901 17561 42935 17595
rect 42935 17561 42944 17595
rect 42892 17552 42944 17561
rect 43904 17484 43956 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4160 17280 4212 17332
rect 18880 17280 18932 17332
rect 21088 17280 21140 17332
rect 22928 17280 22980 17332
rect 38752 17280 38804 17332
rect 41972 17280 42024 17332
rect 42800 17280 42852 17332
rect 2044 17144 2096 17196
rect 5632 17212 5684 17264
rect 14648 17255 14700 17264
rect 14648 17221 14682 17255
rect 14682 17221 14700 17255
rect 14648 17212 14700 17221
rect 17408 17212 17460 17264
rect 3976 17144 4028 17196
rect 4620 17187 4672 17196
rect 4620 17153 4629 17187
rect 4629 17153 4663 17187
rect 4663 17153 4672 17187
rect 4620 17144 4672 17153
rect 16948 17144 17000 17196
rect 22100 17212 22152 17264
rect 37372 17212 37424 17264
rect 43628 17280 43680 17332
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 40040 17144 40092 17196
rect 45192 17212 45244 17264
rect 40316 17144 40368 17196
rect 40776 17144 40828 17196
rect 2228 17076 2280 17128
rect 14280 17076 14332 17128
rect 21088 17119 21140 17128
rect 21088 17085 21097 17119
rect 21097 17085 21131 17119
rect 21131 17085 21140 17119
rect 21088 17076 21140 17085
rect 44548 17144 44600 17196
rect 45560 17144 45612 17196
rect 46572 17187 46624 17196
rect 46572 17153 46581 17187
rect 46581 17153 46615 17187
rect 46615 17153 46624 17187
rect 46572 17144 46624 17153
rect 7380 17008 7432 17060
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 16120 16940 16172 16992
rect 21088 16940 21140 16992
rect 21456 16940 21508 16992
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 43996 17051 44048 17060
rect 43996 17017 44005 17051
rect 44005 17017 44039 17051
rect 44039 17017 44048 17051
rect 43996 17008 44048 17017
rect 42800 16940 42852 16992
rect 46296 16983 46348 16992
rect 46296 16949 46305 16983
rect 46305 16949 46339 16983
rect 46339 16949 46348 16983
rect 46296 16940 46348 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3976 16779 4028 16788
rect 3976 16745 3985 16779
rect 3985 16745 4019 16779
rect 4019 16745 4028 16779
rect 3976 16736 4028 16745
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 21640 16736 21692 16788
rect 40960 16779 41012 16788
rect 40960 16745 40969 16779
rect 40969 16745 41003 16779
rect 41003 16745 41012 16779
rect 40960 16736 41012 16745
rect 46572 16779 46624 16788
rect 46572 16745 46581 16779
rect 46581 16745 46615 16779
rect 46615 16745 46624 16779
rect 46572 16736 46624 16745
rect 20812 16668 20864 16720
rect 14188 16600 14240 16652
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16212 16600 16264 16609
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16488 16532 16540 16584
rect 20812 16532 20864 16584
rect 21088 16600 21140 16652
rect 42800 16600 42852 16652
rect 44548 16600 44600 16652
rect 14096 16464 14148 16516
rect 22192 16532 22244 16584
rect 41144 16532 41196 16584
rect 44456 16575 44508 16584
rect 44456 16541 44465 16575
rect 44465 16541 44499 16575
rect 44499 16541 44508 16575
rect 44456 16532 44508 16541
rect 44640 16532 44692 16584
rect 22376 16464 22428 16516
rect 17776 16396 17828 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 16212 16192 16264 16244
rect 14188 16124 14240 16176
rect 20812 16192 20864 16244
rect 41144 16192 41196 16244
rect 45560 16192 45612 16244
rect 20260 16124 20312 16176
rect 44456 16124 44508 16176
rect 9128 16056 9180 16108
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 20076 16056 20128 16108
rect 14280 15988 14332 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 19984 15988 20036 16040
rect 20904 16056 20956 16108
rect 42800 16056 42852 16108
rect 43812 16056 43864 16108
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 20076 15852 20128 15904
rect 40316 15852 40368 15904
rect 40592 15895 40644 15904
rect 40592 15861 40601 15895
rect 40601 15861 40635 15895
rect 40635 15861 40644 15895
rect 40592 15852 40644 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8208 15648 8260 15700
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 20812 15648 20864 15700
rect 43444 15648 43496 15700
rect 19340 15512 19392 15564
rect 8944 15444 8996 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 16856 15444 16908 15496
rect 19248 15444 19300 15496
rect 22284 15512 22336 15564
rect 40040 15555 40092 15564
rect 40040 15521 40049 15555
rect 40049 15521 40083 15555
rect 40083 15521 40092 15555
rect 40040 15512 40092 15521
rect 41972 15555 42024 15564
rect 41972 15521 41981 15555
rect 41981 15521 42015 15555
rect 42015 15521 42024 15555
rect 41972 15512 42024 15521
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 8024 15419 8076 15428
rect 8024 15385 8033 15419
rect 8033 15385 8067 15419
rect 8067 15385 8076 15419
rect 8024 15376 8076 15385
rect 19340 15376 19392 15428
rect 19984 15376 20036 15428
rect 20904 15419 20956 15428
rect 20904 15385 20913 15419
rect 20913 15385 20947 15419
rect 20947 15385 20956 15419
rect 20904 15376 20956 15385
rect 22100 15376 22152 15428
rect 39580 15444 39632 15496
rect 40592 15444 40644 15496
rect 42156 15487 42208 15496
rect 42156 15453 42165 15487
rect 42165 15453 42199 15487
rect 42199 15453 42208 15487
rect 42156 15444 42208 15453
rect 43720 15487 43772 15496
rect 43720 15453 43729 15487
rect 43729 15453 43763 15487
rect 43763 15453 43772 15487
rect 43720 15444 43772 15453
rect 41880 15419 41932 15428
rect 41880 15385 41889 15419
rect 41889 15385 41923 15419
rect 41923 15385 41932 15419
rect 41880 15376 41932 15385
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 8944 15308 8996 15360
rect 9312 15308 9364 15360
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 22652 15351 22704 15360
rect 22652 15317 22661 15351
rect 22661 15317 22695 15351
rect 22695 15317 22704 15351
rect 22652 15308 22704 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 8944 15147 8996 15156
rect 8944 15113 8953 15147
rect 8953 15113 8987 15147
rect 8987 15113 8996 15147
rect 8944 15104 8996 15113
rect 4620 15036 4672 15088
rect 9312 15079 9364 15088
rect 9312 15045 9321 15079
rect 9321 15045 9355 15079
rect 9355 15045 9364 15079
rect 9312 15036 9364 15045
rect 11152 15036 11204 15088
rect 11796 15036 11848 15088
rect 3608 14968 3660 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 7380 15011 7432 15020
rect 7380 14977 7414 15011
rect 7414 14977 7432 15011
rect 7380 14968 7432 14977
rect 10968 14968 11020 15020
rect 14832 14968 14884 15020
rect 19340 15104 19392 15156
rect 22100 15104 22152 15156
rect 22192 15104 22244 15156
rect 41880 15104 41932 15156
rect 19432 15036 19484 15088
rect 20444 15036 20496 15088
rect 22652 15036 22704 15088
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 39580 15011 39632 15020
rect 39580 14977 39614 15011
rect 39614 14977 39632 15011
rect 39580 14968 39632 14977
rect 43812 15011 43864 15020
rect 43812 14977 43821 15011
rect 43821 14977 43855 15011
rect 43855 14977 43864 15011
rect 43812 14968 43864 14977
rect 45836 14968 45888 15020
rect 20628 14900 20680 14952
rect 39120 14900 39172 14952
rect 8576 14832 8628 14884
rect 13728 14832 13780 14884
rect 5632 14764 5684 14816
rect 9312 14764 9364 14816
rect 11704 14764 11756 14816
rect 13084 14764 13136 14816
rect 14556 14764 14608 14816
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 20260 14764 20312 14816
rect 21916 14764 21968 14816
rect 41144 14807 41196 14816
rect 41144 14773 41153 14807
rect 41153 14773 41187 14807
rect 41187 14773 41196 14807
rect 41144 14764 41196 14773
rect 45560 14764 45612 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3608 14560 3660 14612
rect 7380 14560 7432 14612
rect 8852 14560 8904 14612
rect 11796 14560 11848 14612
rect 17132 14560 17184 14612
rect 20444 14560 20496 14612
rect 20628 14560 20680 14612
rect 21916 14603 21968 14612
rect 9128 14535 9180 14544
rect 9128 14501 9137 14535
rect 9137 14501 9171 14535
rect 9171 14501 9180 14535
rect 9128 14492 9180 14501
rect 4528 14356 4580 14408
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 8208 14424 8260 14476
rect 8576 14467 8628 14476
rect 8576 14433 8585 14467
rect 8585 14433 8619 14467
rect 8619 14433 8628 14467
rect 8576 14424 8628 14433
rect 9220 14424 9272 14476
rect 7656 14356 7708 14408
rect 11796 14424 11848 14476
rect 15108 14424 15160 14476
rect 19800 14492 19852 14544
rect 11336 14356 11388 14408
rect 13084 14399 13136 14408
rect 9312 14331 9364 14340
rect 9312 14297 9339 14331
rect 9339 14297 9364 14331
rect 9312 14288 9364 14297
rect 9588 14288 9640 14340
rect 10508 14288 10560 14340
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 15752 14356 15804 14408
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 8116 14220 8168 14272
rect 11244 14220 11296 14272
rect 11796 14220 11848 14272
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 19340 14424 19392 14476
rect 21916 14569 21925 14603
rect 21925 14569 21959 14603
rect 21959 14569 21968 14603
rect 21916 14560 21968 14569
rect 41972 14560 42024 14612
rect 45836 14603 45888 14612
rect 45836 14569 45845 14603
rect 45845 14569 45879 14603
rect 45879 14569 45888 14603
rect 45836 14560 45888 14569
rect 17776 14356 17828 14365
rect 19156 14356 19208 14408
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 22192 14356 22244 14408
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 39948 14356 40000 14408
rect 40316 14399 40368 14408
rect 40316 14365 40350 14399
rect 40350 14365 40368 14399
rect 40316 14356 40368 14365
rect 43352 14356 43404 14408
rect 43812 14356 43864 14408
rect 45192 14399 45244 14408
rect 45192 14365 45201 14399
rect 45201 14365 45235 14399
rect 45235 14365 45244 14399
rect 45192 14356 45244 14365
rect 19984 14288 20036 14340
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 43720 14288 43772 14340
rect 45284 14220 45336 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4896 14016 4948 14068
rect 5540 14016 5592 14068
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 8852 14059 8904 14068
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 14464 14016 14516 14068
rect 20260 14016 20312 14068
rect 4620 13948 4672 14000
rect 4252 13880 4304 13932
rect 4804 13880 4856 13932
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 10968 13948 11020 14000
rect 11336 13948 11388 14000
rect 9220 13880 9272 13932
rect 8024 13812 8076 13864
rect 11244 13880 11296 13932
rect 12624 13948 12676 14000
rect 14280 13948 14332 14000
rect 14832 13948 14884 14000
rect 19984 13948 20036 14000
rect 20628 13948 20680 14000
rect 12808 13880 12860 13932
rect 15108 13880 15160 13932
rect 20444 13880 20496 13932
rect 42156 14016 42208 14068
rect 44180 14016 44232 14068
rect 41144 13948 41196 14000
rect 45192 13948 45244 14000
rect 43352 13880 43404 13932
rect 44456 13880 44508 13932
rect 45560 13923 45612 13932
rect 45560 13889 45569 13923
rect 45569 13889 45603 13923
rect 45603 13889 45612 13923
rect 45560 13880 45612 13889
rect 11796 13812 11848 13864
rect 20352 13812 20404 13864
rect 39120 13812 39172 13864
rect 39948 13812 40000 13864
rect 11244 13744 11296 13796
rect 11704 13676 11756 13728
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 45284 13719 45336 13728
rect 45284 13685 45293 13719
rect 45293 13685 45327 13719
rect 45327 13685 45336 13719
rect 45284 13676 45336 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 12624 13515 12676 13524
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 17132 13515 17184 13524
rect 17132 13481 17141 13515
rect 17141 13481 17175 13515
rect 17175 13481 17184 13515
rect 17132 13472 17184 13481
rect 20076 13472 20128 13524
rect 21456 13472 21508 13524
rect 5632 13404 5684 13456
rect 5540 13336 5592 13388
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 4896 13268 4948 13320
rect 12532 13404 12584 13456
rect 12900 13404 12952 13456
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 43352 13472 43404 13524
rect 44456 13472 44508 13524
rect 5172 13200 5224 13252
rect 6644 13268 6696 13320
rect 8116 13268 8168 13320
rect 8576 13268 8628 13320
rect 11060 13268 11112 13320
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 11336 13200 11388 13252
rect 12256 13200 12308 13252
rect 16028 13311 16080 13320
rect 16028 13277 16062 13311
rect 16062 13277 16080 13311
rect 16028 13268 16080 13277
rect 12900 13200 12952 13252
rect 20444 13268 20496 13320
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 20536 13200 20588 13252
rect 43260 13243 43312 13252
rect 43260 13209 43294 13243
rect 43294 13209 43312 13243
rect 43260 13200 43312 13209
rect 4988 13132 5040 13184
rect 8208 13132 8260 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 10968 13132 11020 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 5172 12928 5224 12980
rect 8116 12928 8168 12980
rect 11060 12971 11112 12980
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 12808 12971 12860 12980
rect 4896 12792 4948 12801
rect 5632 12792 5684 12844
rect 7380 12792 7432 12844
rect 8024 12792 8076 12844
rect 9036 12860 9088 12912
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 43260 12971 43312 12980
rect 43260 12937 43269 12971
rect 43269 12937 43303 12971
rect 43303 12937 43312 12971
rect 43260 12928 43312 12937
rect 45284 12928 45336 12980
rect 11888 12860 11940 12912
rect 40040 12860 40092 12912
rect 43812 12903 43864 12912
rect 43812 12869 43821 12903
rect 43821 12869 43855 12903
rect 43855 12869 43864 12903
rect 43812 12860 43864 12869
rect 44180 12903 44232 12912
rect 44180 12869 44189 12903
rect 44189 12869 44223 12903
rect 44223 12869 44232 12903
rect 44180 12860 44232 12869
rect 8576 12792 8628 12844
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 10968 12792 11020 12844
rect 12256 12792 12308 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 11796 12724 11848 12776
rect 39120 12767 39172 12776
rect 9404 12656 9456 12708
rect 39120 12733 39129 12767
rect 39129 12733 39163 12767
rect 39163 12733 39172 12767
rect 39120 12724 39172 12733
rect 12256 12656 12308 12708
rect 7748 12588 7800 12640
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 9588 12588 9640 12640
rect 11796 12588 11848 12640
rect 40868 12588 40920 12640
rect 43076 12631 43128 12640
rect 43076 12597 43085 12631
rect 43085 12597 43119 12631
rect 43119 12597 43128 12631
rect 43076 12588 43128 12597
rect 44456 12588 44508 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 8208 12316 8260 12368
rect 9588 12384 9640 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 9404 12316 9456 12368
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 5448 12180 5500 12232
rect 7748 12180 7800 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10784 12223 10836 12232
rect 10784 12189 10818 12223
rect 10818 12189 10836 12223
rect 38844 12223 38896 12232
rect 10784 12180 10836 12189
rect 38844 12189 38853 12223
rect 38853 12189 38887 12223
rect 38887 12189 38896 12223
rect 38844 12180 38896 12189
rect 39304 12223 39356 12232
rect 39304 12189 39313 12223
rect 39313 12189 39347 12223
rect 39347 12189 39356 12223
rect 39304 12180 39356 12189
rect 42892 12223 42944 12232
rect 42892 12189 42901 12223
rect 42901 12189 42935 12223
rect 42935 12189 42944 12223
rect 42892 12180 42944 12189
rect 7288 12112 7340 12164
rect 8392 12112 8444 12164
rect 7104 12044 7156 12096
rect 41604 12087 41656 12096
rect 41604 12053 41613 12087
rect 41613 12053 41647 12087
rect 41647 12053 41656 12087
rect 41604 12044 41656 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 9036 11840 9088 11892
rect 43076 11840 43128 11892
rect 12256 11772 12308 11824
rect 39304 11815 39356 11824
rect 39304 11781 39338 11815
rect 39338 11781 39356 11815
rect 39304 11772 39356 11781
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 39120 11704 39172 11756
rect 39580 11704 39632 11756
rect 41420 11704 41472 11756
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 4712 11568 4764 11620
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 11888 11500 11940 11552
rect 38384 11543 38436 11552
rect 38384 11509 38393 11543
rect 38393 11509 38427 11543
rect 38427 11509 38436 11543
rect 38384 11500 38436 11509
rect 40868 11543 40920 11552
rect 40868 11509 40877 11543
rect 40877 11509 40911 11543
rect 40911 11509 40920 11543
rect 40868 11500 40920 11509
rect 42432 11500 42484 11552
rect 44732 11500 44784 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12256 11296 12308 11348
rect 39580 11296 39632 11348
rect 41420 11339 41472 11348
rect 41420 11305 41429 11339
rect 41429 11305 41463 11339
rect 41463 11305 41472 11339
rect 41420 11296 41472 11305
rect 44456 11339 44508 11348
rect 44456 11305 44465 11339
rect 44465 11305 44499 11339
rect 44499 11305 44508 11339
rect 44456 11296 44508 11305
rect 5448 11160 5500 11212
rect 10508 11160 10560 11212
rect 2688 11092 2740 11144
rect 6460 11092 6512 11144
rect 20352 11135 20404 11144
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 39120 11092 39172 11144
rect 41604 11092 41656 11144
rect 44180 11135 44232 11144
rect 44180 11101 44189 11135
rect 44189 11101 44223 11135
rect 44223 11101 44232 11135
rect 44180 11092 44232 11101
rect 45836 11092 45888 11144
rect 2228 11067 2280 11076
rect 2228 11033 2262 11067
rect 2262 11033 2280 11067
rect 2228 11024 2280 11033
rect 4344 11067 4396 11076
rect 4344 11033 4353 11067
rect 4353 11033 4387 11067
rect 4387 11033 4396 11067
rect 4344 11024 4396 11033
rect 5816 11024 5868 11076
rect 11704 11024 11756 11076
rect 38384 11067 38436 11076
rect 38384 11033 38418 11067
rect 38418 11033 38436 11067
rect 38384 11024 38436 11033
rect 38844 11024 38896 11076
rect 42432 11067 42484 11076
rect 42432 11033 42466 11067
rect 42466 11033 42484 11067
rect 42432 11024 42484 11033
rect 42524 11024 42576 11076
rect 43996 11067 44048 11076
rect 43996 11033 44005 11067
rect 44005 11033 44039 11067
rect 44039 11033 44048 11067
rect 43996 11024 44048 11033
rect 3332 10999 3384 11008
rect 3332 10965 3341 10999
rect 3341 10965 3375 10999
rect 3375 10965 3384 10999
rect 3332 10956 3384 10965
rect 6920 10956 6972 11008
rect 20260 10956 20312 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 9772 10752 9824 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 43996 10795 44048 10804
rect 43996 10761 44005 10795
rect 44005 10761 44039 10795
rect 44039 10761 44048 10795
rect 43996 10752 44048 10761
rect 45836 10795 45888 10804
rect 45836 10761 45845 10795
rect 45845 10761 45879 10795
rect 45879 10761 45888 10795
rect 45836 10752 45888 10761
rect 2688 10616 2740 10668
rect 4344 10684 4396 10736
rect 5448 10684 5500 10736
rect 9496 10684 9548 10736
rect 44732 10727 44784 10736
rect 3976 10616 4028 10668
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 2780 10548 2832 10600
rect 4620 10548 4672 10600
rect 7656 10616 7708 10668
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 40132 10659 40184 10668
rect 40132 10625 40141 10659
rect 40141 10625 40175 10659
rect 40175 10625 40184 10659
rect 40132 10616 40184 10625
rect 42524 10616 42576 10668
rect 44732 10693 44766 10727
rect 44766 10693 44784 10727
rect 44732 10684 44784 10693
rect 44456 10591 44508 10600
rect 44456 10557 44465 10591
rect 44465 10557 44499 10591
rect 44499 10557 44508 10591
rect 44456 10548 44508 10557
rect 4068 10412 4120 10464
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 8208 10412 8260 10464
rect 40592 10412 40644 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2688 10208 2740 10260
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 4620 10208 4672 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 44180 10208 44232 10260
rect 4712 10072 4764 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 42524 10115 42576 10124
rect 42524 10081 42533 10115
rect 42533 10081 42567 10115
rect 42567 10081 42576 10115
rect 42524 10072 42576 10081
rect 44456 10072 44508 10124
rect 3332 10004 3384 10056
rect 4804 10004 4856 10056
rect 5724 10047 5776 10056
rect 5724 10013 5758 10047
rect 5758 10013 5776 10047
rect 5724 10004 5776 10013
rect 20260 10047 20312 10056
rect 20260 10013 20294 10047
rect 20294 10013 20312 10047
rect 20260 10004 20312 10013
rect 45284 10004 45336 10056
rect 4988 9936 5040 9988
rect 42800 9979 42852 9988
rect 42800 9945 42834 9979
rect 42834 9945 42852 9979
rect 42800 9936 42852 9945
rect 1860 9868 1912 9920
rect 22008 9868 22060 9920
rect 57520 9868 57572 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 5816 9528 5868 9580
rect 42524 9596 42576 9648
rect 40592 9528 40644 9580
rect 42800 9571 42852 9580
rect 42800 9537 42809 9571
rect 42809 9537 42843 9571
rect 42843 9537 42852 9571
rect 42800 9528 42852 9537
rect 42616 9324 42668 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 57520 3723 57572 3732
rect 57520 3689 57529 3723
rect 57529 3689 57563 3723
rect 57563 3689 57572 3723
rect 57520 3680 57572 3689
rect 57520 3476 57572 3528
rect 58256 3383 58308 3392
rect 58256 3349 58265 3383
rect 58265 3349 58299 3383
rect 58299 3349 58308 3383
rect 58256 3340 58308 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 42616 2431 42668 2440
rect 42616 2397 42625 2431
rect 42625 2397 42659 2431
rect 42659 2397 42668 2431
rect 42616 2388 42668 2397
rect 20 2252 72 2304
rect 21272 2252 21324 2304
rect 42524 2252 42576 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 6458 59200 6514 59800
rect 28354 59200 28410 59800
rect 49606 59200 49662 59800
rect 6472 57594 6500 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 28368 57594 28396 59200
rect 49620 57610 49648 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 49620 57594 49740 57610
rect 6460 57588 6512 57594
rect 6460 57530 6512 57536
rect 28356 57588 28408 57594
rect 49620 57588 49752 57594
rect 49620 57582 49700 57588
rect 28356 57530 28408 57536
rect 49700 57530 49752 57536
rect 6644 57452 6696 57458
rect 6644 57394 6696 57400
rect 28540 57452 28592 57458
rect 28540 57394 28592 57400
rect 46572 57452 46624 57458
rect 46572 57394 46624 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 6656 46170 6684 57394
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 6644 46164 6696 46170
rect 6644 46106 6696 46112
rect 6736 45960 6788 45966
rect 6736 45902 6788 45908
rect 5816 45892 5868 45898
rect 5816 45834 5868 45840
rect 5828 45626 5856 45834
rect 5816 45620 5868 45626
rect 5816 45562 5868 45568
rect 6748 45354 6776 45902
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 9128 45552 9180 45558
rect 9128 45494 9180 45500
rect 7104 45484 7156 45490
rect 7104 45426 7156 45432
rect 8300 45484 8352 45490
rect 8300 45426 8352 45432
rect 6736 45348 6788 45354
rect 6736 45290 6788 45296
rect 6920 45348 6972 45354
rect 6920 45290 6972 45296
rect 6460 45280 6512 45286
rect 6460 45222 6512 45228
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 3436 27878 3464 44911
rect 6472 44878 6500 45222
rect 6748 44946 6776 45290
rect 6736 44940 6788 44946
rect 6736 44882 6788 44888
rect 6460 44872 6512 44878
rect 6460 44814 6512 44820
rect 6828 44872 6880 44878
rect 6828 44814 6880 44820
rect 5908 44736 5960 44742
rect 5908 44678 5960 44684
rect 5920 44402 5948 44678
rect 5908 44396 5960 44402
rect 5908 44338 5960 44344
rect 5632 44260 5684 44266
rect 5632 44202 5684 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 5644 43382 5672 44202
rect 5920 43994 5948 44338
rect 6840 44334 6868 44814
rect 6828 44328 6880 44334
rect 6828 44270 6880 44276
rect 5908 43988 5960 43994
rect 5908 43930 5960 43936
rect 6840 43722 6868 44270
rect 6276 43716 6328 43722
rect 6276 43658 6328 43664
rect 6828 43716 6880 43722
rect 6828 43658 6880 43664
rect 5632 43376 5684 43382
rect 5632 43318 5684 43324
rect 6288 43314 6316 43658
rect 6276 43308 6328 43314
rect 6276 43250 6328 43256
rect 5908 43104 5960 43110
rect 5908 43046 5960 43052
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 5724 42628 5776 42634
rect 5724 42570 5776 42576
rect 5736 42362 5764 42570
rect 5724 42356 5776 42362
rect 5724 42298 5776 42304
rect 5920 42226 5948 43046
rect 6288 42906 6316 43250
rect 6276 42900 6328 42906
rect 6276 42842 6328 42848
rect 6736 42900 6788 42906
rect 6736 42842 6788 42848
rect 6748 42226 6776 42842
rect 6932 42702 6960 45290
rect 7012 44736 7064 44742
rect 7012 44678 7064 44684
rect 7024 44470 7052 44678
rect 7116 44538 7144 45426
rect 7380 45416 7432 45422
rect 7380 45358 7432 45364
rect 7288 44872 7340 44878
rect 7288 44814 7340 44820
rect 7104 44532 7156 44538
rect 7104 44474 7156 44480
rect 7300 44470 7328 44814
rect 7012 44464 7064 44470
rect 7012 44406 7064 44412
rect 7288 44464 7340 44470
rect 7288 44406 7340 44412
rect 7024 43382 7052 44406
rect 7104 43648 7156 43654
rect 7104 43590 7156 43596
rect 7012 43376 7064 43382
rect 7012 43318 7064 43324
rect 7116 43314 7144 43590
rect 7104 43308 7156 43314
rect 7104 43250 7156 43256
rect 7116 42922 7144 43250
rect 7024 42894 7144 42922
rect 6920 42696 6972 42702
rect 6920 42638 6972 42644
rect 7024 42634 7052 42894
rect 7104 42696 7156 42702
rect 7104 42638 7156 42644
rect 7288 42696 7340 42702
rect 7288 42638 7340 42644
rect 7012 42628 7064 42634
rect 7012 42570 7064 42576
rect 7024 42226 7052 42570
rect 7116 42226 7144 42638
rect 7196 42560 7248 42566
rect 7196 42502 7248 42508
rect 5908 42220 5960 42226
rect 5908 42162 5960 42168
rect 6736 42220 6788 42226
rect 6736 42162 6788 42168
rect 7012 42220 7064 42226
rect 7012 42162 7064 42168
rect 7104 42220 7156 42226
rect 7104 42162 7156 42168
rect 5908 42016 5960 42022
rect 5908 41958 5960 41964
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 5920 41614 5948 41958
rect 7116 41818 7144 42162
rect 7104 41812 7156 41818
rect 7104 41754 7156 41760
rect 7208 41614 7236 42502
rect 7300 41682 7328 42638
rect 7392 42566 7420 45358
rect 7656 45280 7708 45286
rect 7656 45222 7708 45228
rect 7668 45082 7696 45222
rect 8312 45082 8340 45426
rect 7656 45076 7708 45082
rect 7656 45018 7708 45024
rect 8300 45076 8352 45082
rect 8300 45018 8352 45024
rect 9036 45076 9088 45082
rect 9036 45018 9088 45024
rect 9048 44470 9076 45018
rect 9140 44538 9168 45494
rect 9680 45484 9732 45490
rect 9680 45426 9732 45432
rect 27252 45484 27304 45490
rect 27252 45426 27304 45432
rect 9692 44742 9720 45426
rect 10784 45008 10836 45014
rect 10784 44950 10836 44956
rect 10048 44804 10100 44810
rect 10048 44746 10100 44752
rect 9680 44736 9732 44742
rect 9956 44736 10008 44742
rect 9732 44684 9904 44690
rect 9680 44678 9904 44684
rect 9956 44678 10008 44684
rect 9692 44662 9904 44678
rect 9128 44532 9180 44538
rect 9128 44474 9180 44480
rect 9036 44464 9088 44470
rect 9036 44406 9088 44412
rect 9680 44396 9732 44402
rect 9680 44338 9732 44344
rect 9692 43994 9720 44338
rect 9772 44328 9824 44334
rect 9772 44270 9824 44276
rect 9680 43988 9732 43994
rect 9680 43930 9732 43936
rect 9784 43790 9812 44270
rect 9876 43858 9904 44662
rect 9968 44538 9996 44678
rect 9956 44532 10008 44538
rect 9956 44474 10008 44480
rect 9864 43852 9916 43858
rect 9864 43794 9916 43800
rect 9772 43784 9824 43790
rect 9968 43738 9996 44474
rect 10060 44198 10088 44746
rect 10048 44192 10100 44198
rect 10048 44134 10100 44140
rect 10508 44192 10560 44198
rect 10508 44134 10560 44140
rect 9772 43726 9824 43732
rect 9128 43716 9180 43722
rect 9128 43658 9180 43664
rect 9140 43382 9168 43658
rect 7656 43376 7708 43382
rect 7656 43318 7708 43324
rect 9128 43376 9180 43382
rect 9128 43318 9180 43324
rect 7668 42838 7696 43318
rect 8760 43308 8812 43314
rect 8760 43250 8812 43256
rect 7656 42832 7708 42838
rect 7656 42774 7708 42780
rect 7380 42560 7432 42566
rect 7380 42502 7432 42508
rect 7668 41818 7696 42774
rect 8300 42628 8352 42634
rect 8300 42570 8352 42576
rect 8312 42226 8340 42570
rect 8300 42220 8352 42226
rect 8300 42162 8352 42168
rect 7656 41812 7708 41818
rect 7656 41754 7708 41760
rect 7288 41676 7340 41682
rect 7288 41618 7340 41624
rect 5264 41608 5316 41614
rect 5264 41550 5316 41556
rect 5908 41608 5960 41614
rect 5908 41550 5960 41556
rect 7196 41608 7248 41614
rect 7196 41550 7248 41556
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 5276 40594 5304 41550
rect 5540 40928 5592 40934
rect 5540 40870 5592 40876
rect 5264 40588 5316 40594
rect 5264 40530 5316 40536
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 5276 39506 5304 40530
rect 5552 40526 5580 40870
rect 5540 40520 5592 40526
rect 5540 40462 5592 40468
rect 6920 40384 6972 40390
rect 6920 40326 6972 40332
rect 6644 39976 6696 39982
rect 6644 39918 6696 39924
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 5264 39500 5316 39506
rect 5264 39442 5316 39448
rect 5276 38826 5304 39442
rect 5552 39438 5580 39782
rect 6656 39642 6684 39918
rect 6932 39846 6960 40326
rect 7208 40186 7236 41550
rect 8576 41064 8628 41070
rect 8576 41006 8628 41012
rect 8588 40730 8616 41006
rect 8576 40724 8628 40730
rect 8576 40666 8628 40672
rect 7196 40180 7248 40186
rect 7196 40122 7248 40128
rect 8772 40050 8800 43250
rect 9140 42906 9168 43318
rect 9784 43110 9812 43726
rect 9876 43710 9996 43738
rect 9876 43654 9904 43710
rect 9864 43648 9916 43654
rect 9864 43590 9916 43596
rect 9772 43104 9824 43110
rect 9772 43046 9824 43052
rect 9128 42900 9180 42906
rect 9128 42842 9180 42848
rect 9036 42628 9088 42634
rect 9036 42570 9088 42576
rect 9048 42362 9076 42570
rect 9036 42356 9088 42362
rect 9036 42298 9088 42304
rect 9140 42226 9168 42842
rect 9784 42702 9812 43046
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9128 42220 9180 42226
rect 9128 42162 9180 42168
rect 9784 41682 9812 42638
rect 9876 42158 9904 43590
rect 10520 42566 10548 44134
rect 10796 43722 10824 44950
rect 11152 44872 11204 44878
rect 11152 44814 11204 44820
rect 11164 44538 11192 44814
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 11152 44532 11204 44538
rect 11152 44474 11204 44480
rect 24860 44192 24912 44198
rect 24860 44134 24912 44140
rect 24872 43790 24900 44134
rect 24584 43784 24636 43790
rect 24584 43726 24636 43732
rect 24860 43784 24912 43790
rect 24860 43726 24912 43732
rect 10784 43716 10836 43722
rect 10784 43658 10836 43664
rect 10968 43716 11020 43722
rect 10968 43658 11020 43664
rect 12348 43716 12400 43722
rect 12348 43658 12400 43664
rect 10980 43450 11008 43658
rect 10968 43444 11020 43450
rect 10968 43386 11020 43392
rect 12360 43314 12388 43658
rect 13268 43648 13320 43654
rect 13268 43590 13320 43596
rect 10968 43308 11020 43314
rect 10968 43250 11020 43256
rect 12348 43308 12400 43314
rect 12348 43250 12400 43256
rect 10508 42560 10560 42566
rect 10508 42502 10560 42508
rect 10520 42294 10548 42502
rect 10980 42362 11008 43250
rect 10968 42356 11020 42362
rect 10968 42298 11020 42304
rect 10508 42288 10560 42294
rect 10508 42230 10560 42236
rect 9864 42152 9916 42158
rect 9864 42094 9916 42100
rect 12072 42016 12124 42022
rect 12072 41958 12124 41964
rect 9128 41676 9180 41682
rect 9128 41618 9180 41624
rect 9772 41676 9824 41682
rect 9772 41618 9824 41624
rect 9140 41138 9168 41618
rect 9404 41608 9456 41614
rect 9404 41550 9456 41556
rect 9128 41132 9180 41138
rect 9128 41074 9180 41080
rect 9140 40594 9168 41074
rect 9128 40588 9180 40594
rect 9128 40530 9180 40536
rect 9416 40526 9444 41550
rect 11152 41540 11204 41546
rect 11152 41482 11204 41488
rect 11164 41138 11192 41482
rect 11152 41132 11204 41138
rect 11152 41074 11204 41080
rect 11152 40928 11204 40934
rect 11152 40870 11204 40876
rect 9404 40520 9456 40526
rect 9404 40462 9456 40468
rect 7656 40044 7708 40050
rect 7656 39986 7708 39992
rect 8760 40044 8812 40050
rect 8760 39986 8812 39992
rect 6920 39840 6972 39846
rect 6920 39782 6972 39788
rect 7668 39642 7696 39986
rect 11060 39908 11112 39914
rect 11060 39850 11112 39856
rect 9220 39840 9272 39846
rect 9220 39782 9272 39788
rect 6644 39636 6696 39642
rect 6644 39578 6696 39584
rect 7288 39636 7340 39642
rect 7288 39578 7340 39584
rect 7656 39636 7708 39642
rect 7656 39578 7708 39584
rect 5540 39432 5592 39438
rect 5540 39374 5592 39380
rect 7196 39364 7248 39370
rect 7196 39306 7248 39312
rect 5264 38820 5316 38826
rect 5264 38762 5316 38768
rect 6920 38820 6972 38826
rect 6920 38762 6972 38768
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 5276 38418 5304 38762
rect 5540 38752 5592 38758
rect 5540 38694 5592 38700
rect 5264 38412 5316 38418
rect 5264 38354 5316 38360
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5276 37330 5304 38354
rect 5552 38350 5580 38694
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 6932 38010 6960 38762
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 6920 38004 6972 38010
rect 6920 37946 6972 37952
rect 7024 37874 7052 38694
rect 7012 37868 7064 37874
rect 7012 37810 7064 37816
rect 5816 37664 5868 37670
rect 5816 37606 5868 37612
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5828 37262 5856 37606
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 7208 37126 7236 39306
rect 7300 38486 7328 39578
rect 7380 39500 7432 39506
rect 7380 39442 7432 39448
rect 7288 38480 7340 38486
rect 7288 38422 7340 38428
rect 7392 38010 7420 39442
rect 9232 39438 9260 39782
rect 7472 39432 7524 39438
rect 7472 39374 7524 39380
rect 8392 39432 8444 39438
rect 8392 39374 8444 39380
rect 8760 39432 8812 39438
rect 8760 39374 8812 39380
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 7484 38554 7512 39374
rect 7472 38548 7524 38554
rect 7472 38490 7524 38496
rect 8404 38350 8432 39374
rect 8772 38758 8800 39374
rect 11072 39098 11100 39850
rect 11164 39642 11192 40870
rect 12084 40526 12112 41958
rect 13280 41818 13308 43590
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 24216 42696 24268 42702
rect 24216 42638 24268 42644
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 24228 42294 24256 42638
rect 24216 42288 24268 42294
rect 24216 42230 24268 42236
rect 23388 42152 23440 42158
rect 23388 42094 23440 42100
rect 15292 42016 15344 42022
rect 15292 41958 15344 41964
rect 23020 42016 23072 42022
rect 23020 41958 23072 41964
rect 13268 41812 13320 41818
rect 13268 41754 13320 41760
rect 13176 41608 13228 41614
rect 13176 41550 13228 41556
rect 13268 41608 13320 41614
rect 13268 41550 13320 41556
rect 14924 41608 14976 41614
rect 14924 41550 14976 41556
rect 12440 41472 12492 41478
rect 12440 41414 12492 41420
rect 11796 40520 11848 40526
rect 11796 40462 11848 40468
rect 12072 40520 12124 40526
rect 12072 40462 12124 40468
rect 11244 40384 11296 40390
rect 11244 40326 11296 40332
rect 11152 39636 11204 39642
rect 11152 39578 11204 39584
rect 11256 39438 11284 40326
rect 11244 39432 11296 39438
rect 11244 39374 11296 39380
rect 11060 39092 11112 39098
rect 11060 39034 11112 39040
rect 8760 38752 8812 38758
rect 8760 38694 8812 38700
rect 8772 38350 8800 38694
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8760 38344 8812 38350
rect 8760 38286 8812 38292
rect 9772 38344 9824 38350
rect 9772 38286 9824 38292
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 7380 38004 7432 38010
rect 7380 37946 7432 37952
rect 8772 37942 8800 38286
rect 8760 37936 8812 37942
rect 8760 37878 8812 37884
rect 9784 37806 9812 38286
rect 10612 37942 10640 38286
rect 10600 37936 10652 37942
rect 10600 37878 10652 37884
rect 9772 37800 9824 37806
rect 9772 37742 9824 37748
rect 9784 37262 9812 37742
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3424 27872 3476 27878
rect 3424 27814 3476 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 11072 23594 11100 39034
rect 11704 38752 11756 38758
rect 11704 38694 11756 38700
rect 11716 38282 11744 38694
rect 11808 38350 11836 40462
rect 12452 40186 12480 41414
rect 13188 40730 13216 41550
rect 13280 41274 13308 41550
rect 13452 41472 13504 41478
rect 13452 41414 13504 41420
rect 13268 41268 13320 41274
rect 13268 41210 13320 41216
rect 13176 40724 13228 40730
rect 13176 40666 13228 40672
rect 12440 40180 12492 40186
rect 12440 40122 12492 40128
rect 13176 40044 13228 40050
rect 13176 39986 13228 39992
rect 13188 39642 13216 39986
rect 13464 39846 13492 41414
rect 14936 41070 14964 41550
rect 15200 41132 15252 41138
rect 15200 41074 15252 41080
rect 13820 41064 13872 41070
rect 13820 41006 13872 41012
rect 14924 41064 14976 41070
rect 14924 41006 14976 41012
rect 13832 40594 13860 41006
rect 13820 40588 13872 40594
rect 13820 40530 13872 40536
rect 14924 40588 14976 40594
rect 14924 40530 14976 40536
rect 13832 40458 13860 40530
rect 13820 40452 13872 40458
rect 13820 40394 13872 40400
rect 13832 40118 13860 40394
rect 13820 40112 13872 40118
rect 13820 40054 13872 40060
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13176 39636 13228 39642
rect 13176 39578 13228 39584
rect 13556 38554 13584 39918
rect 14936 39506 14964 40530
rect 15212 39642 15240 41074
rect 15200 39636 15252 39642
rect 15200 39578 15252 39584
rect 14924 39500 14976 39506
rect 14924 39442 14976 39448
rect 15304 39438 15332 41958
rect 22100 41608 22152 41614
rect 22100 41550 22152 41556
rect 21088 41540 21140 41546
rect 21088 41482 21140 41488
rect 16764 41472 16816 41478
rect 16764 41414 16816 41420
rect 16776 40730 16804 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 21100 41138 21128 41482
rect 22112 41274 22140 41550
rect 22744 41472 22796 41478
rect 22744 41414 22796 41420
rect 22100 41268 22152 41274
rect 22100 41210 22152 41216
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 16856 40928 16908 40934
rect 16856 40870 16908 40876
rect 16764 40724 16816 40730
rect 16764 40666 16816 40672
rect 16868 40594 16896 40870
rect 22112 40594 22140 41210
rect 22756 41206 22784 41414
rect 22744 41200 22796 41206
rect 22744 41142 22796 41148
rect 22928 41064 22980 41070
rect 22928 41006 22980 41012
rect 22284 40928 22336 40934
rect 22284 40870 22336 40876
rect 16856 40588 16908 40594
rect 16856 40530 16908 40536
rect 22100 40588 22152 40594
rect 22100 40530 22152 40536
rect 16764 40452 16816 40458
rect 16764 40394 16816 40400
rect 16776 39642 16804 40394
rect 17224 40384 17276 40390
rect 17224 40326 17276 40332
rect 17236 40118 17264 40326
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 17224 40112 17276 40118
rect 17224 40054 17276 40060
rect 22112 40050 22140 40530
rect 22296 40050 22324 40870
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 16764 39636 16816 39642
rect 16764 39578 16816 39584
rect 22112 39506 22140 39986
rect 22100 39500 22152 39506
rect 22100 39442 22152 39448
rect 15292 39432 15344 39438
rect 15292 39374 15344 39380
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 22112 38962 22140 39442
rect 22480 39438 22508 40462
rect 22940 40186 22968 41006
rect 23032 40934 23060 41958
rect 23400 41274 23428 42094
rect 24596 41682 24624 43726
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 24768 42220 24820 42226
rect 24768 42162 24820 42168
rect 24584 41676 24636 41682
rect 24584 41618 24636 41624
rect 23388 41268 23440 41274
rect 23388 41210 23440 41216
rect 24492 41132 24544 41138
rect 24492 41074 24544 41080
rect 23572 41064 23624 41070
rect 23572 41006 23624 41012
rect 23020 40928 23072 40934
rect 23020 40870 23072 40876
rect 23204 40928 23256 40934
rect 23204 40870 23256 40876
rect 23216 40526 23244 40870
rect 23204 40520 23256 40526
rect 23204 40462 23256 40468
rect 22928 40180 22980 40186
rect 22928 40122 22980 40128
rect 23584 39642 23612 41006
rect 24504 40730 24532 41074
rect 24492 40724 24544 40730
rect 24492 40666 24544 40672
rect 24780 40458 24808 42162
rect 25228 41608 25280 41614
rect 25228 41550 25280 41556
rect 24216 40452 24268 40458
rect 24216 40394 24268 40400
rect 24768 40452 24820 40458
rect 24768 40394 24820 40400
rect 24228 39846 24256 40394
rect 25240 40050 25268 41550
rect 25516 40934 25544 43590
rect 25596 42016 25648 42022
rect 25596 41958 25648 41964
rect 25608 41070 25636 41958
rect 27264 41818 27292 45426
rect 28552 45354 28580 57394
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 45560 49224 45612 49230
rect 45560 49166 45612 49172
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 40500 45960 40552 45966
rect 40500 45902 40552 45908
rect 44272 45960 44324 45966
rect 44272 45902 44324 45908
rect 40512 45558 40540 45902
rect 29000 45552 29052 45558
rect 29000 45494 29052 45500
rect 40500 45552 40552 45558
rect 40500 45494 40552 45500
rect 28540 45348 28592 45354
rect 28540 45290 28592 45296
rect 29012 42090 29040 45494
rect 44284 45490 44312 45902
rect 44272 45484 44324 45490
rect 44272 45426 44324 45432
rect 44456 45484 44508 45490
rect 44456 45426 44508 45432
rect 40132 45416 40184 45422
rect 40132 45358 40184 45364
rect 37740 45280 37792 45286
rect 37740 45222 37792 45228
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 36268 44804 36320 44810
rect 36268 44746 36320 44752
rect 37280 44804 37332 44810
rect 37280 44746 37332 44752
rect 36280 44402 36308 44746
rect 36268 44396 36320 44402
rect 36268 44338 36320 44344
rect 37292 44334 37320 44746
rect 37752 44402 37780 45222
rect 40144 44878 40172 45358
rect 41512 45280 41564 45286
rect 41512 45222 41564 45228
rect 40132 44872 40184 44878
rect 40132 44814 40184 44820
rect 41052 44872 41104 44878
rect 41052 44814 41104 44820
rect 38476 44736 38528 44742
rect 38476 44678 38528 44684
rect 37740 44396 37792 44402
rect 37740 44338 37792 44344
rect 37280 44328 37332 44334
rect 37280 44270 37332 44276
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 37292 43790 37320 44270
rect 37740 44192 37792 44198
rect 37740 44134 37792 44140
rect 37280 43784 37332 43790
rect 37280 43726 37332 43732
rect 37292 43246 37320 43726
rect 37752 43382 37780 44134
rect 38488 43994 38516 44678
rect 40144 44402 40172 44814
rect 40132 44396 40184 44402
rect 40132 44338 40184 44344
rect 38752 44192 38804 44198
rect 38752 44134 38804 44140
rect 38476 43988 38528 43994
rect 38476 43930 38528 43936
rect 38660 43852 38712 43858
rect 38660 43794 38712 43800
rect 38672 43450 38700 43794
rect 38764 43790 38792 44134
rect 40144 43790 40172 44338
rect 41064 44266 41092 44814
rect 41052 44260 41104 44266
rect 41052 44202 41104 44208
rect 40316 44192 40368 44198
rect 40316 44134 40368 44140
rect 40328 43790 40356 44134
rect 41524 43994 41552 45222
rect 43996 44804 44048 44810
rect 43996 44746 44048 44752
rect 42156 44736 42208 44742
rect 42156 44678 42208 44684
rect 43168 44736 43220 44742
rect 43168 44678 43220 44684
rect 41972 44192 42024 44198
rect 41972 44134 42024 44140
rect 41512 43988 41564 43994
rect 41512 43930 41564 43936
rect 41984 43858 42012 44134
rect 41972 43852 42024 43858
rect 41972 43794 42024 43800
rect 42168 43790 42196 44678
rect 38752 43784 38804 43790
rect 38752 43726 38804 43732
rect 40132 43784 40184 43790
rect 40132 43726 40184 43732
rect 40316 43784 40368 43790
rect 40316 43726 40368 43732
rect 42156 43784 42208 43790
rect 42156 43726 42208 43732
rect 43180 43722 43208 44678
rect 43260 44192 43312 44198
rect 43260 44134 43312 44140
rect 43272 43790 43300 44134
rect 44008 43994 44036 44746
rect 44180 44328 44232 44334
rect 44180 44270 44232 44276
rect 43996 43988 44048 43994
rect 43996 43930 44048 43936
rect 43260 43784 43312 43790
rect 43260 43726 43312 43732
rect 43168 43716 43220 43722
rect 43168 43658 43220 43664
rect 43628 43716 43680 43722
rect 43628 43658 43680 43664
rect 40960 43648 41012 43654
rect 40960 43590 41012 43596
rect 42340 43648 42392 43654
rect 42340 43590 42392 43596
rect 38660 43444 38712 43450
rect 38660 43386 38712 43392
rect 40972 43382 41000 43590
rect 42352 43382 42380 43590
rect 43640 43450 43668 43658
rect 43628 43444 43680 43450
rect 43628 43386 43680 43392
rect 37740 43376 37792 43382
rect 37740 43318 37792 43324
rect 40960 43376 41012 43382
rect 40960 43318 41012 43324
rect 42340 43376 42392 43382
rect 42340 43318 42392 43324
rect 41328 43308 41380 43314
rect 41328 43250 41380 43256
rect 37280 43240 37332 43246
rect 37280 43182 37332 43188
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 33876 42696 33928 42702
rect 33876 42638 33928 42644
rect 35072 42696 35124 42702
rect 35072 42638 35124 42644
rect 32404 42288 32456 42294
rect 32404 42230 32456 42236
rect 29000 42084 29052 42090
rect 29000 42026 29052 42032
rect 27252 41812 27304 41818
rect 27252 41754 27304 41760
rect 29012 41682 29040 42026
rect 29000 41676 29052 41682
rect 29000 41618 29052 41624
rect 27068 41608 27120 41614
rect 27068 41550 27120 41556
rect 27436 41608 27488 41614
rect 27436 41550 27488 41556
rect 25780 41472 25832 41478
rect 25780 41414 25832 41420
rect 25792 41138 25820 41414
rect 25780 41132 25832 41138
rect 25780 41074 25832 41080
rect 25596 41064 25648 41070
rect 25596 41006 25648 41012
rect 25504 40928 25556 40934
rect 25504 40870 25556 40876
rect 25688 40928 25740 40934
rect 25688 40870 25740 40876
rect 25700 40526 25728 40870
rect 27080 40730 27108 41550
rect 27344 41540 27396 41546
rect 27344 41482 27396 41488
rect 27356 41274 27384 41482
rect 27344 41268 27396 41274
rect 27344 41210 27396 41216
rect 26332 40724 26384 40730
rect 26332 40666 26384 40672
rect 27068 40724 27120 40730
rect 27068 40666 27120 40672
rect 25688 40520 25740 40526
rect 25688 40462 25740 40468
rect 25228 40044 25280 40050
rect 25228 39986 25280 39992
rect 24216 39840 24268 39846
rect 24216 39782 24268 39788
rect 23572 39636 23624 39642
rect 23572 39578 23624 39584
rect 22468 39432 22520 39438
rect 22468 39374 22520 39380
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 13544 38548 13596 38554
rect 13544 38490 13596 38496
rect 13176 38412 13228 38418
rect 13176 38354 13228 38360
rect 11796 38344 11848 38350
rect 11796 38286 11848 38292
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 11704 38276 11756 38282
rect 11704 38218 11756 38224
rect 12544 37874 12572 38286
rect 13084 38276 13136 38282
rect 13084 38218 13136 38224
rect 13096 38010 13124 38218
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 12532 37868 12584 37874
rect 12532 37810 12584 37816
rect 13188 37466 13216 38354
rect 13912 38344 13964 38350
rect 13912 38286 13964 38292
rect 13924 38010 13952 38286
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 13912 38004 13964 38010
rect 13912 37946 13964 37952
rect 23308 37874 23336 38898
rect 23492 38554 23520 38898
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23584 37942 23612 38286
rect 23572 37936 23624 37942
rect 23572 37878 23624 37884
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 13176 37460 13228 37466
rect 13176 37402 13228 37408
rect 23308 37262 23336 37810
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 11888 37188 11940 37194
rect 11888 37130 11940 37136
rect 22928 37188 22980 37194
rect 22928 37130 22980 37136
rect 11900 36786 11928 37130
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 22940 36786 22968 37130
rect 11888 36780 11940 36786
rect 11888 36722 11940 36728
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23480 36712 23532 36718
rect 23480 36654 23532 36660
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 20088 34746 20116 35226
rect 21364 35080 21416 35086
rect 21416 35028 21588 35034
rect 21364 35022 21588 35028
rect 21376 35006 21588 35022
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 21560 34542 21588 35006
rect 22020 34678 22048 35430
rect 23492 35154 23520 36654
rect 23768 36378 23796 36722
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23584 35290 23612 35634
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23480 35148 23532 35154
rect 23480 35090 23532 35096
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23308 34746 23336 35022
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 22008 34672 22060 34678
rect 22008 34614 22060 34620
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21560 34066 21588 34478
rect 22296 34202 22324 34546
rect 23400 34202 23428 35022
rect 23492 34474 23520 35090
rect 23480 34468 23532 34474
rect 23480 34410 23532 34416
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 21548 34060 21600 34066
rect 21548 34002 21600 34008
rect 22008 33924 22060 33930
rect 22008 33866 22060 33872
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 22020 33522 22048 33866
rect 24228 33522 24256 39782
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24596 37466 24624 38694
rect 26240 38208 26292 38214
rect 26240 38150 26292 38156
rect 24676 37664 24728 37670
rect 24676 37606 24728 37612
rect 24584 37460 24636 37466
rect 24584 37402 24636 37408
rect 24688 37330 24716 37606
rect 24676 37324 24728 37330
rect 24676 37266 24728 37272
rect 24860 37256 24912 37262
rect 24860 37198 24912 37204
rect 24872 36922 24900 37198
rect 26252 37194 26280 38150
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 24860 36916 24912 36922
rect 24860 36858 24912 36864
rect 25608 35494 25636 37062
rect 26344 35834 26372 40666
rect 27448 40526 27476 41550
rect 27988 41268 28040 41274
rect 27988 41210 28040 41216
rect 28000 40526 28028 41210
rect 29012 41138 29040 41618
rect 28264 41132 28316 41138
rect 28264 41074 28316 41080
rect 29000 41132 29052 41138
rect 29000 41074 29052 41080
rect 30380 41132 30432 41138
rect 30380 41074 30432 41080
rect 27436 40520 27488 40526
rect 27436 40462 27488 40468
rect 27988 40520 28040 40526
rect 27988 40462 28040 40468
rect 27528 40452 27580 40458
rect 27528 40394 27580 40400
rect 26700 40384 26752 40390
rect 26700 40326 26752 40332
rect 26712 40118 26740 40326
rect 26700 40112 26752 40118
rect 26700 40054 26752 40060
rect 27540 39914 27568 40394
rect 27620 40044 27672 40050
rect 27620 39986 27672 39992
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 27528 39908 27580 39914
rect 27528 39850 27580 39856
rect 27540 39098 27568 39850
rect 27528 39092 27580 39098
rect 27528 39034 27580 39040
rect 27436 38956 27488 38962
rect 27436 38898 27488 38904
rect 27448 38350 27476 38898
rect 27632 38486 27660 39986
rect 27724 39030 27752 39986
rect 28000 39982 28028 40462
rect 28276 40186 28304 41074
rect 30104 40928 30156 40934
rect 30104 40870 30156 40876
rect 30116 40526 30144 40870
rect 29736 40520 29788 40526
rect 29736 40462 29788 40468
rect 30104 40520 30156 40526
rect 30104 40462 30156 40468
rect 28448 40384 28500 40390
rect 28448 40326 28500 40332
rect 28264 40180 28316 40186
rect 28264 40122 28316 40128
rect 28460 40050 28488 40326
rect 28448 40044 28500 40050
rect 28448 39986 28500 39992
rect 27988 39976 28040 39982
rect 27988 39918 28040 39924
rect 27712 39024 27764 39030
rect 27712 38966 27764 38972
rect 28172 38956 28224 38962
rect 28172 38898 28224 38904
rect 27712 38548 27764 38554
rect 27712 38490 27764 38496
rect 27620 38480 27672 38486
rect 27620 38422 27672 38428
rect 27436 38344 27488 38350
rect 27436 38286 27488 38292
rect 27068 37664 27120 37670
rect 27068 37606 27120 37612
rect 27080 36174 27108 37606
rect 27448 37466 27476 38286
rect 27528 37936 27580 37942
rect 27528 37878 27580 37884
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 27172 36786 27200 37062
rect 27540 36922 27568 37878
rect 27724 37670 27752 38490
rect 28184 38214 28212 38898
rect 28356 38888 28408 38894
rect 28356 38830 28408 38836
rect 28368 38350 28396 38830
rect 28460 38554 28488 39986
rect 28448 38548 28500 38554
rect 28448 38490 28500 38496
rect 28908 38548 28960 38554
rect 28908 38490 28960 38496
rect 28356 38344 28408 38350
rect 28356 38286 28408 38292
rect 28368 38214 28396 38286
rect 28172 38208 28224 38214
rect 28172 38150 28224 38156
rect 28356 38208 28408 38214
rect 28356 38150 28408 38156
rect 28184 37874 28212 38150
rect 28368 37874 28396 38150
rect 28172 37868 28224 37874
rect 28172 37810 28224 37816
rect 28356 37868 28408 37874
rect 28356 37810 28408 37816
rect 27712 37664 27764 37670
rect 27712 37606 27764 37612
rect 27804 37188 27856 37194
rect 27804 37130 27856 37136
rect 27528 36916 27580 36922
rect 27528 36858 27580 36864
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27264 36378 27292 36722
rect 27252 36372 27304 36378
rect 27252 36314 27304 36320
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 26332 35828 26384 35834
rect 26332 35770 26384 35776
rect 27068 35692 27120 35698
rect 27068 35634 27120 35640
rect 25596 35488 25648 35494
rect 25596 35430 25648 35436
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24596 34610 24624 35090
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 24584 34604 24636 34610
rect 24584 34546 24636 34552
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24596 34066 24624 34546
rect 24584 34060 24636 34066
rect 24584 34002 24636 34008
rect 24596 33658 24624 34002
rect 24872 33998 24900 34546
rect 26620 34202 26648 34886
rect 26700 34740 26752 34746
rect 26700 34682 26752 34688
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26712 34066 26740 34682
rect 27080 34202 27108 35634
rect 27068 34196 27120 34202
rect 27068 34138 27120 34144
rect 27816 34066 27844 37130
rect 28184 36854 28212 37810
rect 28368 37738 28396 37810
rect 28356 37732 28408 37738
rect 28356 37674 28408 37680
rect 28368 37466 28396 37674
rect 28816 37664 28868 37670
rect 28920 37652 28948 38490
rect 29644 38276 29696 38282
rect 29644 38218 29696 38224
rect 29656 37670 29684 38218
rect 28868 37624 28948 37652
rect 29644 37664 29696 37670
rect 28816 37606 28868 37612
rect 29644 37606 29696 37612
rect 28828 37466 28856 37606
rect 28356 37460 28408 37466
rect 28356 37402 28408 37408
rect 28816 37460 28868 37466
rect 28816 37402 28868 37408
rect 28172 36848 28224 36854
rect 28172 36790 28224 36796
rect 28368 36582 28396 37402
rect 29748 37262 29776 40462
rect 30392 40186 30420 41074
rect 31208 40384 31260 40390
rect 31208 40326 31260 40332
rect 30380 40180 30432 40186
rect 30380 40122 30432 40128
rect 31220 40050 31248 40326
rect 30564 40044 30616 40050
rect 30564 39986 30616 39992
rect 31208 40044 31260 40050
rect 31208 39986 31260 39992
rect 30576 38962 30604 39986
rect 30564 38956 30616 38962
rect 30564 38898 30616 38904
rect 30840 38956 30892 38962
rect 30840 38898 30892 38904
rect 30012 38208 30064 38214
rect 30012 38150 30064 38156
rect 29736 37256 29788 37262
rect 28644 37194 28948 37210
rect 29736 37198 29788 37204
rect 28632 37188 28960 37194
rect 28684 37182 28908 37188
rect 28632 37130 28684 37136
rect 28908 37130 28960 37136
rect 29748 36922 29776 37198
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 30024 35834 30052 38150
rect 30576 38010 30604 38898
rect 30748 38752 30800 38758
rect 30748 38694 30800 38700
rect 30760 38282 30788 38694
rect 30748 38276 30800 38282
rect 30748 38218 30800 38224
rect 30564 38004 30616 38010
rect 30564 37946 30616 37952
rect 30380 37868 30432 37874
rect 30380 37810 30432 37816
rect 30288 37732 30340 37738
rect 30288 37674 30340 37680
rect 30300 37262 30328 37674
rect 30288 37256 30340 37262
rect 30288 37198 30340 37204
rect 30300 36394 30328 37198
rect 30208 36378 30328 36394
rect 30196 36372 30328 36378
rect 30248 36366 30328 36372
rect 30196 36314 30248 36320
rect 30012 35828 30064 35834
rect 30012 35770 30064 35776
rect 30208 35698 30236 36314
rect 30392 35834 30420 37810
rect 30576 37482 30604 37946
rect 30852 37942 30880 38898
rect 31760 38480 31812 38486
rect 31760 38422 31812 38428
rect 30932 38208 30984 38214
rect 30932 38150 30984 38156
rect 30944 38010 30972 38150
rect 30932 38004 30984 38010
rect 30932 37946 30984 37952
rect 30840 37936 30892 37942
rect 30840 37878 30892 37884
rect 31116 37868 31168 37874
rect 31116 37810 31168 37816
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 30576 37466 30696 37482
rect 31128 37466 31156 37810
rect 30576 37460 30708 37466
rect 30576 37454 30656 37460
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 30576 35698 30604 37454
rect 30656 37402 30708 37408
rect 31116 37460 31168 37466
rect 31116 37402 31168 37408
rect 31496 37398 31524 37810
rect 31484 37392 31536 37398
rect 31484 37334 31536 37340
rect 31116 36916 31168 36922
rect 31116 36858 31168 36864
rect 31128 36242 31156 36858
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 28172 34400 28224 34406
rect 28172 34342 28224 34348
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 26700 34060 26752 34066
rect 26700 34002 26752 34008
rect 27804 34060 27856 34066
rect 27804 34002 27856 34008
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 26240 33924 26292 33930
rect 26240 33866 26292 33872
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 24216 33516 24268 33522
rect 24216 33458 24268 33464
rect 24596 32978 24624 33594
rect 26160 33454 26188 33866
rect 26148 33448 26200 33454
rect 26148 33390 26200 33396
rect 26252 33114 26280 33866
rect 28184 33590 28212 34342
rect 28828 33998 28856 34342
rect 31128 34082 31156 36178
rect 31772 36174 31800 38422
rect 31852 38208 31904 38214
rect 31852 38150 31904 38156
rect 31864 37942 31892 38150
rect 31852 37936 31904 37942
rect 31852 37878 31904 37884
rect 32312 37800 32364 37806
rect 32312 37742 32364 37748
rect 31852 37664 31904 37670
rect 31852 37606 31904 37612
rect 31864 37330 31892 37606
rect 31852 37324 31904 37330
rect 31852 37266 31904 37272
rect 32324 36922 32352 37742
rect 32416 36922 32444 42230
rect 33888 42226 33916 42638
rect 35084 42226 35112 42638
rect 33876 42220 33928 42226
rect 33876 42162 33928 42168
rect 35072 42220 35124 42226
rect 35072 42162 35124 42168
rect 37292 42158 37320 43182
rect 37372 42696 37424 42702
rect 37372 42638 37424 42644
rect 33324 42152 33376 42158
rect 33324 42094 33376 42100
rect 37280 42152 37332 42158
rect 37280 42094 37332 42100
rect 33336 41546 33364 42094
rect 34796 42016 34848 42022
rect 34796 41958 34848 41964
rect 35348 42016 35400 42022
rect 35348 41958 35400 41964
rect 34808 41682 34836 41958
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41818 35388 41958
rect 35348 41812 35400 41818
rect 35348 41754 35400 41760
rect 34796 41676 34848 41682
rect 34796 41618 34848 41624
rect 37188 41608 37240 41614
rect 37292 41562 37320 42094
rect 37384 41614 37412 42638
rect 38108 42560 38160 42566
rect 38108 42502 38160 42508
rect 38120 42294 38148 42502
rect 38108 42288 38160 42294
rect 38108 42230 38160 42236
rect 39212 42288 39264 42294
rect 39212 42230 39264 42236
rect 38568 42152 38620 42158
rect 38568 42094 38620 42100
rect 38580 41750 38608 42094
rect 38568 41744 38620 41750
rect 38568 41686 38620 41692
rect 38660 41676 38712 41682
rect 38660 41618 38712 41624
rect 37240 41556 37320 41562
rect 37188 41550 37320 41556
rect 37372 41608 37424 41614
rect 37372 41550 37424 41556
rect 33324 41540 33376 41546
rect 33324 41482 33376 41488
rect 35072 41540 35124 41546
rect 37200 41534 37320 41550
rect 35072 41482 35124 41488
rect 33336 41138 33364 41482
rect 34980 41472 35032 41478
rect 34980 41414 35032 41420
rect 34992 41138 35020 41414
rect 35084 41274 35112 41482
rect 35072 41268 35124 41274
rect 35072 41210 35124 41216
rect 33324 41132 33376 41138
rect 33324 41074 33376 41080
rect 33508 41132 33560 41138
rect 33508 41074 33560 41080
rect 34980 41132 35032 41138
rect 34980 41074 35032 41080
rect 33520 40730 33548 41074
rect 37292 41070 37320 41534
rect 37740 41132 37792 41138
rect 37740 41074 37792 41080
rect 37280 41064 37332 41070
rect 37280 41006 37332 41012
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 33508 40724 33560 40730
rect 33508 40666 33560 40672
rect 37292 40458 37320 41006
rect 37280 40452 37332 40458
rect 37280 40394 37332 40400
rect 37292 39982 37320 40394
rect 37280 39976 37332 39982
rect 37280 39918 37332 39924
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 36636 38752 36688 38758
rect 36636 38694 36688 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 36648 37874 36676 38694
rect 37292 38350 37320 39918
rect 37752 39642 37780 41074
rect 37740 39636 37792 39642
rect 37740 39578 37792 39584
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 37292 37874 37320 38286
rect 38292 38208 38344 38214
rect 38292 38150 38344 38156
rect 36636 37868 36688 37874
rect 36636 37810 36688 37816
rect 37280 37868 37332 37874
rect 37280 37810 37332 37816
rect 37740 37868 37792 37874
rect 37740 37810 37792 37816
rect 37464 37800 37516 37806
rect 37464 37742 37516 37748
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 37476 37262 37504 37742
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 37464 37256 37516 37262
rect 37464 37198 37516 37204
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32324 36242 32352 36858
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 32312 36236 32364 36242
rect 32312 36178 32364 36184
rect 32956 36236 33008 36242
rect 32956 36178 33008 36184
rect 31760 36168 31812 36174
rect 31760 36110 31812 36116
rect 32968 35698 32996 36178
rect 33244 36174 33272 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 36188 36242 36216 37198
rect 36636 37188 36688 37194
rect 36636 37130 36688 37136
rect 36648 36786 36676 37130
rect 37752 36786 37780 37810
rect 38200 37664 38252 37670
rect 38200 37606 38252 37612
rect 38212 37466 38240 37606
rect 38200 37460 38252 37466
rect 38200 37402 38252 37408
rect 38304 37330 38332 38150
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 38672 37126 38700 41618
rect 39120 41540 39172 41546
rect 39120 41482 39172 41488
rect 38752 41472 38804 41478
rect 38752 41414 38804 41420
rect 38764 40730 38792 41414
rect 39028 40928 39080 40934
rect 39028 40870 39080 40876
rect 38752 40724 38804 40730
rect 38752 40666 38804 40672
rect 39040 40526 39068 40870
rect 39132 40730 39160 41482
rect 39120 40724 39172 40730
rect 39120 40666 39172 40672
rect 39028 40520 39080 40526
rect 39028 40462 39080 40468
rect 38844 40452 38896 40458
rect 38844 40394 38896 40400
rect 38856 40186 38884 40394
rect 38844 40180 38896 40186
rect 38844 40122 38896 40128
rect 39224 38554 39252 42230
rect 39304 42084 39356 42090
rect 39304 42026 39356 42032
rect 39316 41614 39344 42026
rect 40684 42016 40736 42022
rect 40684 41958 40736 41964
rect 40696 41614 40724 41958
rect 41340 41818 41368 43250
rect 44008 43246 44036 43930
rect 44192 43450 44220 44270
rect 44284 43790 44312 45426
rect 44364 45008 44416 45014
rect 44364 44950 44416 44956
rect 44376 44266 44404 44950
rect 44364 44260 44416 44266
rect 44364 44202 44416 44208
rect 44272 43784 44324 43790
rect 44272 43726 44324 43732
rect 44180 43444 44232 43450
rect 44180 43386 44232 43392
rect 43996 43240 44048 43246
rect 43996 43182 44048 43188
rect 42616 43172 42668 43178
rect 42616 43114 42668 43120
rect 41328 41812 41380 41818
rect 41328 41754 41380 41760
rect 39304 41608 39356 41614
rect 39304 41550 39356 41556
rect 40684 41608 40736 41614
rect 40684 41550 40736 41556
rect 42156 41472 42208 41478
rect 42156 41414 42208 41420
rect 41328 41132 41380 41138
rect 41328 41074 41380 41080
rect 40316 41064 40368 41070
rect 40316 41006 40368 41012
rect 40132 40928 40184 40934
rect 40132 40870 40184 40876
rect 40144 40118 40172 40870
rect 40328 40526 40356 41006
rect 40316 40520 40368 40526
rect 40316 40462 40368 40468
rect 40132 40112 40184 40118
rect 40132 40054 40184 40060
rect 40328 39982 40356 40462
rect 40592 40452 40644 40458
rect 40592 40394 40644 40400
rect 40316 39976 40368 39982
rect 40316 39918 40368 39924
rect 40604 39642 40632 40394
rect 40684 39840 40736 39846
rect 40684 39782 40736 39788
rect 40592 39636 40644 39642
rect 40592 39578 40644 39584
rect 39212 38548 39264 38554
rect 39212 38490 39264 38496
rect 39224 37942 39252 38490
rect 40696 38350 40724 39782
rect 41340 39642 41368 41074
rect 42168 40730 42196 41414
rect 42432 40928 42484 40934
rect 42432 40870 42484 40876
rect 42156 40724 42208 40730
rect 42156 40666 42208 40672
rect 42444 40526 42472 40870
rect 42628 40730 42656 43114
rect 44008 42702 44036 43182
rect 44192 42702 44220 43386
rect 44376 43110 44404 44202
rect 44364 43104 44416 43110
rect 44364 43046 44416 43052
rect 43996 42696 44048 42702
rect 43996 42638 44048 42644
rect 44180 42696 44232 42702
rect 44180 42638 44232 42644
rect 44364 42696 44416 42702
rect 44364 42638 44416 42644
rect 44008 42226 44036 42638
rect 44180 42288 44232 42294
rect 44180 42230 44232 42236
rect 43996 42220 44048 42226
rect 43996 42162 44048 42168
rect 43444 42016 43496 42022
rect 43444 41958 43496 41964
rect 43456 41546 43484 41958
rect 43444 41540 43496 41546
rect 43444 41482 43496 41488
rect 44192 41274 44220 42230
rect 44376 42226 44404 42638
rect 44364 42220 44416 42226
rect 44364 42162 44416 42168
rect 44180 41268 44232 41274
rect 44180 41210 44232 41216
rect 42616 40724 42668 40730
rect 42616 40666 42668 40672
rect 41788 40520 41840 40526
rect 41788 40462 41840 40468
rect 42432 40520 42484 40526
rect 42432 40462 42484 40468
rect 41800 40186 41828 40462
rect 41788 40180 41840 40186
rect 41788 40122 41840 40128
rect 41328 39636 41380 39642
rect 41328 39578 41380 39584
rect 40776 38956 40828 38962
rect 40776 38898 40828 38904
rect 41604 38956 41656 38962
rect 41604 38898 41656 38904
rect 40132 38344 40184 38350
rect 40132 38286 40184 38292
rect 40684 38344 40736 38350
rect 40684 38286 40736 38292
rect 39212 37936 39264 37942
rect 39212 37878 39264 37884
rect 39396 37936 39448 37942
rect 39396 37878 39448 37884
rect 38844 37664 38896 37670
rect 38844 37606 38896 37612
rect 38856 37262 38884 37606
rect 38844 37256 38896 37262
rect 38844 37198 38896 37204
rect 39304 37256 39356 37262
rect 39304 37198 39356 37204
rect 38660 37120 38712 37126
rect 38660 37062 38712 37068
rect 36636 36780 36688 36786
rect 36636 36722 36688 36728
rect 37740 36780 37792 36786
rect 37740 36722 37792 36728
rect 39316 36650 39344 37198
rect 39304 36644 39356 36650
rect 39304 36586 39356 36592
rect 36176 36236 36228 36242
rect 36176 36178 36228 36184
rect 33232 36168 33284 36174
rect 33232 36110 33284 36116
rect 38108 36100 38160 36106
rect 38108 36042 38160 36048
rect 34796 36032 34848 36038
rect 34796 35974 34848 35980
rect 37648 36032 37700 36038
rect 37648 35974 37700 35980
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32968 35154 32996 35634
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 34520 35488 34572 35494
rect 34520 35430 34572 35436
rect 32956 35148 33008 35154
rect 32956 35090 33008 35096
rect 34440 35086 34468 35430
rect 34532 35154 34560 35430
rect 34808 35290 34836 35974
rect 36544 35488 36596 35494
rect 36544 35430 36596 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 35284 34848 35290
rect 34796 35226 34848 35232
rect 34520 35148 34572 35154
rect 34520 35090 34572 35096
rect 36556 35086 36584 35430
rect 34428 35080 34480 35086
rect 34428 35022 34480 35028
rect 35164 35080 35216 35086
rect 35164 35022 35216 35028
rect 36268 35080 36320 35086
rect 36268 35022 36320 35028
rect 36544 35080 36596 35086
rect 36544 35022 36596 35028
rect 35176 34746 35204 35022
rect 35164 34740 35216 34746
rect 35164 34682 35216 34688
rect 33876 34604 33928 34610
rect 33876 34546 33928 34552
rect 32312 34468 32364 34474
rect 32312 34410 32364 34416
rect 31208 34400 31260 34406
rect 31208 34342 31260 34348
rect 31036 34054 31156 34082
rect 31036 33998 31064 34054
rect 31220 33998 31248 34342
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 31024 33992 31076 33998
rect 31024 33934 31076 33940
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 29736 33856 29788 33862
rect 29736 33798 29788 33804
rect 28172 33584 28224 33590
rect 28172 33526 28224 33532
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26436 33114 26464 33458
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26424 33108 26476 33114
rect 26424 33050 26476 33056
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 23308 31346 23336 32914
rect 24596 31890 24624 32914
rect 27816 32910 27844 33390
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 29276 33312 29328 33318
rect 29276 33254 29328 33260
rect 27908 32910 27936 33254
rect 29288 32910 29316 33254
rect 29748 33114 29776 33798
rect 30484 33658 30512 33934
rect 30472 33652 30524 33658
rect 30472 33594 30524 33600
rect 31036 33590 31064 33934
rect 31760 33924 31812 33930
rect 31760 33866 31812 33872
rect 31772 33658 31800 33866
rect 31760 33652 31812 33658
rect 31760 33594 31812 33600
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 30932 33516 30984 33522
rect 30932 33458 30984 33464
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 29276 32904 29328 32910
rect 29276 32846 29328 32852
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 24872 32434 24900 32778
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 27620 32224 27672 32230
rect 27620 32166 27672 32172
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 27632 31822 27660 32166
rect 27816 32026 27844 32846
rect 28908 32836 28960 32842
rect 28908 32778 28960 32784
rect 28920 32026 28948 32778
rect 30944 32434 30972 33458
rect 32324 33454 32352 34410
rect 33888 34202 33916 34546
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 33048 34196 33100 34202
rect 33048 34138 33100 34144
rect 33876 34196 33928 34202
rect 33876 34138 33928 34144
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 32312 33448 32364 33454
rect 32312 33390 32364 33396
rect 31392 33312 31444 33318
rect 31392 33254 31444 33260
rect 31116 32904 31168 32910
rect 31116 32846 31168 32852
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 27804 32020 27856 32026
rect 27804 31962 27856 31968
rect 28908 32020 28960 32026
rect 28908 31962 28960 31968
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 23308 30190 23336 31282
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23584 30326 23612 30670
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 22848 29238 22876 29990
rect 23308 29646 23336 30126
rect 24596 29714 24624 31078
rect 25148 30258 25176 31282
rect 30840 31136 30892 31142
rect 30840 31078 30892 31084
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30392 30258 30420 30670
rect 30852 30666 30880 31078
rect 31128 30734 31156 32846
rect 31404 32842 31432 33254
rect 32324 32910 32352 33390
rect 32508 33114 32536 33934
rect 33060 33658 33088 34138
rect 36280 33998 36308 35022
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 37476 34678 37504 34886
rect 37464 34672 37516 34678
rect 37464 34614 37516 34620
rect 37556 34536 37608 34542
rect 37556 34478 37608 34484
rect 36452 34400 36504 34406
rect 36452 34342 36504 34348
rect 36268 33992 36320 33998
rect 36268 33934 36320 33940
rect 36464 33930 36492 34342
rect 37568 34202 37596 34478
rect 37660 34406 37688 35974
rect 38120 35290 38148 36042
rect 38108 35284 38160 35290
rect 38108 35226 38160 35232
rect 37740 34944 37792 34950
rect 37740 34886 37792 34892
rect 37752 34610 37780 34886
rect 37740 34604 37792 34610
rect 37740 34546 37792 34552
rect 39304 34536 39356 34542
rect 39304 34478 39356 34484
rect 37648 34400 37700 34406
rect 37648 34342 37700 34348
rect 38016 34400 38068 34406
rect 38016 34342 38068 34348
rect 37556 34196 37608 34202
rect 37556 34138 37608 34144
rect 38028 33998 38056 34342
rect 39316 34202 39344 34478
rect 39304 34196 39356 34202
rect 39304 34138 39356 34144
rect 38016 33992 38068 33998
rect 38016 33934 38068 33940
rect 38200 33992 38252 33998
rect 38200 33934 38252 33940
rect 36452 33924 36504 33930
rect 36452 33866 36504 33872
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 33244 33114 33272 33798
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 38212 33114 38240 33934
rect 38384 33924 38436 33930
rect 38384 33866 38436 33872
rect 38396 33454 38424 33866
rect 39304 33856 39356 33862
rect 39304 33798 39356 33804
rect 39316 33658 39344 33798
rect 39304 33652 39356 33658
rect 39304 33594 39356 33600
rect 39212 33516 39264 33522
rect 39212 33458 39264 33464
rect 38384 33448 38436 33454
rect 38384 33390 38436 33396
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 33232 33108 33284 33114
rect 33232 33050 33284 33056
rect 38200 33108 38252 33114
rect 38200 33050 38252 33056
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 31392 32836 31444 32842
rect 31392 32778 31444 32784
rect 32496 31408 32548 31414
rect 32496 31350 32548 31356
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 30840 30660 30892 30666
rect 30840 30602 30892 30608
rect 31404 30394 31432 30670
rect 31392 30388 31444 30394
rect 31392 30330 31444 30336
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24688 29850 24716 29990
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 22836 29232 22888 29238
rect 22836 29174 22888 29180
rect 23308 29170 23336 29582
rect 24872 29306 24900 29582
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 17328 28558 17356 28902
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 16960 28014 16988 28494
rect 18340 28150 18368 28902
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 20088 28082 20116 28358
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 16948 28008 17000 28014
rect 16948 27950 17000 27956
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16776 27062 16804 27814
rect 16960 27470 16988 27950
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17328 27470 17356 27814
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16960 26994 16988 27406
rect 19352 27130 19380 28018
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 20352 27872 20404 27878
rect 20352 27814 20404 27820
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 19904 27606 19932 27814
rect 19892 27600 19944 27606
rect 19892 27542 19944 27548
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13372 25974 13400 26182
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13556 25498 13584 26318
rect 16960 26234 16988 26930
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 16960 26206 17080 26234
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13452 25424 13504 25430
rect 13452 25366 13504 25372
rect 13464 24954 13492 25366
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12084 23730 12112 24142
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23798 12296 24074
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 12084 23050 12112 23666
rect 12268 23322 12296 23734
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 12360 23118 12388 24006
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22710 2912 22918
rect 12084 22778 12112 22986
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 13004 22710 13032 24550
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 2964 22568 3016 22574
rect 1766 22536 1822 22545
rect 2964 22510 3016 22516
rect 1766 22471 1822 22480
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22030 1624 22374
rect 1780 22234 1808 22471
rect 1768 22228 1820 22234
rect 1768 22170 1820 22176
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2136 20868 2188 20874
rect 2136 20810 2188 20816
rect 2148 20466 2176 20810
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2332 19854 2360 21286
rect 2608 20942 2636 21626
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2608 20466 2636 20878
rect 2884 20534 2912 22102
rect 2976 21690 3004 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 13188 21894 13216 24754
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 22030 13308 24006
rect 13372 22234 13400 24550
rect 13464 24342 13492 24890
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13464 21962 13492 24278
rect 13556 24206 13584 24754
rect 13832 24206 13860 25638
rect 14016 25294 14044 25638
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 13912 25220 13964 25226
rect 13912 25162 13964 25168
rect 13924 24818 13952 25162
rect 14016 24886 14044 25230
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 14568 24954 14596 25094
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 15856 24886 15884 25774
rect 17052 25294 17080 26206
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17328 25294 17356 25638
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17052 24886 17080 25230
rect 14004 24880 14056 24886
rect 14004 24822 14056 24828
rect 15844 24880 15896 24886
rect 15844 24822 15896 24828
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13832 23186 13860 24142
rect 13924 24138 13952 24754
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 14016 24070 14044 24822
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14464 24064 14516 24070
rect 14648 24064 14700 24070
rect 14516 24012 14596 24018
rect 14464 24006 14596 24012
rect 14648 24006 14700 24012
rect 14476 23990 14596 24006
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13832 22778 13860 23122
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13832 22642 13860 22714
rect 14016 22642 14044 23462
rect 14568 23118 14596 23990
rect 14660 23186 14688 24006
rect 15212 23730 15240 24550
rect 15396 24138 15424 24550
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15856 23730 15884 24822
rect 17052 24274 17080 24822
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17144 24206 17172 24550
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 16040 23730 16068 24142
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16224 23798 16252 24074
rect 16868 23798 16896 24142
rect 16212 23792 16264 23798
rect 16212 23734 16264 23740
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 15212 23050 15240 23462
rect 15488 23254 15516 23666
rect 15672 23322 15700 23666
rect 16224 23322 16252 23734
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 4632 21554 4660 21830
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 3436 20058 3464 20810
rect 3988 20602 4016 21082
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4264 20602 4292 20878
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 2056 18834 2084 19790
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18290 2084 18770
rect 2332 18766 2360 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3528 18426 3556 18634
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2056 17746 2084 18226
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 2056 17202 2084 17682
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2240 17134 2268 18226
rect 3896 17882 3924 18770
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 18170 4200 18702
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4080 18142 4200 18170
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17678 4016 18022
rect 4080 17864 4108 18142
rect 4448 18086 4476 18566
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4080 17836 4200 17864
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4172 17338 4200 17836
rect 4632 17678 4660 21490
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4724 18358 4752 20742
rect 5552 20534 5580 21286
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5828 19378 5856 20334
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 19786 12756 20198
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 13648 19378 13676 20878
rect 13832 20534 13860 22578
rect 14016 21554 14044 22578
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21554 14412 21830
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13832 19922 13860 20470
rect 13924 20466 13952 20878
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13832 19446 13860 19858
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4816 18290 4844 18566
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4632 17202 4660 17478
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 3988 16794 4016 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15094 4660 17138
rect 5092 16574 5120 18022
rect 5644 17270 5672 18702
rect 6564 18290 6592 19314
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18970 7972 19110
rect 14568 18970 14596 19722
rect 14752 19514 14780 20334
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14844 19378 14872 21490
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 20534 16620 21286
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15212 20058 15240 20402
rect 15672 20058 15700 20402
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 16684 19786 16712 22374
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16764 20936 16816 20942
rect 16960 20924 16988 21490
rect 16816 20896 16988 20924
rect 16764 20878 16816 20884
rect 16960 20466 16988 20896
rect 17052 20874 17080 21966
rect 17604 21622 17632 21966
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16960 19786 16988 20402
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 7024 17882 7052 18702
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 6564 16998 6592 17614
rect 7116 17610 7144 18294
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 5092 16546 5212 16574
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3620 14618 3648 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13938 4292 14214
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4540 13818 4568 14350
rect 4632 14006 4660 15030
rect 4712 14408 4764 14414
rect 4896 14408 4948 14414
rect 4764 14368 4844 14396
rect 4712 14350 4764 14356
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4816 13938 4844 14368
rect 4896 14350 4948 14356
rect 4908 14074 4936 14350
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4540 13790 4660 13818
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 12986 4660 13790
rect 4816 13326 4844 13874
rect 4908 13326 4936 14010
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4816 12850 4844 13262
rect 4908 12850 4936 13262
rect 5184 13258 5212 16546
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14074 5580 14350
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5644 13954 5672 14758
rect 5552 13938 5672 13954
rect 5540 13932 5672 13938
rect 5592 13926 5672 13932
rect 5540 13874 5592 13880
rect 5552 13394 5580 13874
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11082 2268 11494
rect 2700 11150 2728 11630
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2700 10674 2728 11086
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10266 2728 10610
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 2446 1900 9862
rect 2792 9586 2820 10542
rect 3344 10062 3372 10950
rect 3988 10674 4016 12174
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 10742 4384 11018
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10266 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 10542
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4724 10130 4752 11562
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4816 10062 4844 10406
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 5000 9994 5028 13126
rect 5184 12986 5212 13194
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5644 12850 5672 13398
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11218 5488 12174
rect 6564 11898 6592 16934
rect 7116 15026 7144 17546
rect 7392 17066 7420 18634
rect 7944 18426 7972 18702
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8404 17610 8432 18022
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 14660 17270 14688 17614
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14108 16114 14136 16458
rect 14200 16182 14228 16594
rect 14292 16590 14320 17070
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14618 7420 14962
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7668 14414 7696 15302
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 8036 14074 8064 15370
rect 8220 14482 8248 15642
rect 8956 15502 8984 15846
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15162 8984 15302
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8588 14482 8616 14826
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8128 13938 8156 14214
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6564 11234 6592 11834
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 6472 11206 6592 11234
rect 5460 10742 5488 11154
rect 6472 11150 6500 11206
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5460 10130 5488 10678
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5736 10062 5764 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5828 9586 5856 11018
rect 6656 10810 6684 13262
rect 8036 13258 8064 13806
rect 8128 13326 8156 13874
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12850 8064 13194
rect 8128 12986 8156 13262
rect 8220 13190 8248 14418
rect 8864 14074 8892 14554
rect 9140 14550 9168 16050
rect 14292 16046 14320 16526
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 15094 9352 15302
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9324 14906 9352 15030
rect 9232 14878 9352 14906
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9232 14482 9260 14878
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 9232 13938 9260 14418
rect 9324 14346 9352 14758
rect 10520 14346 10548 15438
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7392 12646 7420 12786
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7760 12434 7788 12582
rect 7668 12406 7788 12434
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11762 7144 12038
rect 7300 11898 7328 12106
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6932 10674 6960 10950
rect 7668 10674 7696 12406
rect 8220 12374 8248 13126
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11762 7788 12174
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8220 10470 8248 12310
rect 8404 12170 8432 13126
rect 8588 12850 8616 13262
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8588 12442 8616 12786
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 9048 11898 9076 12854
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 12374 9444 12650
rect 9600 12646 9628 14282
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9508 10742 9536 12582
rect 9600 12442 9628 12582
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 10520 12238 10548 14282
rect 10980 14006 11008 14962
rect 11164 14074 11192 15030
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10980 13190 11008 13942
rect 11256 13938 11284 14214
rect 11348 14006 11376 14350
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11256 13802 11284 13874
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10796 12238 10824 13126
rect 10980 12850 11008 13126
rect 11072 12986 11100 13262
rect 11348 13258 11376 13942
rect 11716 13734 11744 14758
rect 11808 14618 11836 15030
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11808 14278 11836 14418
rect 13096 14414 13124 14758
rect 13740 14414 13768 14826
rect 14568 14822 14596 15982
rect 14844 15026 14872 19314
rect 16856 18760 16908 18766
rect 16960 18714 16988 19722
rect 17972 19378 18000 26250
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20364 25906 20392 27814
rect 21008 27470 21036 27814
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 20640 26926 20668 27406
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20640 26586 20668 26862
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23662 18736 24006
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18892 23526 18920 25094
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19168 23730 19196 24550
rect 19352 23866 19380 25774
rect 20640 25362 20668 26522
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20364 24818 20392 25230
rect 20640 24886 20668 25298
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 21008 24138 21036 25638
rect 21100 25294 21128 25638
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 22020 24954 22048 25842
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22112 24410 22140 25774
rect 22204 25498 22232 25842
rect 22296 25702 22324 27270
rect 23216 27062 23244 27406
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24596 26450 24624 26862
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 23112 26308 23164 26314
rect 23112 26250 23164 26256
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 23124 24818 23152 26250
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 24596 24682 24624 26386
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 24596 24274 24624 24618
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 20996 24132 21048 24138
rect 20996 24074 21048 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 23032 23050 23060 24142
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23308 23730 23336 24006
rect 24044 23730 24072 24142
rect 24596 23798 24624 24210
rect 24688 24138 24716 27814
rect 24872 26382 24900 28494
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24964 25974 24992 26726
rect 24952 25968 25004 25974
rect 24952 25910 25004 25916
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24872 25702 24900 25842
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 24596 23186 24624 23734
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 24872 23118 24900 25230
rect 24964 23866 24992 25774
rect 25056 25702 25084 27270
rect 25148 25906 25176 29446
rect 30300 29170 30328 29582
rect 30392 29238 30420 30194
rect 31404 29714 31432 30330
rect 31496 30326 31524 31078
rect 31760 30796 31812 30802
rect 31760 30738 31812 30744
rect 31484 30320 31536 30326
rect 31484 30262 31536 30268
rect 31772 30122 31800 30738
rect 32404 30660 32456 30666
rect 32404 30602 32456 30608
rect 31760 30116 31812 30122
rect 31760 30058 31812 30064
rect 31944 30048 31996 30054
rect 31944 29990 31996 29996
rect 31392 29708 31444 29714
rect 31392 29650 31444 29656
rect 31956 29646 31984 29990
rect 31944 29640 31996 29646
rect 31944 29582 31996 29588
rect 32416 29306 32444 30602
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 30380 29232 30432 29238
rect 30380 29174 30432 29180
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 32508 28762 32536 31350
rect 33152 30938 33180 32846
rect 33244 32570 33272 32846
rect 33232 32564 33284 32570
rect 33232 32506 33284 32512
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 34716 31346 34744 31758
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34808 31278 34836 31758
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 33140 30932 33192 30938
rect 33140 30874 33192 30880
rect 34808 30734 34836 31214
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 32680 30728 32732 30734
rect 32680 30670 32732 30676
rect 34796 30728 34848 30734
rect 34796 30670 34848 30676
rect 32692 29850 32720 30670
rect 34808 30394 34836 30670
rect 35360 30666 35388 32166
rect 35452 31822 35480 32846
rect 36912 32496 36964 32502
rect 36912 32438 36964 32444
rect 35808 32428 35860 32434
rect 35808 32370 35860 32376
rect 36452 32428 36504 32434
rect 36452 32370 36504 32376
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35348 30660 35400 30666
rect 35348 30602 35400 30608
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 32680 29844 32732 29850
rect 32680 29786 32732 29792
rect 31760 28756 31812 28762
rect 31760 28698 31812 28704
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 30656 28416 30708 28422
rect 30656 28358 30708 28364
rect 30668 27946 30696 28358
rect 30656 27940 30708 27946
rect 30656 27882 30708 27888
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 25608 27062 25636 27814
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27344 27396 27396 27402
rect 27344 27338 27396 27344
rect 25596 27056 25648 27062
rect 25596 26998 25648 27004
rect 25320 26784 25372 26790
rect 25320 26726 25372 26732
rect 25228 26240 25280 26246
rect 25228 26182 25280 26188
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25240 25838 25268 26182
rect 25332 25906 25360 26726
rect 27356 26586 27384 27338
rect 27724 26994 27752 27406
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 27724 26450 27752 26930
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27724 25974 27752 26386
rect 27712 25968 27764 25974
rect 27712 25910 27764 25916
rect 27908 25906 27936 26726
rect 28644 26382 28672 27814
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 29104 25906 29132 27270
rect 31220 27130 31248 27406
rect 31208 27124 31260 27130
rect 31208 27066 31260 27072
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 29092 25900 29144 25906
rect 29092 25842 29144 25848
rect 29840 25838 29868 26726
rect 31772 26382 31800 28698
rect 34808 28558 34836 30330
rect 35820 30054 35848 32370
rect 35992 32360 36044 32366
rect 35992 32302 36044 32308
rect 36004 30938 36032 32302
rect 36084 32224 36136 32230
rect 36084 32166 36136 32172
rect 36096 32026 36124 32166
rect 36084 32020 36136 32026
rect 36084 31962 36136 31968
rect 36464 31482 36492 32370
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36452 31476 36504 31482
rect 36452 31418 36504 31424
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 36740 30326 36768 31758
rect 36924 31414 36952 32438
rect 38396 32230 38424 33390
rect 39224 33114 39252 33458
rect 39212 33108 39264 33114
rect 39212 33050 39264 33056
rect 39408 32502 39436 37878
rect 40040 37664 40092 37670
rect 40040 37606 40092 37612
rect 40052 37330 40080 37606
rect 40040 37324 40092 37330
rect 40040 37266 40092 37272
rect 39488 36780 39540 36786
rect 39488 36722 39540 36728
rect 39500 34202 39528 36722
rect 40052 35494 40080 37266
rect 40144 36922 40172 38286
rect 40316 38208 40368 38214
rect 40316 38150 40368 38156
rect 40224 37460 40276 37466
rect 40224 37402 40276 37408
rect 40132 36916 40184 36922
rect 40132 36858 40184 36864
rect 40236 36106 40264 37402
rect 40328 37262 40356 38150
rect 40696 37670 40724 38286
rect 40684 37664 40736 37670
rect 40684 37606 40736 37612
rect 40316 37256 40368 37262
rect 40316 37198 40368 37204
rect 40316 36916 40368 36922
rect 40316 36858 40368 36864
rect 40328 36378 40356 36858
rect 40788 36650 40816 38898
rect 41616 38214 41644 38898
rect 41972 38752 42024 38758
rect 41972 38694 42024 38700
rect 41604 38208 41656 38214
rect 41604 38150 41656 38156
rect 41616 37806 41644 38150
rect 41604 37800 41656 37806
rect 41604 37742 41656 37748
rect 41616 37194 41644 37742
rect 41880 37732 41932 37738
rect 41880 37674 41932 37680
rect 41892 37194 41920 37674
rect 41984 37194 42012 38694
rect 44468 38554 44496 45426
rect 45572 45354 45600 49166
rect 46584 46170 46612 57394
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 58256 49088 58308 49094
rect 58254 49056 58256 49065
rect 58308 49056 58310 49065
rect 50294 48988 50602 48997
rect 58254 48991 58310 49000
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 46572 46164 46624 46170
rect 46572 46106 46624 46112
rect 45836 45892 45888 45898
rect 45836 45834 45888 45840
rect 45560 45348 45612 45354
rect 45560 45290 45612 45296
rect 45848 45082 45876 45834
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 45836 45076 45888 45082
rect 45836 45018 45888 45024
rect 45468 44872 45520 44878
rect 45468 44814 45520 44820
rect 45192 44736 45244 44742
rect 45192 44678 45244 44684
rect 44548 44396 44600 44402
rect 44548 44338 44600 44344
rect 42800 38548 42852 38554
rect 42800 38490 42852 38496
rect 44456 38548 44508 38554
rect 44456 38490 44508 38496
rect 42064 38344 42116 38350
rect 42064 38286 42116 38292
rect 42076 38010 42104 38286
rect 42708 38276 42760 38282
rect 42708 38218 42760 38224
rect 42064 38004 42116 38010
rect 42064 37946 42116 37952
rect 42720 37466 42748 38218
rect 42812 37942 42840 38490
rect 44560 37942 44588 44338
rect 45008 43784 45060 43790
rect 45008 43726 45060 43732
rect 44824 43648 44876 43654
rect 44824 43590 44876 43596
rect 44836 42906 44864 43590
rect 45020 43314 45048 43726
rect 45204 43382 45232 44678
rect 45480 44538 45508 44814
rect 45560 44804 45612 44810
rect 45560 44746 45612 44752
rect 45468 44532 45520 44538
rect 45468 44474 45520 44480
rect 45376 44260 45428 44266
rect 45376 44202 45428 44208
rect 45388 43994 45416 44202
rect 45572 43994 45600 44746
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 45376 43988 45428 43994
rect 45376 43930 45428 43936
rect 45560 43988 45612 43994
rect 45560 43930 45612 43936
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 45192 43376 45244 43382
rect 45192 43318 45244 43324
rect 45008 43308 45060 43314
rect 45008 43250 45060 43256
rect 44824 42900 44876 42906
rect 44824 42842 44876 42848
rect 44640 42084 44692 42090
rect 44640 42026 44692 42032
rect 44652 41818 44680 42026
rect 44640 41812 44692 41818
rect 44640 41754 44692 41760
rect 45020 41478 45048 43250
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 45100 42016 45152 42022
rect 45100 41958 45152 41964
rect 45008 41472 45060 41478
rect 45008 41414 45060 41420
rect 45020 41138 45048 41414
rect 45112 41206 45140 41958
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 45100 41200 45152 41206
rect 45100 41142 45152 41148
rect 45008 41132 45060 41138
rect 45008 41074 45060 41080
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 42800 37936 42852 37942
rect 42800 37878 42852 37884
rect 44548 37936 44600 37942
rect 44548 37878 44600 37884
rect 42708 37460 42760 37466
rect 42708 37402 42760 37408
rect 41604 37188 41656 37194
rect 41604 37130 41656 37136
rect 41880 37188 41932 37194
rect 41880 37130 41932 37136
rect 41972 37188 42024 37194
rect 41972 37130 42024 37136
rect 41420 37120 41472 37126
rect 41420 37062 41472 37068
rect 41432 36786 41460 37062
rect 41892 36922 41920 37130
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 41880 36916 41932 36922
rect 41880 36858 41932 36864
rect 41420 36780 41472 36786
rect 41420 36722 41472 36728
rect 40776 36644 40828 36650
rect 40776 36586 40828 36592
rect 40316 36372 40368 36378
rect 40316 36314 40368 36320
rect 40224 36100 40276 36106
rect 40224 36042 40276 36048
rect 40132 36032 40184 36038
rect 40132 35974 40184 35980
rect 40040 35488 40092 35494
rect 40040 35430 40092 35436
rect 40144 35086 40172 35974
rect 40224 35760 40276 35766
rect 40224 35702 40276 35708
rect 40236 35290 40264 35702
rect 40224 35284 40276 35290
rect 40224 35226 40276 35232
rect 40132 35080 40184 35086
rect 40132 35022 40184 35028
rect 39764 34604 39816 34610
rect 39764 34546 39816 34552
rect 39948 34604 40000 34610
rect 39948 34546 40000 34552
rect 39488 34196 39540 34202
rect 39488 34138 39540 34144
rect 39776 34066 39804 34546
rect 39856 34536 39908 34542
rect 39856 34478 39908 34484
rect 39764 34060 39816 34066
rect 39764 34002 39816 34008
rect 39396 32496 39448 32502
rect 39396 32438 39448 32444
rect 39868 32434 39896 34478
rect 39960 33658 39988 34546
rect 40224 34400 40276 34406
rect 40224 34342 40276 34348
rect 40236 34202 40264 34342
rect 40224 34196 40276 34202
rect 40224 34138 40276 34144
rect 40328 33998 40356 36314
rect 41144 36168 41196 36174
rect 41144 36110 41196 36116
rect 41156 35834 41184 36110
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 41144 35828 41196 35834
rect 41144 35770 41196 35776
rect 40500 35488 40552 35494
rect 40500 35430 40552 35436
rect 40316 33992 40368 33998
rect 40316 33934 40368 33940
rect 40132 33924 40184 33930
rect 40132 33866 40184 33872
rect 40040 33856 40092 33862
rect 40040 33798 40092 33804
rect 39948 33652 40000 33658
rect 39948 33594 40000 33600
rect 40052 32978 40080 33798
rect 40040 32972 40092 32978
rect 40040 32914 40092 32920
rect 40144 32842 40172 33866
rect 40316 33856 40368 33862
rect 40316 33798 40368 33804
rect 40328 33114 40356 33798
rect 40512 33522 40540 35430
rect 41156 34626 41184 35770
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 41064 34598 41184 34626
rect 41064 34542 41092 34598
rect 41052 34536 41104 34542
rect 41052 34478 41104 34484
rect 41064 33998 41092 34478
rect 41052 33992 41104 33998
rect 41052 33934 41104 33940
rect 41236 33992 41288 33998
rect 41236 33934 41288 33940
rect 43444 33992 43496 33998
rect 43444 33934 43496 33940
rect 41248 33658 41276 33934
rect 43260 33856 43312 33862
rect 43260 33798 43312 33804
rect 41236 33652 41288 33658
rect 41236 33594 41288 33600
rect 40500 33516 40552 33522
rect 40500 33458 40552 33464
rect 40776 33516 40828 33522
rect 40776 33458 40828 33464
rect 40788 33114 40816 33458
rect 40316 33108 40368 33114
rect 40316 33050 40368 33056
rect 40776 33108 40828 33114
rect 40776 33050 40828 33056
rect 40132 32836 40184 32842
rect 40132 32778 40184 32784
rect 40224 32768 40276 32774
rect 40224 32710 40276 32716
rect 41144 32768 41196 32774
rect 41144 32710 41196 32716
rect 40236 32570 40264 32710
rect 40224 32564 40276 32570
rect 40224 32506 40276 32512
rect 41156 32434 41184 32710
rect 39856 32428 39908 32434
rect 39856 32370 39908 32376
rect 41144 32428 41196 32434
rect 41144 32370 41196 32376
rect 41248 32366 41276 33594
rect 43272 33590 43300 33798
rect 43260 33584 43312 33590
rect 43260 33526 43312 33532
rect 42800 33448 42852 33454
rect 42800 33390 42852 33396
rect 42812 33130 42840 33390
rect 42628 33102 42840 33130
rect 43456 33114 43484 33934
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 44364 33312 44416 33318
rect 44364 33254 44416 33260
rect 43444 33108 43496 33114
rect 42064 32836 42116 32842
rect 42064 32778 42116 32784
rect 42076 32570 42104 32778
rect 42524 32768 42576 32774
rect 42524 32710 42576 32716
rect 42536 32570 42564 32710
rect 42064 32564 42116 32570
rect 42064 32506 42116 32512
rect 42524 32564 42576 32570
rect 42524 32506 42576 32512
rect 41236 32360 41288 32366
rect 41236 32302 41288 32308
rect 38384 32224 38436 32230
rect 38384 32166 38436 32172
rect 41788 32224 41840 32230
rect 41788 32166 41840 32172
rect 36912 31408 36964 31414
rect 36912 31350 36964 31356
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 38396 30190 38424 32166
rect 41800 31754 41828 32166
rect 41788 31748 41840 31754
rect 41788 31690 41840 31696
rect 42628 31686 42656 33102
rect 43444 33050 43496 33056
rect 43352 33040 43404 33046
rect 43352 32982 43404 32988
rect 42708 32564 42760 32570
rect 42708 32506 42760 32512
rect 42720 32366 42748 32506
rect 42800 32428 42852 32434
rect 42800 32370 42852 32376
rect 42708 32360 42760 32366
rect 42708 32302 42760 32308
rect 42812 32026 42840 32370
rect 42800 32020 42852 32026
rect 42800 31962 42852 31968
rect 42892 31884 42944 31890
rect 42892 31826 42944 31832
rect 42616 31680 42668 31686
rect 42616 31622 42668 31628
rect 41880 31340 41932 31346
rect 41880 31282 41932 31288
rect 41892 30394 41920 31282
rect 42628 31210 42656 31622
rect 42616 31204 42668 31210
rect 42616 31146 42668 31152
rect 42628 30734 42656 31146
rect 42708 31136 42760 31142
rect 42708 31078 42760 31084
rect 42720 30734 42748 31078
rect 42616 30728 42668 30734
rect 42616 30670 42668 30676
rect 42708 30728 42760 30734
rect 42708 30670 42760 30676
rect 41880 30388 41932 30394
rect 41880 30330 41932 30336
rect 38384 30184 38436 30190
rect 38384 30126 38436 30132
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 35072 28552 35124 28558
rect 35072 28494 35124 28500
rect 35084 28082 35112 28494
rect 35072 28076 35124 28082
rect 35072 28018 35124 28024
rect 31944 27872 31996 27878
rect 31944 27814 31996 27820
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 31956 27402 31984 27814
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 31944 27396 31996 27402
rect 31944 27338 31996 27344
rect 32324 27062 32352 27406
rect 32312 27056 32364 27062
rect 32312 26998 32364 27004
rect 32324 26926 32352 26998
rect 32968 26994 32996 27814
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35452 27470 35480 28970
rect 36176 28960 36228 28966
rect 36176 28902 36228 28908
rect 36188 28490 36216 28902
rect 36176 28484 36228 28490
rect 36176 28426 36228 28432
rect 37648 28416 37700 28422
rect 37648 28358 37700 28364
rect 37660 28082 37688 28358
rect 38396 28082 38424 30126
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 37648 28076 37700 28082
rect 37648 28018 37700 28024
rect 37740 28076 37792 28082
rect 37740 28018 37792 28024
rect 38384 28076 38436 28082
rect 38384 28018 38436 28024
rect 37464 27872 37516 27878
rect 37464 27814 37516 27820
rect 37476 27606 37504 27814
rect 37464 27600 37516 27606
rect 37464 27542 37516 27548
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 37004 27464 37056 27470
rect 37004 27406 37056 27412
rect 33416 27328 33468 27334
rect 33416 27270 33468 27276
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 32312 26920 32364 26926
rect 32312 26862 32364 26868
rect 32324 26382 32352 26862
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 30012 26240 30064 26246
rect 30012 26182 30064 26188
rect 29920 25968 29972 25974
rect 29920 25910 29972 25916
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 25044 25696 25096 25702
rect 25044 25638 25096 25644
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29644 24608 29696 24614
rect 29644 24550 29696 24556
rect 29656 24206 29684 24550
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 23322 25636 23666
rect 25792 23662 25820 24006
rect 25872 23724 25924 23730
rect 25872 23666 25924 23672
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25884 23322 25912 23666
rect 25596 23316 25648 23322
rect 25596 23258 25648 23264
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20364 21622 20392 21966
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18064 20058 18092 21490
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 21146 18736 21286
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18800 20330 18828 21422
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 19378 18460 19654
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 16908 18708 16988 18714
rect 16856 18702 16988 18708
rect 16304 18692 16356 18698
rect 16868 18686 16988 18702
rect 16304 18634 16356 18640
rect 16316 18290 16344 18634
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16960 18222 16988 18686
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16960 17746 16988 18158
rect 17052 17882 17080 18226
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16960 17202 16988 17682
rect 17420 17270 17448 19110
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18616 17610 18644 18702
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18800 18358 18828 18566
rect 18984 18426 19012 20334
rect 19076 20262 19104 21286
rect 20088 20942 20116 21422
rect 21008 20942 21036 21966
rect 28920 21486 28948 23054
rect 29196 23050 29224 24142
rect 29840 23730 29868 24754
rect 29932 24614 29960 25910
rect 30024 25906 30052 26182
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 31772 25702 31800 26318
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32600 25906 32628 26250
rect 33336 25906 33364 26726
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 33428 25702 33456 27270
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 33612 25838 33640 26726
rect 34532 26382 34560 27406
rect 37016 26994 37044 27406
rect 37752 27130 37780 28018
rect 37924 27872 37976 27878
rect 37924 27814 37976 27820
rect 37740 27124 37792 27130
rect 37740 27066 37792 27072
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 37832 26444 37884 26450
rect 37832 26386 37884 26392
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 33692 26240 33744 26246
rect 33692 26182 33744 26188
rect 33704 25974 33732 26182
rect 33692 25968 33744 25974
rect 33692 25910 33744 25916
rect 33600 25832 33652 25838
rect 33600 25774 33652 25780
rect 31576 25696 31628 25702
rect 31576 25638 31628 25644
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 33232 25696 33284 25702
rect 33232 25638 33284 25644
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 31588 25294 31616 25638
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29932 24274 29960 24550
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 29932 23730 29960 24210
rect 30668 23798 30696 25230
rect 31772 24886 31800 25638
rect 33244 25498 33272 25638
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 31760 24880 31812 24886
rect 31760 24822 31812 24828
rect 31668 24200 31720 24206
rect 31668 24142 31720 24148
rect 31680 23866 31708 24142
rect 31668 23860 31720 23866
rect 31668 23802 31720 23808
rect 30656 23792 30708 23798
rect 30656 23734 30708 23740
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21468 21146 21496 21286
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20466 20024 20878
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20088 20398 20116 20878
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18892 17338 18920 18158
rect 19076 17882 19104 18226
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16132 16794 16160 16934
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 16250 16252 16594
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16500 15706 16528 16526
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16868 15502 16896 15846
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14822 14872 14962
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 11808 13870 11836 14214
rect 14292 14006 14320 14214
rect 14476 14074 14504 14350
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14844 14006 14872 14758
rect 15120 14482 15148 15438
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11716 12594 11744 13670
rect 11808 13190 11836 13806
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13462 12572 13670
rect 12636 13530 12664 13942
rect 15120 13938 15148 14418
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11808 12782 11836 13126
rect 11900 12918 11928 13126
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11796 12640 11848 12646
rect 11716 12588 11796 12594
rect 11716 12582 11848 12588
rect 11716 12566 11836 12582
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 10810 9812 11698
rect 10520 11218 10548 12174
rect 11808 11626 11836 12566
rect 11900 12442 11928 12854
rect 12268 12850 12296 13194
rect 12820 12986 12848 13874
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12912 13258 12940 13398
rect 15764 13394 15792 14350
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 16040 13326 16068 13670
rect 17144 13530 17172 14554
rect 17788 14414 17816 16390
rect 19352 15586 19380 20198
rect 20088 19854 20116 20334
rect 22020 19854 22048 21286
rect 28920 20942 28948 21422
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20058 22140 20810
rect 22388 20602 22416 20878
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22572 20466 22600 20742
rect 27908 20466 27936 20878
rect 29932 20466 29960 20878
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 28276 20058 28304 20402
rect 30024 20058 30052 20402
rect 30484 20058 30512 20742
rect 30760 20602 30788 21490
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 30852 21146 30880 21422
rect 30840 21140 30892 21146
rect 30840 21082 30892 21088
rect 31036 20602 31064 21490
rect 31772 21350 31800 24822
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31864 24274 31892 24550
rect 33152 24410 33180 25298
rect 33968 25288 34020 25294
rect 33968 25230 34020 25236
rect 33876 25152 33928 25158
rect 33876 25094 33928 25100
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 31852 24268 31904 24274
rect 31852 24210 31904 24216
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 31852 24132 31904 24138
rect 31852 24074 31904 24080
rect 31864 23322 31892 24074
rect 32968 23730 32996 24142
rect 32956 23724 33008 23730
rect 32956 23666 33008 23672
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33520 23322 33548 23666
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 32864 22160 32916 22166
rect 32864 22102 32916 22108
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 32588 21344 32640 21350
rect 32588 21286 32640 21292
rect 31772 20874 31800 21286
rect 32600 20942 32628 21286
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 31024 20596 31076 20602
rect 31024 20538 31076 20544
rect 32324 20398 32352 20878
rect 32876 20534 32904 22102
rect 33888 22030 33916 25094
rect 33980 24206 34008 25230
rect 34532 24614 34560 26318
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 34704 25220 34756 25226
rect 34704 25162 34756 25168
rect 34520 24608 34572 24614
rect 34520 24550 34572 24556
rect 34716 24342 34744 25162
rect 36084 24880 36136 24886
rect 36084 24822 36136 24828
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 35900 24608 35952 24614
rect 35900 24550 35952 24556
rect 34704 24336 34756 24342
rect 34704 24278 34756 24284
rect 34808 24274 34836 24550
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24268 34848 24274
rect 34796 24210 34848 24216
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34624 23866 34652 24142
rect 34612 23860 34664 23866
rect 34612 23802 34664 23808
rect 35912 23798 35940 24550
rect 36096 24138 36124 24822
rect 36280 24818 36308 25230
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 36084 24132 36136 24138
rect 36084 24074 36136 24080
rect 35900 23792 35952 23798
rect 35900 23734 35952 23740
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35912 22098 35940 23734
rect 36372 23730 36400 25230
rect 36912 24812 36964 24818
rect 36912 24754 36964 24760
rect 36924 23866 36952 24754
rect 37844 24682 37872 26386
rect 37936 26382 37964 27814
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 38120 27062 38148 27406
rect 38672 27062 38700 28970
rect 38752 28552 38804 28558
rect 38752 28494 38804 28500
rect 38764 28150 38792 28494
rect 38752 28144 38804 28150
rect 38752 28086 38804 28092
rect 42628 28082 42656 30670
rect 42904 30326 42932 31826
rect 42892 30320 42944 30326
rect 42892 30262 42944 30268
rect 43076 30252 43128 30258
rect 43076 30194 43128 30200
rect 43088 29170 43116 30194
rect 43364 30054 43392 32982
rect 44376 32842 44404 33254
rect 43628 32836 43680 32842
rect 43628 32778 43680 32784
rect 44364 32836 44416 32842
rect 44364 32778 44416 32784
rect 44548 32836 44600 32842
rect 44548 32778 44600 32784
rect 43640 32434 43668 32778
rect 43720 32564 43772 32570
rect 43720 32506 43772 32512
rect 43628 32428 43680 32434
rect 43628 32370 43680 32376
rect 43640 32298 43668 32370
rect 43628 32292 43680 32298
rect 43628 32234 43680 32240
rect 43536 32224 43588 32230
rect 43536 32166 43588 32172
rect 43548 31414 43576 32166
rect 43640 31822 43668 32234
rect 43732 31890 43760 32506
rect 44456 32496 44508 32502
rect 44456 32438 44508 32444
rect 44088 32292 44140 32298
rect 44088 32234 44140 32240
rect 44100 31890 44128 32234
rect 43720 31884 43772 31890
rect 43720 31826 43772 31832
rect 44088 31884 44140 31890
rect 44088 31826 44140 31832
rect 43628 31816 43680 31822
rect 43628 31758 43680 31764
rect 43536 31408 43588 31414
rect 43536 31350 43588 31356
rect 43628 31136 43680 31142
rect 43628 31078 43680 31084
rect 43640 30258 43668 31078
rect 44100 30938 44128 31826
rect 44468 31414 44496 32438
rect 44560 32026 44588 32778
rect 45376 32768 45428 32774
rect 45376 32710 45428 32716
rect 46020 32768 46072 32774
rect 46020 32710 46072 32716
rect 45388 32026 45416 32710
rect 44548 32020 44600 32026
rect 44548 31962 44600 31968
rect 45376 32020 45428 32026
rect 45376 31962 45428 31968
rect 46032 31822 46060 32710
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 46204 32428 46256 32434
rect 46204 32370 46256 32376
rect 46216 32026 46244 32370
rect 46480 32360 46532 32366
rect 46480 32302 46532 32308
rect 46204 32020 46256 32026
rect 46204 31962 46256 31968
rect 46020 31816 46072 31822
rect 46020 31758 46072 31764
rect 44456 31408 44508 31414
rect 44456 31350 44508 31356
rect 44468 30938 44496 31350
rect 46492 31210 46520 32302
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 46480 31204 46532 31210
rect 46480 31146 46532 31152
rect 44088 30932 44140 30938
rect 44088 30874 44140 30880
rect 44456 30932 44508 30938
rect 44456 30874 44508 30880
rect 43628 30252 43680 30258
rect 43628 30194 43680 30200
rect 43352 30048 43404 30054
rect 43352 29990 43404 29996
rect 43076 29164 43128 29170
rect 43076 29106 43128 29112
rect 42892 28960 42944 28966
rect 42892 28902 42944 28908
rect 42800 28416 42852 28422
rect 42800 28358 42852 28364
rect 41880 28076 41932 28082
rect 41880 28018 41932 28024
rect 42616 28076 42668 28082
rect 42616 28018 42668 28024
rect 40040 27872 40092 27878
rect 40040 27814 40092 27820
rect 40132 27872 40184 27878
rect 40132 27814 40184 27820
rect 39488 27328 39540 27334
rect 39488 27270 39540 27276
rect 39500 27062 39528 27270
rect 38108 27056 38160 27062
rect 38108 26998 38160 27004
rect 38660 27056 38712 27062
rect 38660 26998 38712 27004
rect 39488 27056 39540 27062
rect 39488 26998 39540 27004
rect 37924 26376 37976 26382
rect 37924 26318 37976 26324
rect 38120 24818 38148 26998
rect 40052 26790 40080 27814
rect 40144 27402 40172 27814
rect 41892 27674 41920 28018
rect 41880 27668 41932 27674
rect 41880 27610 41932 27616
rect 42064 27464 42116 27470
rect 42064 27406 42116 27412
rect 40132 27396 40184 27402
rect 40132 27338 40184 27344
rect 40316 27396 40368 27402
rect 40316 27338 40368 27344
rect 40328 27062 40356 27338
rect 40500 27328 40552 27334
rect 40500 27270 40552 27276
rect 40316 27056 40368 27062
rect 40316 26998 40368 27004
rect 40512 26994 40540 27270
rect 40500 26988 40552 26994
rect 40500 26930 40552 26936
rect 40040 26784 40092 26790
rect 40040 26726 40092 26732
rect 40684 26784 40736 26790
rect 40684 26726 40736 26732
rect 40696 26586 40724 26726
rect 40684 26580 40736 26586
rect 40684 26522 40736 26528
rect 42076 26382 42104 27406
rect 42812 27402 42840 28358
rect 42904 27674 42932 28902
rect 42984 28552 43036 28558
rect 42984 28494 43036 28500
rect 42996 28218 43024 28494
rect 43088 28490 43116 29106
rect 43260 29096 43312 29102
rect 43260 29038 43312 29044
rect 43272 28558 43300 29038
rect 43364 28966 43392 29990
rect 46492 29646 46520 31146
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 43904 29640 43956 29646
rect 43904 29582 43956 29588
rect 46480 29640 46532 29646
rect 46480 29582 46532 29588
rect 43916 29306 43944 29582
rect 44640 29504 44692 29510
rect 44640 29446 44692 29452
rect 43904 29300 43956 29306
rect 43904 29242 43956 29248
rect 44652 29186 44680 29446
rect 44560 29170 44680 29186
rect 45284 29232 45336 29238
rect 45284 29174 45336 29180
rect 45376 29232 45428 29238
rect 45376 29174 45428 29180
rect 44548 29164 44680 29170
rect 44600 29158 44680 29164
rect 44548 29106 44600 29112
rect 43352 28960 43404 28966
rect 43352 28902 43404 28908
rect 44652 28626 44680 29158
rect 44732 29164 44784 29170
rect 44732 29106 44784 29112
rect 44640 28620 44692 28626
rect 44640 28562 44692 28568
rect 44744 28558 44772 29106
rect 43260 28552 43312 28558
rect 43260 28494 43312 28500
rect 43720 28552 43772 28558
rect 43720 28494 43772 28500
rect 44732 28552 44784 28558
rect 44732 28494 44784 28500
rect 43076 28484 43128 28490
rect 43076 28426 43128 28432
rect 42984 28212 43036 28218
rect 42984 28154 43036 28160
rect 42892 27668 42944 27674
rect 42892 27610 42944 27616
rect 42800 27396 42852 27402
rect 42800 27338 42852 27344
rect 42064 26376 42116 26382
rect 42064 26318 42116 26324
rect 42708 26376 42760 26382
rect 42708 26318 42760 26324
rect 41880 26308 41932 26314
rect 41880 26250 41932 26256
rect 41892 26042 41920 26250
rect 41880 26036 41932 26042
rect 41880 25978 41932 25984
rect 42720 25974 42748 26318
rect 42708 25968 42760 25974
rect 42708 25910 42760 25916
rect 42064 25900 42116 25906
rect 42064 25842 42116 25848
rect 40316 25696 40368 25702
rect 40316 25638 40368 25644
rect 40328 25294 40356 25638
rect 38568 25288 38620 25294
rect 38568 25230 38620 25236
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40316 25288 40368 25294
rect 40316 25230 40368 25236
rect 38580 24886 38608 25230
rect 40052 24886 40080 25230
rect 40224 25220 40276 25226
rect 40224 25162 40276 25168
rect 38568 24880 38620 24886
rect 38568 24822 38620 24828
rect 40040 24880 40092 24886
rect 40040 24822 40092 24828
rect 38108 24812 38160 24818
rect 38108 24754 38160 24760
rect 37832 24676 37884 24682
rect 37832 24618 37884 24624
rect 38120 24274 38148 24754
rect 38200 24744 38252 24750
rect 38200 24686 38252 24692
rect 38108 24268 38160 24274
rect 38108 24210 38160 24216
rect 38120 23866 38148 24210
rect 38212 23866 38240 24686
rect 36912 23860 36964 23866
rect 36912 23802 36964 23808
rect 38108 23860 38160 23866
rect 38108 23802 38160 23808
rect 38200 23860 38252 23866
rect 38200 23802 38252 23808
rect 40052 23730 40080 24822
rect 40236 24818 40264 25162
rect 41696 25152 41748 25158
rect 41696 25094 41748 25100
rect 41420 24880 41472 24886
rect 41420 24822 41472 24828
rect 40224 24812 40276 24818
rect 40224 24754 40276 24760
rect 40868 24608 40920 24614
rect 40868 24550 40920 24556
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 37924 23724 37976 23730
rect 37924 23666 37976 23672
rect 40040 23724 40092 23730
rect 40040 23666 40092 23672
rect 40316 23724 40368 23730
rect 40316 23666 40368 23672
rect 37936 23322 37964 23666
rect 40328 23322 40356 23666
rect 37924 23316 37976 23322
rect 37924 23258 37976 23264
rect 40316 23316 40368 23322
rect 40316 23258 40368 23264
rect 40880 23118 40908 24550
rect 41432 24410 41460 24822
rect 41604 24608 41656 24614
rect 41604 24550 41656 24556
rect 41420 24404 41472 24410
rect 41420 24346 41472 24352
rect 41144 24064 41196 24070
rect 41144 24006 41196 24012
rect 40868 23112 40920 23118
rect 40868 23054 40920 23060
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 38200 22636 38252 22642
rect 38200 22578 38252 22584
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 33232 21412 33284 21418
rect 33232 21354 33284 21360
rect 32864 20528 32916 20534
rect 32864 20470 32916 20476
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30472 20052 30524 20058
rect 30472 19994 30524 20000
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 19174 20116 19790
rect 32140 19446 32168 19790
rect 32128 19440 32180 19446
rect 32128 19382 32180 19388
rect 32324 19378 32352 20334
rect 33244 19854 33272 21354
rect 33508 20800 33560 20806
rect 33508 20742 33560 20748
rect 33520 20058 33548 20742
rect 34072 20058 34100 21966
rect 35912 21622 35940 22034
rect 36636 21956 36688 21962
rect 36636 21898 36688 21904
rect 35900 21616 35952 21622
rect 35900 21558 35952 21564
rect 34152 21548 34204 21554
rect 34152 21490 34204 21496
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 34164 21146 34192 21490
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34532 19922 34560 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20810
rect 35452 20602 35480 21490
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 35544 20534 35572 21490
rect 35912 20942 35940 21558
rect 36268 21480 36320 21486
rect 36268 21422 36320 21428
rect 36280 21146 36308 21422
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 35532 20528 35584 20534
rect 35532 20470 35584 20476
rect 35912 20466 35940 20878
rect 36648 20602 36676 21898
rect 37568 21894 37596 22578
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37556 21888 37608 21894
rect 37556 21830 37608 21836
rect 37384 21418 37412 21830
rect 37568 21622 37596 21830
rect 37556 21616 37608 21622
rect 37556 21558 37608 21564
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 37372 21412 37424 21418
rect 37372 21354 37424 21360
rect 36820 21344 36872 21350
rect 36820 21286 36872 21292
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 36740 20534 36768 20878
rect 36728 20528 36780 20534
rect 36728 20470 36780 20476
rect 36832 20466 36860 21286
rect 37384 21078 37412 21354
rect 37372 21072 37424 21078
rect 37372 21014 37424 21020
rect 37752 20602 37780 21490
rect 37936 21010 37964 22374
rect 38212 21962 38240 22578
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 38200 21956 38252 21962
rect 38200 21898 38252 21904
rect 38212 21690 38240 21898
rect 38384 21888 38436 21894
rect 38384 21830 38436 21836
rect 38200 21684 38252 21690
rect 38200 21626 38252 21632
rect 38396 21146 38424 21830
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38856 21078 38884 21966
rect 39040 21146 39068 21966
rect 39212 21888 39264 21894
rect 39212 21830 39264 21836
rect 39120 21344 39172 21350
rect 39120 21286 39172 21292
rect 39028 21140 39080 21146
rect 39028 21082 39080 21088
rect 38844 21072 38896 21078
rect 38844 21014 38896 21020
rect 37924 21004 37976 21010
rect 37924 20946 37976 20952
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37936 20466 37964 20742
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 36820 20460 36872 20466
rect 36820 20402 36872 20408
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 38856 20330 38884 21014
rect 39132 21010 39160 21286
rect 39120 21004 39172 21010
rect 39120 20946 39172 20952
rect 39132 20534 39160 20946
rect 39224 20942 39252 21830
rect 39396 21548 39448 21554
rect 39396 21490 39448 21496
rect 39408 21146 39436 21490
rect 40776 21344 40828 21350
rect 40776 21286 40828 21292
rect 39396 21140 39448 21146
rect 39396 21082 39448 21088
rect 40788 20942 40816 21286
rect 39212 20936 39264 20942
rect 39212 20878 39264 20884
rect 40776 20936 40828 20942
rect 40776 20878 40828 20884
rect 39120 20528 39172 20534
rect 39120 20470 39172 20476
rect 38844 20324 38896 20330
rect 38844 20266 38896 20272
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 34520 19916 34572 19922
rect 34520 19858 34572 19864
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33704 19514 33732 19790
rect 33692 19508 33744 19514
rect 33692 19450 33744 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18222 20116 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20088 17610 20116 18158
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20732 16794 20760 18226
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 16726 20852 18702
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 17542 21036 18566
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21100 17338 21128 18702
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 21468 18086 21496 18226
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21100 16998 21128 17070
rect 21468 16998 21496 18022
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20824 16590 20852 16662
rect 21100 16658 21128 16934
rect 21652 16794 21680 17546
rect 22112 17542 22140 18226
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17270 22140 17478
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 22204 16590 22232 18022
rect 22940 17814 22968 18226
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 22928 17808 22980 17814
rect 22928 17750 22980 17756
rect 22940 17338 22968 17750
rect 36924 17610 36952 18022
rect 36912 17604 36964 17610
rect 36912 17546 36964 17552
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 37384 17270 37412 18702
rect 37476 18222 37504 18702
rect 37844 18698 37872 19110
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37476 17678 37504 18158
rect 38844 18080 38896 18086
rect 38844 18022 38896 18028
rect 38752 17876 38804 17882
rect 38752 17818 38804 17824
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 17264 37424 17270
rect 37372 17206 37424 17212
rect 37476 17202 37504 17614
rect 38764 17338 38792 17818
rect 38856 17746 38884 18022
rect 38844 17740 38896 17746
rect 38844 17682 38896 17688
rect 38948 17678 38976 18566
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 38752 17332 38804 17338
rect 38752 17274 38804 17280
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20824 16250 20852 16526
rect 22388 16522 22416 16934
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19168 15570 19380 15586
rect 19168 15564 19392 15570
rect 19168 15558 19340 15564
rect 19168 14414 19196 15558
rect 19340 15506 19392 15512
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19260 15042 19288 15438
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 15162 19380 15370
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19444 15094 19472 15846
rect 19996 15434 20024 15982
rect 20088 15910 20116 16050
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15144 20024 15370
rect 19812 15116 20024 15144
rect 19432 15088 19484 15094
rect 19260 15014 19380 15042
rect 19432 15030 19484 15036
rect 19352 14482 19380 15014
rect 19812 14550 19840 15116
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14006 20024 14282
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12850 12940 13194
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12268 12714 12296 12786
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12268 11830 12296 12650
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 10810 11744 11018
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 11900 10674 11928 11494
rect 12268 11354 12296 11766
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 6840 10266 6868 10406
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 19996 10130 20024 13942
rect 20088 13530 20116 15846
rect 20272 14822 20300 16118
rect 20824 15706 20852 16186
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20916 15434 20944 16050
rect 22388 15722 22416 16458
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 22296 15694 22416 15722
rect 22296 15570 22324 15694
rect 40052 15570 40080 17138
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 40040 15564 40092 15570
rect 40040 15506 40092 15512
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 20904 15428 20956 15434
rect 20904 15370 20956 15376
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20272 14074 20300 14758
rect 20456 14618 20484 15030
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20456 13938 20484 14554
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20364 11150 20392 13806
rect 20456 13326 20484 13874
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20548 13258 20576 15302
rect 20916 15026 20944 15370
rect 22112 15162 22140 15370
rect 22204 15162 22232 15438
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14618 20668 14894
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 21928 14618 21956 14758
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 20640 14006 20668 14554
rect 22204 14414 22232 15098
rect 22296 14414 22324 15506
rect 39580 15496 39632 15502
rect 39580 15438 39632 15444
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 15094 22692 15302
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 39592 15026 39620 15438
rect 39580 15020 39632 15026
rect 39580 14962 39632 14968
rect 39120 14952 39172 14958
rect 39120 14894 39172 14900
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 21468 13530 21496 14350
rect 39132 13870 39160 14894
rect 39948 14408 40000 14414
rect 39948 14350 40000 14356
rect 39960 13870 39988 14350
rect 39120 13864 39172 13870
rect 39120 13806 39172 13812
rect 39948 13864 40000 13870
rect 39948 13806 40000 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 39132 12782 39160 13806
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40052 12918 40080 13262
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39120 12776 39172 12782
rect 39120 12718 39172 12724
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 38844 12232 38896 12238
rect 38844 12174 38896 12180
rect 38384 11552 38436 11558
rect 38384 11494 38436 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 38396 11082 38424 11494
rect 38856 11082 38884 12174
rect 39132 11762 39160 12718
rect 39304 12232 39356 12238
rect 39304 12174 39356 12180
rect 39316 11830 39344 12174
rect 39304 11824 39356 11830
rect 39304 11766 39356 11772
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 39580 11756 39632 11762
rect 39580 11698 39632 11704
rect 39132 11150 39160 11698
rect 39592 11354 39620 11698
rect 39580 11348 39632 11354
rect 39580 11290 39632 11296
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 38844 11076 38896 11082
rect 38844 11018 38896 11024
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 20272 10062 20300 10950
rect 40144 10674 40172 20198
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40972 18766 41000 19110
rect 40776 18760 40828 18766
rect 40776 18702 40828 18708
rect 40960 18760 41012 18766
rect 40960 18702 41012 18708
rect 40788 18290 40816 18702
rect 40776 18284 40828 18290
rect 40776 18226 40828 18232
rect 40960 18284 41012 18290
rect 40960 18226 41012 18232
rect 40316 18080 40368 18086
rect 40316 18022 40368 18028
rect 40328 17202 40356 18022
rect 40788 17202 40816 18226
rect 40316 17196 40368 17202
rect 40316 17138 40368 17144
rect 40776 17196 40828 17202
rect 40776 17138 40828 17144
rect 40972 16794 41000 18226
rect 41156 17610 41184 24006
rect 41432 22030 41460 24346
rect 41512 23520 41564 23526
rect 41512 23462 41564 23468
rect 41524 23322 41552 23462
rect 41512 23316 41564 23322
rect 41512 23258 41564 23264
rect 41616 23186 41644 24550
rect 41604 23180 41656 23186
rect 41604 23122 41656 23128
rect 41708 23118 41736 25094
rect 42076 24954 42104 25842
rect 42720 25294 42748 25910
rect 42904 25770 42932 27610
rect 42996 26926 43024 28154
rect 43088 28150 43116 28426
rect 43076 28144 43128 28150
rect 43076 28086 43128 28092
rect 43088 27656 43116 28086
rect 43168 27668 43220 27674
rect 43088 27628 43168 27656
rect 43088 26994 43116 27628
rect 43168 27610 43220 27616
rect 43732 27402 43760 28494
rect 45192 28416 45244 28422
rect 45192 28358 45244 28364
rect 43904 28212 43956 28218
rect 43904 28154 43956 28160
rect 43916 27402 43944 28154
rect 44916 28144 44968 28150
rect 44916 28086 44968 28092
rect 44928 27470 44956 28086
rect 45204 28082 45232 28358
rect 45192 28076 45244 28082
rect 45192 28018 45244 28024
rect 45296 27606 45324 29174
rect 45388 28218 45416 29174
rect 46296 28960 46348 28966
rect 46296 28902 46348 28908
rect 46308 28558 46336 28902
rect 46492 28558 46520 29582
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 46296 28552 46348 28558
rect 46296 28494 46348 28500
rect 46480 28552 46532 28558
rect 46480 28494 46532 28500
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 45376 28212 45428 28218
rect 45376 28154 45428 28160
rect 45376 28076 45428 28082
rect 45376 28018 45428 28024
rect 45284 27600 45336 27606
rect 45284 27542 45336 27548
rect 45388 27470 45416 28018
rect 44916 27464 44968 27470
rect 44916 27406 44968 27412
rect 45376 27464 45428 27470
rect 45376 27406 45428 27412
rect 43720 27396 43772 27402
rect 43720 27338 43772 27344
rect 43904 27396 43956 27402
rect 43904 27338 43956 27344
rect 43732 27062 43760 27338
rect 43916 27130 43944 27338
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 43904 27124 43956 27130
rect 43904 27066 43956 27072
rect 43720 27056 43772 27062
rect 43720 26998 43772 27004
rect 43076 26988 43128 26994
rect 43076 26930 43128 26936
rect 43732 26926 43760 26998
rect 58072 26988 58124 26994
rect 58072 26930 58124 26936
rect 42984 26920 43036 26926
rect 42984 26862 43036 26868
rect 43720 26920 43772 26926
rect 43720 26862 43772 26868
rect 43444 26852 43496 26858
rect 43444 26794 43496 26800
rect 43352 26784 43404 26790
rect 43352 26726 43404 26732
rect 43168 26580 43220 26586
rect 43168 26522 43220 26528
rect 43180 26382 43208 26522
rect 43168 26376 43220 26382
rect 43168 26318 43220 26324
rect 43180 25838 43208 26318
rect 43168 25832 43220 25838
rect 43168 25774 43220 25780
rect 42892 25764 42944 25770
rect 42892 25706 42944 25712
rect 42708 25288 42760 25294
rect 42708 25230 42760 25236
rect 42064 24948 42116 24954
rect 42064 24890 42116 24896
rect 42720 24410 42748 25230
rect 42904 24954 42932 25706
rect 42892 24948 42944 24954
rect 42892 24890 42944 24896
rect 42984 24880 43036 24886
rect 42984 24822 43036 24828
rect 42708 24404 42760 24410
rect 42708 24346 42760 24352
rect 42996 23866 43024 24822
rect 43180 24614 43208 25774
rect 43364 24818 43392 26726
rect 43456 26586 43484 26794
rect 44364 26784 44416 26790
rect 44364 26726 44416 26732
rect 43444 26580 43496 26586
rect 43444 26522 43496 26528
rect 43996 26376 44048 26382
rect 43996 26318 44048 26324
rect 44008 25906 44036 26318
rect 44180 26308 44232 26314
rect 44180 26250 44232 26256
rect 44192 25906 44220 26250
rect 44376 25906 44404 26726
rect 45560 26580 45612 26586
rect 45560 26522 45612 26528
rect 45572 25974 45600 26522
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 45560 25968 45612 25974
rect 45560 25910 45612 25916
rect 43444 25900 43496 25906
rect 43444 25842 43496 25848
rect 43996 25900 44048 25906
rect 43996 25842 44048 25848
rect 44180 25900 44232 25906
rect 44180 25842 44232 25848
rect 44364 25900 44416 25906
rect 44364 25842 44416 25848
rect 43456 24886 43484 25842
rect 44192 25498 44220 25842
rect 44180 25492 44232 25498
rect 44180 25434 44232 25440
rect 43812 25220 43864 25226
rect 43812 25162 43864 25168
rect 43824 24954 43852 25162
rect 43812 24948 43864 24954
rect 43812 24890 43864 24896
rect 43444 24880 43496 24886
rect 43444 24822 43496 24828
rect 44192 24818 44220 25434
rect 43352 24812 43404 24818
rect 43352 24754 43404 24760
rect 44180 24812 44232 24818
rect 44180 24754 44232 24760
rect 44376 24682 44404 25842
rect 58084 25702 58112 26930
rect 58256 26784 58308 26790
rect 58256 26726 58308 26732
rect 58268 26625 58296 26726
rect 58254 26616 58310 26625
rect 58254 26551 58310 26560
rect 58072 25696 58124 25702
rect 58072 25638 58124 25644
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 44364 24676 44416 24682
rect 44364 24618 44416 24624
rect 43168 24608 43220 24614
rect 43168 24550 43220 24556
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 42984 23860 43036 23866
rect 42984 23802 43036 23808
rect 42616 23724 42668 23730
rect 42616 23666 42668 23672
rect 43628 23724 43680 23730
rect 43628 23666 43680 23672
rect 42628 23254 42656 23666
rect 42616 23248 42668 23254
rect 42616 23190 42668 23196
rect 41696 23112 41748 23118
rect 41696 23054 41748 23060
rect 41604 22432 41656 22438
rect 41604 22374 41656 22380
rect 42616 22432 42668 22438
rect 42616 22374 42668 22380
rect 41616 22030 41644 22374
rect 41420 22024 41472 22030
rect 41420 21966 41472 21972
rect 41604 22024 41656 22030
rect 41604 21966 41656 21972
rect 41432 21554 41460 21966
rect 41880 21956 41932 21962
rect 41880 21898 41932 21904
rect 41420 21548 41472 21554
rect 41420 21490 41472 21496
rect 41432 21146 41460 21490
rect 41892 21146 41920 21898
rect 42340 21548 42392 21554
rect 42340 21490 42392 21496
rect 41420 21140 41472 21146
rect 41420 21082 41472 21088
rect 41880 21140 41932 21146
rect 41880 21082 41932 21088
rect 42352 21010 42380 21490
rect 42340 21004 42392 21010
rect 42340 20946 42392 20952
rect 42628 20942 42656 22374
rect 42892 22160 42944 22166
rect 42892 22102 42944 22108
rect 42904 21554 42932 22102
rect 43352 22024 43404 22030
rect 43352 21966 43404 21972
rect 43364 21690 43392 21966
rect 43640 21894 43668 23666
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 43720 22024 43772 22030
rect 43720 21966 43772 21972
rect 43628 21888 43680 21894
rect 43628 21830 43680 21836
rect 43352 21684 43404 21690
rect 43352 21626 43404 21632
rect 42892 21548 42944 21554
rect 42892 21490 42944 21496
rect 43732 21146 43760 21966
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 43720 21140 43772 21146
rect 43720 21082 43772 21088
rect 42616 20936 42668 20942
rect 42616 20878 42668 20884
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 42800 19168 42852 19174
rect 42800 19110 42852 19116
rect 42616 18624 42668 18630
rect 42616 18566 42668 18572
rect 41972 18284 42024 18290
rect 41972 18226 42024 18232
rect 41144 17604 41196 17610
rect 41144 17546 41196 17552
rect 40960 16788 41012 16794
rect 40960 16730 41012 16736
rect 41156 16590 41184 17546
rect 41984 17338 42012 18226
rect 42628 18086 42656 18566
rect 42616 18080 42668 18086
rect 42616 18022 42668 18028
rect 42812 17338 42840 19110
rect 44456 18760 44508 18766
rect 44456 18702 44508 18708
rect 44468 18358 44496 18702
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 44456 18352 44508 18358
rect 44456 18294 44508 18300
rect 43996 18284 44048 18290
rect 43996 18226 44048 18232
rect 43352 18080 43404 18086
rect 43352 18022 43404 18028
rect 43364 17882 43392 18022
rect 43352 17876 43404 17882
rect 43352 17818 43404 17824
rect 43444 17740 43496 17746
rect 43444 17682 43496 17688
rect 42892 17604 42944 17610
rect 42892 17546 42944 17552
rect 41972 17332 42024 17338
rect 41972 17274 42024 17280
rect 42800 17332 42852 17338
rect 42800 17274 42852 17280
rect 42800 16992 42852 16998
rect 42800 16934 42852 16940
rect 42812 16658 42840 16934
rect 42800 16652 42852 16658
rect 42800 16594 42852 16600
rect 41144 16584 41196 16590
rect 41144 16526 41196 16532
rect 41156 16250 41184 16526
rect 41144 16244 41196 16250
rect 41144 16186 41196 16192
rect 42812 16114 42840 16594
rect 42800 16108 42852 16114
rect 42800 16050 42852 16056
rect 40316 15904 40368 15910
rect 40316 15846 40368 15852
rect 40592 15904 40644 15910
rect 40592 15846 40644 15852
rect 40328 14414 40356 15846
rect 40604 15502 40632 15846
rect 41972 15564 42024 15570
rect 41972 15506 42024 15512
rect 40592 15496 40644 15502
rect 40592 15438 40644 15444
rect 41880 15428 41932 15434
rect 41880 15370 41932 15376
rect 41892 15162 41920 15370
rect 41880 15156 41932 15162
rect 41880 15098 41932 15104
rect 41144 14816 41196 14822
rect 41144 14758 41196 14764
rect 40316 14408 40368 14414
rect 40316 14350 40368 14356
rect 41156 14006 41184 14758
rect 41984 14618 42012 15506
rect 42156 15496 42208 15502
rect 42156 15438 42208 15444
rect 41972 14612 42024 14618
rect 41972 14554 42024 14560
rect 42168 14074 42196 15438
rect 42156 14068 42208 14074
rect 42156 14010 42208 14016
rect 41144 14000 41196 14006
rect 41144 13942 41196 13948
rect 40868 12640 40920 12646
rect 40868 12582 40920 12588
rect 40880 11558 40908 12582
rect 42904 12238 42932 17546
rect 43456 15706 43484 17682
rect 43628 17672 43680 17678
rect 43628 17614 43680 17620
rect 43640 17338 43668 17614
rect 43904 17536 43956 17542
rect 43904 17478 43956 17484
rect 43628 17332 43680 17338
rect 43628 17274 43680 17280
rect 43812 16108 43864 16114
rect 43812 16050 43864 16056
rect 43444 15700 43496 15706
rect 43444 15642 43496 15648
rect 43720 15496 43772 15502
rect 43720 15438 43772 15444
rect 43352 14408 43404 14414
rect 43352 14350 43404 14356
rect 43364 13938 43392 14350
rect 43732 14346 43760 15438
rect 43824 15026 43852 16050
rect 43812 15020 43864 15026
rect 43812 14962 43864 14968
rect 43824 14414 43852 14962
rect 43812 14408 43864 14414
rect 43812 14350 43864 14356
rect 43720 14340 43772 14346
rect 43720 14282 43772 14288
rect 43916 14090 43944 17478
rect 44008 17066 44036 18226
rect 44548 18080 44600 18086
rect 44548 18022 44600 18028
rect 46296 18080 46348 18086
rect 46296 18022 46348 18028
rect 44560 17202 44588 18022
rect 44640 17672 44692 17678
rect 44640 17614 44692 17620
rect 45192 17672 45244 17678
rect 45192 17614 45244 17620
rect 44548 17196 44600 17202
rect 44548 17138 44600 17144
rect 43996 17060 44048 17066
rect 43996 17002 44048 17008
rect 44560 16658 44588 17138
rect 44548 16652 44600 16658
rect 44548 16594 44600 16600
rect 44652 16590 44680 17614
rect 45204 17270 45232 17614
rect 45192 17264 45244 17270
rect 45192 17206 45244 17212
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 44456 16584 44508 16590
rect 44456 16526 44508 16532
rect 44640 16584 44692 16590
rect 44640 16526 44692 16532
rect 44468 16182 44496 16526
rect 45572 16250 45600 17138
rect 46308 16998 46336 18022
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 46572 17196 46624 17202
rect 46572 17138 46624 17144
rect 46296 16992 46348 16998
rect 46296 16934 46348 16940
rect 46584 16794 46612 17138
rect 46572 16788 46624 16794
rect 46572 16730 46624 16736
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 45560 16244 45612 16250
rect 45560 16186 45612 16192
rect 44456 16176 44508 16182
rect 44456 16118 44508 16124
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 45836 15020 45888 15026
rect 45836 14962 45888 14968
rect 45560 14816 45612 14822
rect 45560 14758 45612 14764
rect 45192 14408 45244 14414
rect 45192 14350 45244 14356
rect 43824 14062 43944 14090
rect 44180 14068 44232 14074
rect 43352 13932 43404 13938
rect 43352 13874 43404 13880
rect 43364 13530 43392 13874
rect 43352 13524 43404 13530
rect 43352 13466 43404 13472
rect 43260 13252 43312 13258
rect 43260 13194 43312 13200
rect 43272 12986 43300 13194
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 43824 12918 43852 14062
rect 44180 14010 44232 14016
rect 44192 12918 44220 14010
rect 45204 14006 45232 14350
rect 45284 14272 45336 14278
rect 45284 14214 45336 14220
rect 45192 14000 45244 14006
rect 45192 13942 45244 13948
rect 44456 13932 44508 13938
rect 44456 13874 44508 13880
rect 44468 13530 44496 13874
rect 45296 13734 45324 14214
rect 45572 13938 45600 14758
rect 45848 14618 45876 14962
rect 45836 14612 45888 14618
rect 45836 14554 45888 14560
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 45560 13932 45612 13938
rect 45560 13874 45612 13880
rect 45284 13728 45336 13734
rect 45284 13670 45336 13676
rect 44456 13524 44508 13530
rect 44456 13466 44508 13472
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 45284 12980 45336 12986
rect 45284 12922 45336 12928
rect 43812 12912 43864 12918
rect 43812 12854 43864 12860
rect 44180 12912 44232 12918
rect 44180 12854 44232 12860
rect 43076 12640 43128 12646
rect 43076 12582 43128 12588
rect 44456 12640 44508 12646
rect 44456 12582 44508 12588
rect 42892 12232 42944 12238
rect 42892 12174 42944 12180
rect 41604 12096 41656 12102
rect 41604 12038 41656 12044
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 40868 11552 40920 11558
rect 40868 11494 40920 11500
rect 41432 11354 41460 11698
rect 41420 11348 41472 11354
rect 41420 11290 41472 11296
rect 41616 11150 41644 12038
rect 43088 11898 43116 12582
rect 43076 11892 43128 11898
rect 43076 11834 43128 11840
rect 42432 11552 42484 11558
rect 42432 11494 42484 11500
rect 41604 11144 41656 11150
rect 41604 11086 41656 11092
rect 42444 11082 42472 11494
rect 44468 11354 44496 12582
rect 44732 11552 44784 11558
rect 44732 11494 44784 11500
rect 44456 11348 44508 11354
rect 44456 11290 44508 11296
rect 44180 11144 44232 11150
rect 44180 11086 44232 11092
rect 42432 11076 42484 11082
rect 42432 11018 42484 11024
rect 42524 11076 42576 11082
rect 42524 11018 42576 11024
rect 43996 11076 44048 11082
rect 43996 11018 44048 11024
rect 42536 10674 42564 11018
rect 44008 10810 44036 11018
rect 43996 10804 44048 10810
rect 43996 10746 44048 10752
rect 40132 10668 40184 10674
rect 40132 10610 40184 10616
rect 42524 10668 42576 10674
rect 42524 10610 42576 10616
rect 40592 10464 40644 10470
rect 40592 10406 40644 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 22020 2446 22048 9862
rect 40604 9586 40632 10406
rect 42536 10130 42564 10610
rect 44192 10266 44220 11086
rect 44744 10742 44772 11494
rect 44732 10736 44784 10742
rect 44732 10678 44784 10684
rect 44456 10600 44508 10606
rect 44456 10542 44508 10548
rect 44180 10260 44232 10266
rect 44180 10202 44232 10208
rect 44468 10130 44496 10542
rect 42524 10124 42576 10130
rect 42524 10066 42576 10072
rect 44456 10124 44508 10130
rect 44456 10066 44508 10072
rect 42536 9654 42564 10066
rect 45296 10062 45324 12922
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 45836 11144 45888 11150
rect 45836 11086 45888 11092
rect 45848 10810 45876 11086
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 45836 10804 45888 10810
rect 45836 10746 45888 10752
rect 45284 10056 45336 10062
rect 45284 9998 45336 10004
rect 42800 9988 42852 9994
rect 42800 9930 42852 9936
rect 42524 9648 42576 9654
rect 42524 9590 42576 9596
rect 42812 9586 42840 9930
rect 57520 9920 57572 9926
rect 57520 9862 57572 9868
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 40592 9580 40644 9586
rect 40592 9522 40644 9528
rect 42800 9580 42852 9586
rect 42800 9522 42852 9528
rect 42616 9376 42668 9382
rect 42616 9318 42668 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 42628 2446 42656 9318
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 57532 3738 57560 9862
rect 57520 3732 57572 3738
rect 57520 3674 57572 3680
rect 57532 3534 57560 3674
rect 57520 3528 57572 3534
rect 57520 3470 57572 3476
rect 58254 3496 58310 3505
rect 58254 3431 58310 3440
rect 58268 3398 58296 3431
rect 58256 3392 58308 3398
rect 58256 3334 58308 3340
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 42616 2440 42668 2446
rect 42616 2382 42668 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 32 800 60 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2246
rect 42536 800 42564 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 18 200 74 800
rect 21270 200 21326 800
rect 42522 200 42578 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 3422 44920 3478 44976
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1766 22480 1822 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 58254 49036 58256 49056
rect 58256 49036 58308 49056
rect 58308 49036 58310 49056
rect 58254 49000 58310 49036
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 58254 26560 58310 26616
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 58254 3440 58310 3496
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 58249 49058 58315 49061
rect 59200 49058 59800 49088
rect 58249 49056 59800 49058
rect 58249 49000 58254 49056
rect 58310 49000 59800 49056
rect 58249 48998 59800 49000
rect 58249 48995 58315 48998
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 59200 48968 59800 48998
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 200 44978 800 45008
rect 3417 44978 3483 44981
rect 200 44976 3483 44978
rect 200 44920 3422 44976
rect 3478 44920 3483 44976
rect 200 44918 3483 44920
rect 200 44888 800 44918
rect 3417 44915 3483 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58249 26618 58315 26621
rect 59200 26618 59800 26648
rect 58249 26616 59800 26618
rect 58249 26560 58254 26616
rect 58310 26560 59800 26616
rect 58249 26558 59800 26560
rect 58249 26555 58315 26558
rect 59200 26528 59800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 58249 3498 58315 3501
rect 59200 3498 59800 3528
rect 58249 3496 59800 3498
rect 58249 3440 58254 3496
rect 58310 3440 59800 3496
rect 58249 3438 59800 3440
rect 58249 3435 58315 3438
rect 59200 3408 59800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23000 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1666464484
transform -1 0 16284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1666464484
transform -1 0 30820 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_clk_A
timestamp 1666464484
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_clk_A
timestamp 1666464484
transform 1 0 4416 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_clk_A
timestamp 1666464484
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_clk_A
timestamp 1666464484
transform 1 0 18768 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_clk_A
timestamp 1666464484
transform 1 0 9476 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_clk_A
timestamp 1666464484
transform 1 0 15824 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_clk_A
timestamp 1666464484
transform 1 0 24104 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_clk_A
timestamp 1666464484
transform 1 0 26404 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_clk_A
timestamp 1666464484
transform 1 0 32292 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_clk_A
timestamp 1666464484
transform 1 0 31004 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_clk_A
timestamp 1666464484
transform -1 0 38272 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_clk_A
timestamp 1666464484
transform 1 0 39192 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_clk_A
timestamp 1666464484
transform -1 0 44620 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_clk_A
timestamp 1666464484
transform 1 0 36800 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_clk_A
timestamp 1666464484
transform 1 0 32292 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_clk_A
timestamp 1666464484
transform 1 0 31648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_clk_A
timestamp 1666464484
transform 1 0 38272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_clk_A
timestamp 1666464484
transform 1 0 40940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_clk_A
timestamp 1666464484
transform -1 0 41400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_clk_A
timestamp 1666464484
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_clk_A
timestamp 1666464484
transform 1 0 23092 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_clk_A
timestamp 1666464484
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_clk_A
timestamp 1666464484
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_clk_A
timestamp 1666464484
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_clk_A
timestamp 1666464484
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_opt_1_0_clk_A
timestamp 1666464484
transform 1 0 10948 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_opt_2_0_clk_A
timestamp 1666464484
transform 1 0 42596 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_opt_3_0_clk_A
timestamp 1666464484
transform 1 0 40572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output1_A
timestamp 1666464484
transform 1 0 57500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_231
timestamp 1666464484
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1666464484
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1666464484
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1666464484
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1666464484
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1666464484
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1666464484
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1666464484
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1666464484
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1666464484
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1666464484
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_455
timestamp 1666464484
transform 1 0 42964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1666464484
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1666464484
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1666464484
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1666464484
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1666464484
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1666464484
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1666464484
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1666464484
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1666464484
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1666464484
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1666464484
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1666464484
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1666464484
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1666464484
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1666464484
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1666464484
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1666464484
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1666464484
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1666464484
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1666464484
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1666464484
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1666464484
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1666464484
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1666464484
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1666464484
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1666464484
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1666464484
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1666464484
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1666464484
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1666464484
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1666464484
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1666464484
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666464484
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1666464484
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1666464484
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1666464484
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1666464484
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1666464484
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1666464484
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1666464484
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1666464484
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1666464484
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1666464484
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1666464484
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1666464484
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1666464484
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1666464484
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1666464484
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1666464484
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_615
timestamp 1666464484
transform 1 0 57684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_623
timestamp 1666464484
transform 1 0 58420 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1666464484
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666464484
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666464484
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666464484
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666464484
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666464484
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666464484
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666464484
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1666464484
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1666464484
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1666464484
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1666464484
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1666464484
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1666464484
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1666464484
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1666464484
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666464484
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666464484
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666464484
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666464484
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666464484
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666464484
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666464484
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1666464484
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1666464484
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1666464484
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1666464484
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1666464484
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1666464484
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1666464484
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666464484
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666464484
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666464484
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666464484
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666464484
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666464484
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666464484
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1666464484
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1666464484
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1666464484
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1666464484
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1666464484
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666464484
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666464484
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1666464484
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1666464484
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1666464484
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666464484
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1666464484
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1666464484
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1666464484
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666464484
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666464484
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1666464484
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1666464484
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1666464484
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1666464484
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666464484
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666464484
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666464484
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666464484
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666464484
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1666464484
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1666464484
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1666464484
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666464484
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666464484
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666464484
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666464484
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666464484
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666464484
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666464484
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666464484
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1666464484
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1666464484
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1666464484
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666464484
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666464484
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666464484
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666464484
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666464484
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666464484
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1666464484
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1666464484
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1666464484
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1666464484
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_21
timestamp 1666464484
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1666464484
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_45
timestamp 1666464484
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666464484
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666464484
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666464484
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_425
timestamp 1666464484
transform 1 0 40204 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1666464484
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_456
timestamp 1666464484
transform 1 0 43056 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_468
timestamp 1666464484
transform 1 0 44160 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_480
timestamp 1666464484
transform 1 0 45264 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_492
timestamp 1666464484
transform 1 0 46368 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1666464484
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1666464484
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1666464484
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1666464484
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_38
timestamp 1666464484
transform 1 0 4600 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_63
timestamp 1666464484
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1666464484
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666464484
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666464484
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666464484
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666464484
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666464484
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_445
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_449
timestamp 1666464484
transform 1 0 42412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_466
timestamp 1666464484
transform 1 0 43976 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1666464484
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_495
timestamp 1666464484
transform 1 0 46644 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_507
timestamp 1666464484
transform 1 0 47748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_519
timestamp 1666464484
transform 1 0 48852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1666464484
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1666464484
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1666464484
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1666464484
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1666464484
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_65
timestamp 1666464484
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_71
timestamp 1666464484
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_79
timestamp 1666464484
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_91
timestamp 1666464484
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_103
timestamp 1666464484
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_118
timestamp 1666464484
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_130
timestamp 1666464484
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_142
timestamp 1666464484
transform 1 0 14168 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_154
timestamp 1666464484
transform 1 0 15272 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666464484
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666464484
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666464484
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666464484
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_417
timestamp 1666464484
transform 1 0 39468 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_423
timestamp 1666464484
transform 1 0 40020 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1666464484
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_439
timestamp 1666464484
transform 1 0 41492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1666464484
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_467
timestamp 1666464484
transform 1 0 44068 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_487
timestamp 1666464484
transform 1 0 45908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1666464484
transform 1 0 47012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1666464484
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1666464484
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1666464484
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1666464484
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1666464484
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1666464484
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1666464484
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_210
timestamp 1666464484
transform 1 0 20424 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_222
timestamp 1666464484
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_234
timestamp 1666464484
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1666464484
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666464484
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666464484
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1666464484
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1666464484
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_439
timestamp 1666464484
transform 1 0 41492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_462
timestamp 1666464484
transform 1 0 43608 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_472
timestamp 1666464484
transform 1 0 44528 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1666464484
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1666464484
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1666464484
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_33
timestamp 1666464484
transform 1 0 4140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_37
timestamp 1666464484
transform 1 0 4508 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_41
timestamp 1666464484
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1666464484
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_61
timestamp 1666464484
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1666464484
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1666464484
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_95
timestamp 1666464484
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1666464484
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_133
timestamp 1666464484
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_145
timestamp 1666464484
transform 1 0 14444 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_157
timestamp 1666464484
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1666464484
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666464484
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666464484
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666464484
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_408
timestamp 1666464484
transform 1 0 38640 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_428
timestamp 1666464484
transform 1 0 40480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_438
timestamp 1666464484
transform 1 0 41400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1666464484
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_454
timestamp 1666464484
transform 1 0 42872 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1666464484
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_34
timestamp 1666464484
transform 1 0 4232 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_46
timestamp 1666464484
transform 1 0 5336 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1666464484
transform 1 0 6440 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_94
timestamp 1666464484
transform 1 0 9752 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_118
timestamp 1666464484
transform 1 0 11960 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1666464484
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666464484
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1666464484
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_407
timestamp 1666464484
transform 1 0 38548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_411
timestamp 1666464484
transform 1 0 38916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1666464484
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_433
timestamp 1666464484
transform 1 0 40940 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_455
timestamp 1666464484
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_467
timestamp 1666464484
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1666464484
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1666464484
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_35
timestamp 1666464484
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1666464484
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1666464484
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1666464484
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1666464484
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1666464484
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_92
timestamp 1666464484
transform 1 0 9568 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_100
timestamp 1666464484
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1666464484
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1666464484
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_129
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_141
timestamp 1666464484
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1666464484
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1666464484
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666464484
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666464484
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666464484
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_405
timestamp 1666464484
transform 1 0 38364 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666464484
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_460
timestamp 1666464484
transform 1 0 43424 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_469
timestamp 1666464484
transform 1 0 44252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_481
timestamp 1666464484
transform 1 0 45356 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_493
timestamp 1666464484
transform 1 0 46460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_501
timestamp 1666464484
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1666464484
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1666464484
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_60
timestamp 1666464484
transform 1 0 6624 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 1666464484
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1666464484
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1666464484
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 1666464484
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1666464484
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_175
timestamp 1666464484
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1666464484
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_220
timestamp 1666464484
transform 1 0 21344 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_232
timestamp 1666464484
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1666464484
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666464484
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666464484
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666464484
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666464484
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666464484
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_426
timestamp 1666464484
transform 1 0 40296 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_438
timestamp 1666464484
transform 1 0 41400 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_450
timestamp 1666464484
transform 1 0 42504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_454
timestamp 1666464484
transform 1 0 42872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_471
timestamp 1666464484
transform 1 0 44436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1666464484
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1666464484
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1666464484
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1666464484
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1666464484
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_85
timestamp 1666464484
transform 1 0 8924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_97
timestamp 1666464484
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1666464484
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_140
timestamp 1666464484
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_152
timestamp 1666464484
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1666464484
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1666464484
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1666464484
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1666464484
transform 1 0 20516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666464484
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666464484
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666464484
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666464484
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666464484
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_417
timestamp 1666464484
transform 1 0 39468 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_439
timestamp 1666464484
transform 1 0 41492 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_457
timestamp 1666464484
transform 1 0 43148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_476
timestamp 1666464484
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_486
timestamp 1666464484
transform 1 0 45816 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_498
timestamp 1666464484
transform 1 0 46920 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1666464484
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1666464484
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1666464484
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1666464484
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_51
timestamp 1666464484
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_63
timestamp 1666464484
transform 1 0 6900 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1666464484
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1666464484
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_92
timestamp 1666464484
transform 1 0 9568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1666464484
transform 1 0 10672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1666464484
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1666464484
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_146
timestamp 1666464484
transform 1 0 14536 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1666464484
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_190
timestamp 1666464484
transform 1 0 18584 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1666464484
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1666464484
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_231
timestamp 1666464484
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1666464484
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666464484
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666464484
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666464484
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666464484
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666464484
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666464484
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666464484
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_439
timestamp 1666464484
transform 1 0 41492 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_451
timestamp 1666464484
transform 1 0 42596 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1666464484
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_482
timestamp 1666464484
transform 1 0 45448 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666464484
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1666464484
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1666464484
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1666464484
transform 1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1666464484
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1666464484
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_100
timestamp 1666464484
transform 1 0 10304 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_120
timestamp 1666464484
transform 1 0 12144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1666464484
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_150
timestamp 1666464484
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1666464484
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1666464484
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_207
timestamp 1666464484
transform 1 0 20148 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1666464484
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_243
timestamp 1666464484
transform 1 0 23460 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_255
timestamp 1666464484
transform 1 0 24564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_267
timestamp 1666464484
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666464484
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666464484
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666464484
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666464484
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666464484
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_405
timestamp 1666464484
transform 1 0 38364 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_413
timestamp 1666464484
transform 1 0 39100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_431
timestamp 1666464484
transform 1 0 40756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 1666464484
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1666464484
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_461
timestamp 1666464484
transform 1 0 43516 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_480
timestamp 1666464484
transform 1 0 45264 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_492
timestamp 1666464484
transform 1 0 46368 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1666464484
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_103
timestamp 1666464484
transform 1 0 10580 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_115
timestamp 1666464484
transform 1 0 11684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_127
timestamp 1666464484
transform 1 0 12788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1666464484
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_168
timestamp 1666464484
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_180
timestamp 1666464484
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1666464484
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1666464484
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_216
timestamp 1666464484
transform 1 0 20976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_224
timestamp 1666464484
transform 1 0 21712 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1666464484
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_237
timestamp 1666464484
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1666464484
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666464484
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666464484
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666464484
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666464484
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666464484
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_413
timestamp 1666464484
transform 1 0 39100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1666464484
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_439
timestamp 1666464484
transform 1 0 41492 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_449
timestamp 1666464484
transform 1 0 42412 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_461
timestamp 1666464484
transform 1 0 43516 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_466
timestamp 1666464484
transform 1 0 43976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1666464484
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666464484
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666464484
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1666464484
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1666464484
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_86
timestamp 1666464484
transform 1 0 9016 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_98
timestamp 1666464484
transform 1 0 10120 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1666464484
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1666464484
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_174
timestamp 1666464484
transform 1 0 17112 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_186
timestamp 1666464484
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_198
timestamp 1666464484
transform 1 0 19320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1666464484
transform 1 0 19780 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_210
timestamp 1666464484
transform 1 0 20424 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1666464484
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666464484
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666464484
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666464484
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666464484
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_417
timestamp 1666464484
transform 1 0 39468 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_421
timestamp 1666464484
transform 1 0 39836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_425
timestamp 1666464484
transform 1 0 40204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_432
timestamp 1666464484
transform 1 0 40848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_438
timestamp 1666464484
transform 1 0 41400 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1666464484
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_461
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_483
timestamp 1666464484
transform 1 0 45540 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_495
timestamp 1666464484
transform 1 0 46644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1666464484
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_34
timestamp 1666464484
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1666464484
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1666464484
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1666464484
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1666464484
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_169
timestamp 1666464484
transform 1 0 16652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_181
timestamp 1666464484
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1666464484
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1666464484
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_224
timestamp 1666464484
transform 1 0 21712 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_236
timestamp 1666464484
transform 1 0 22816 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1666464484
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666464484
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666464484
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666464484
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666464484
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666464484
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666464484
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666464484
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_429
timestamp 1666464484
transform 1 0 40572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_434
timestamp 1666464484
transform 1 0 41032 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_458
timestamp 1666464484
transform 1 0 43240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_470
timestamp 1666464484
transform 1 0 44344 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1666464484
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_495
timestamp 1666464484
transform 1 0 46644 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_507
timestamp 1666464484
transform 1 0 47748 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_519
timestamp 1666464484
transform 1 0 48852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1666464484
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1666464484
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_12
timestamp 1666464484
transform 1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_32
timestamp 1666464484
transform 1 0 4048 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_61
timestamp 1666464484
transform 1 0 6716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_73
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1666464484
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_143
timestamp 1666464484
transform 1 0 14260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1666464484
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_189
timestamp 1666464484
transform 1 0 18492 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_201
timestamp 1666464484
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1666464484
transform 1 0 20700 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1666464484
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_232
timestamp 1666464484
transform 1 0 22448 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_244
timestamp 1666464484
transform 1 0 23552 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_256
timestamp 1666464484
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1666464484
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666464484
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666464484
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666464484
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_411
timestamp 1666464484
transform 1 0 38916 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_423
timestamp 1666464484
transform 1 0 40020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666464484
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666464484
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_467
timestamp 1666464484
transform 1 0 44068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_487
timestamp 1666464484
transform 1 0 45908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666464484
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1666464484
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1666464484
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1666464484
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_75
timestamp 1666464484
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_150
timestamp 1666464484
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_162
timestamp 1666464484
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1666464484
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1666464484
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1666464484
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1666464484
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_238
timestamp 1666464484
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1666464484
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666464484
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666464484
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1666464484
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1666464484
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_402
timestamp 1666464484
transform 1 0 38088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1666464484
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_431
timestamp 1666464484
transform 1 0 40756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_455
timestamp 1666464484
transform 1 0 42964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_465
timestamp 1666464484
transform 1 0 43884 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1666464484
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_482
timestamp 1666464484
transform 1 0 45448 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_494
timestamp 1666464484
transform 1 0 46552 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_506
timestamp 1666464484
transform 1 0 47656 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_518
timestamp 1666464484
transform 1 0 48760 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_530
timestamp 1666464484
transform 1 0 49864 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1666464484
transform 1 0 4232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_50
timestamp 1666464484
transform 1 0 5704 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1666464484
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1666464484
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_82
timestamp 1666464484
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_94
timestamp 1666464484
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1666464484
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1666464484
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_198
timestamp 1666464484
transform 1 0 19320 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1666464484
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_231
timestamp 1666464484
transform 1 0 22356 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_243
timestamp 1666464484
transform 1 0 23460 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_255
timestamp 1666464484
transform 1 0 24564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_267
timestamp 1666464484
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666464484
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666464484
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666464484
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_385
timestamp 1666464484
transform 1 0 36524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_411
timestamp 1666464484
transform 1 0 38916 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_418
timestamp 1666464484
transform 1 0 39560 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_422
timestamp 1666464484
transform 1 0 39928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_426
timestamp 1666464484
transform 1 0 40296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1666464484
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_457
timestamp 1666464484
transform 1 0 43148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_465
timestamp 1666464484
transform 1 0 43884 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_484
timestamp 1666464484
transform 1 0 45632 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_496
timestamp 1666464484
transform 1 0 46736 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1666464484
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1666464484
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1666464484
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1666464484
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_37
timestamp 1666464484
transform 1 0 4508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_52
timestamp 1666464484
transform 1 0 5888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_60
timestamp 1666464484
transform 1 0 6624 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_69
timestamp 1666464484
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1666464484
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1666464484
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1666464484
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_186
timestamp 1666464484
transform 1 0 18216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1666464484
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_218
timestamp 1666464484
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_230
timestamp 1666464484
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1666464484
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666464484
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666464484
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666464484
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666464484
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666464484
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666464484
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666464484
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666464484
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_392
timestamp 1666464484
transform 1 0 37168 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_412
timestamp 1666464484
transform 1 0 39008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_429
timestamp 1666464484
transform 1 0 40572 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_446
timestamp 1666464484
transform 1 0 42136 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_458
timestamp 1666464484
transform 1 0 43240 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_470
timestamp 1666464484
transform 1 0 44344 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1666464484
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1666464484
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1666464484
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_18
timestamp 1666464484
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_30
timestamp 1666464484
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_42
timestamp 1666464484
transform 1 0 4968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_50
timestamp 1666464484
transform 1 0 5704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1666464484
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_75
timestamp 1666464484
transform 1 0 8004 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_87
timestamp 1666464484
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_99
timestamp 1666464484
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_180
timestamp 1666464484
transform 1 0 17664 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 1666464484
transform 1 0 18400 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_209
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1666464484
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666464484
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666464484
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666464484
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_355
timestamp 1666464484
transform 1 0 33764 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_367
timestamp 1666464484
transform 1 0 34868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_379
timestamp 1666464484
transform 1 0 35972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_402
timestamp 1666464484
transform 1 0 38088 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_414
timestamp 1666464484
transform 1 0 39192 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_426
timestamp 1666464484
transform 1 0 40296 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_432
timestamp 1666464484
transform 1 0 40848 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_436
timestamp 1666464484
transform 1 0 41216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_443
timestamp 1666464484
transform 1 0 41860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666464484
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666464484
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666464484
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666464484
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666464484
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1666464484
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1666464484
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1666464484
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_159
timestamp 1666464484
transform 1 0 15732 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_167
timestamp 1666464484
transform 1 0 16468 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1666464484
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1666464484
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1666464484
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_223
timestamp 1666464484
transform 1 0 21620 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_235
timestamp 1666464484
transform 1 0 22724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1666464484
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1666464484
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1666464484
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_315
timestamp 1666464484
transform 1 0 30084 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_322
timestamp 1666464484
transform 1 0 30728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_334
timestamp 1666464484
transform 1 0 31832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_338
timestamp 1666464484
transform 1 0 32200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_346
timestamp 1666464484
transform 1 0 32936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1666464484
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_370
timestamp 1666464484
transform 1 0 35144 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_382
timestamp 1666464484
transform 1 0 36248 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_394
timestamp 1666464484
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_406
timestamp 1666464484
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1666464484
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666464484
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666464484
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666464484
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666464484
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666464484
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666464484
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1666464484
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1666464484
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1666464484
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_12
timestamp 1666464484
transform 1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1666464484
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_129
timestamp 1666464484
transform 1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1666464484
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_187
timestamp 1666464484
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_191
timestamp 1666464484
transform 1 0 18676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_198
timestamp 1666464484
transform 1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_289
timestamp 1666464484
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_308
timestamp 1666464484
transform 1 0 29440 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_312
timestamp 1666464484
transform 1 0 29808 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_341
timestamp 1666464484
transform 1 0 32476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_358
timestamp 1666464484
transform 1 0 34040 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_380
timestamp 1666464484
transform 1 0 36064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1666464484
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1666464484
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_401
timestamp 1666464484
transform 1 0 37996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_419
timestamp 1666464484
transform 1 0 39652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1666464484
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1666464484
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666464484
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666464484
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666464484
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1666464484
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1666464484
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1666464484
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1666464484
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1666464484
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_37
timestamp 1666464484
transform 1 0 4508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_49
timestamp 1666464484
transform 1 0 5612 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_61
timestamp 1666464484
transform 1 0 6716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 1666464484
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1666464484
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1666464484
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_146
timestamp 1666464484
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_158
timestamp 1666464484
transform 1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_166
timestamp 1666464484
transform 1 0 16376 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1666464484
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1666464484
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_204
timestamp 1666464484
transform 1 0 19872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1666464484
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1666464484
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1666464484
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1666464484
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_355
timestamp 1666464484
transform 1 0 33764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1666464484
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_383
timestamp 1666464484
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_390
timestamp 1666464484
transform 1 0 36984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_399
timestamp 1666464484
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_410
timestamp 1666464484
transform 1 0 38824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1666464484
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_427
timestamp 1666464484
transform 1 0 40388 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_444
timestamp 1666464484
transform 1 0 41952 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_464
timestamp 1666464484
transform 1 0 43792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666464484
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666464484
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1666464484
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1666464484
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1666464484
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1666464484
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1666464484
transform 1 0 2208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_36
timestamp 1666464484
transform 1 0 4416 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1666464484
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1666464484
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_197
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_230
timestamp 1666464484
transform 1 0 22264 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_242
timestamp 1666464484
transform 1 0 23368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_254
timestamp 1666464484
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1666464484
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1666464484
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_298
timestamp 1666464484
transform 1 0 28520 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1666464484
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_328
timestamp 1666464484
transform 1 0 31280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1666464484
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_342
timestamp 1666464484
transform 1 0 32568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_350
timestamp 1666464484
transform 1 0 33304 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1666464484
transform 1 0 34868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_377
timestamp 1666464484
transform 1 0 35788 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_383
timestamp 1666464484
transform 1 0 36340 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_411
timestamp 1666464484
transform 1 0 38916 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_431
timestamp 1666464484
transform 1 0 40756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1666464484
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1666464484
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_467
timestamp 1666464484
transform 1 0 44068 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_479
timestamp 1666464484
transform 1 0 45172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_491
timestamp 1666464484
transform 1 0 46276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1666464484
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_9
timestamp 1666464484
transform 1 0 1932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_17
timestamp 1666464484
transform 1 0 2668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1666464484
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_35
timestamp 1666464484
transform 1 0 4324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_38
timestamp 1666464484
transform 1 0 4600 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_50
timestamp 1666464484
transform 1 0 5704 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_62
timestamp 1666464484
transform 1 0 6808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1666464484
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_129
timestamp 1666464484
transform 1 0 12972 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1666464484
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_145
timestamp 1666464484
transform 1 0 14444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_157
timestamp 1666464484
transform 1 0 15548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_169
timestamp 1666464484
transform 1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1666464484
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1666464484
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1666464484
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_219
timestamp 1666464484
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1666464484
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666464484
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666464484
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666464484
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666464484
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666464484
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_348
timestamp 1666464484
transform 1 0 33120 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1666464484
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_377
timestamp 1666464484
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_397
timestamp 1666464484
transform 1 0 37628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_406
timestamp 1666464484
transform 1 0 38456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_415
timestamp 1666464484
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666464484
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_429
timestamp 1666464484
transform 1 0 40572 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_433
timestamp 1666464484
transform 1 0 40940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_453
timestamp 1666464484
transform 1 0 42780 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_463
timestamp 1666464484
transform 1 0 43700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666464484
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666464484
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666464484
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1666464484
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1666464484
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1666464484
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1666464484
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1666464484
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1666464484
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1666464484
transform 1 0 12052 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1666464484
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1666464484
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1666464484
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_186
timestamp 1666464484
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_198
timestamp 1666464484
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1666464484
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666464484
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666464484
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666464484
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_402
timestamp 1666464484
transform 1 0 38088 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_414
timestamp 1666464484
transform 1 0 39192 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_426
timestamp 1666464484
transform 1 0 40296 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_438
timestamp 1666464484
transform 1 0 41400 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1666464484
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666464484
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_454
timestamp 1666464484
transform 1 0 42872 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_466
timestamp 1666464484
transform 1 0 43976 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_478
timestamp 1666464484
transform 1 0 45080 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_490
timestamp 1666464484
transform 1 0 46184 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1666464484
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1666464484
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1666464484
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1666464484
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1666464484
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1666464484
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1666464484
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_150
timestamp 1666464484
transform 1 0 14904 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1666464484
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1666464484
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_271
timestamp 1666464484
transform 1 0 26036 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_283
timestamp 1666464484
transform 1 0 27140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_295
timestamp 1666464484
transform 1 0 28244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666464484
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_327
timestamp 1666464484
transform 1 0 31188 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_339
timestamp 1666464484
transform 1 0 32292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_351
timestamp 1666464484
transform 1 0 33396 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1666464484
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_377
timestamp 1666464484
transform 1 0 35788 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_386
timestamp 1666464484
transform 1 0 36616 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_398
timestamp 1666464484
transform 1 0 37720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_410
timestamp 1666464484
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1666464484
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_426
timestamp 1666464484
transform 1 0 40296 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_438
timestamp 1666464484
transform 1 0 41400 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_450
timestamp 1666464484
transform 1 0 42504 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_462
timestamp 1666464484
transform 1 0 43608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1666464484
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1666464484
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1666464484
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1666464484
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1666464484
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1666464484
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_120
timestamp 1666464484
transform 1 0 12144 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_128
timestamp 1666464484
transform 1 0 12880 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1666464484
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_199
timestamp 1666464484
transform 1 0 19412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_211
timestamp 1666464484
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_242
timestamp 1666464484
transform 1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1666464484
transform 1 0 25208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1666464484
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1666464484
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_309
timestamp 1666464484
transform 1 0 29532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_313
timestamp 1666464484
transform 1 0 29900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1666464484
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_365
timestamp 1666464484
transform 1 0 34684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_373
timestamp 1666464484
transform 1 0 35420 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1666464484
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_415
timestamp 1666464484
transform 1 0 39284 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_439
timestamp 1666464484
transform 1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666464484
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_456
timestamp 1666464484
transform 1 0 43056 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_468
timestamp 1666464484
transform 1 0 44160 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_480
timestamp 1666464484
transform 1 0 45264 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_492
timestamp 1666464484
transform 1 0 46368 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1666464484
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1666464484
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1666464484
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_128
timestamp 1666464484
transform 1 0 12880 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1666464484
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_163
timestamp 1666464484
transform 1 0 16100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1666464484
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_229
timestamp 1666464484
transform 1 0 22172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_237
timestamp 1666464484
transform 1 0 22908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_241
timestamp 1666464484
transform 1 0 23276 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1666464484
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_271
timestamp 1666464484
transform 1 0 26036 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_283
timestamp 1666464484
transform 1 0 27140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_295
timestamp 1666464484
transform 1 0 28244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1666464484
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_329
timestamp 1666464484
transform 1 0 31372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_339
timestamp 1666464484
transform 1 0 32292 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_345
timestamp 1666464484
transform 1 0 32844 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1666464484
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_372
timestamp 1666464484
transform 1 0 35328 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_400
timestamp 1666464484
transform 1 0 37904 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_406
timestamp 1666464484
transform 1 0 38456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1666464484
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_435
timestamp 1666464484
transform 1 0 41124 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_459
timestamp 1666464484
transform 1 0 43332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1666464484
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666464484
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1666464484
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1666464484
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1666464484
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1666464484
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1666464484
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_130
timestamp 1666464484
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_134
timestamp 1666464484
transform 1 0 13432 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1666464484
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_143
timestamp 1666464484
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_156
timestamp 1666464484
transform 1 0 15456 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1666464484
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1666464484
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1666464484
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_241
timestamp 1666464484
transform 1 0 23276 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_265
timestamp 1666464484
transform 1 0 25484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1666464484
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_311
timestamp 1666464484
transform 1 0 29716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_343
timestamp 1666464484
transform 1 0 32660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_347
timestamp 1666464484
transform 1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_367
timestamp 1666464484
transform 1 0 34868 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_373
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1666464484
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_400
timestamp 1666464484
transform 1 0 37904 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_420
timestamp 1666464484
transform 1 0 39744 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_440
timestamp 1666464484
transform 1 0 41584 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_460
timestamp 1666464484
transform 1 0 43424 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_470
timestamp 1666464484
transform 1 0 44344 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_482
timestamp 1666464484
transform 1 0 45448 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_494
timestamp 1666464484
transform 1 0 46552 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1666464484
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1666464484
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1666464484
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1666464484
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_129
timestamp 1666464484
transform 1 0 12972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1666464484
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_148
timestamp 1666464484
transform 1 0 14720 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_160
timestamp 1666464484
transform 1 0 15824 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_172
timestamp 1666464484
transform 1 0 16928 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_205
timestamp 1666464484
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1666464484
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_230
timestamp 1666464484
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1666464484
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1666464484
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_258
timestamp 1666464484
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_270
timestamp 1666464484
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_282
timestamp 1666464484
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1666464484
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1666464484
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_324
timestamp 1666464484
transform 1 0 30912 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_336
timestamp 1666464484
transform 1 0 32016 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_344
timestamp 1666464484
transform 1 0 32752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_353
timestamp 1666464484
transform 1 0 33580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1666464484
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 1666464484
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_385
timestamp 1666464484
transform 1 0 36524 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_392
timestamp 1666464484
transform 1 0 37168 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_404
timestamp 1666464484
transform 1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_410
timestamp 1666464484
transform 1 0 38824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_414
timestamp 1666464484
transform 1 0 39192 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1666464484
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_439
timestamp 1666464484
transform 1 0 41492 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_451
timestamp 1666464484
transform 1 0 42596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_468
timestamp 1666464484
transform 1 0 44160 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666464484
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1666464484
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1666464484
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1666464484
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_144
timestamp 1666464484
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_156
timestamp 1666464484
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_175
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_179
timestamp 1666464484
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_199
timestamp 1666464484
transform 1 0 19412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_214
timestamp 1666464484
transform 1 0 20792 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1666464484
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_233
timestamp 1666464484
transform 1 0 22540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1666464484
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1666464484
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_266
timestamp 1666464484
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1666464484
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_289
timestamp 1666464484
transform 1 0 27692 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_306
timestamp 1666464484
transform 1 0 29256 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_310
timestamp 1666464484
transform 1 0 29624 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666464484
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1666464484
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_342
timestamp 1666464484
transform 1 0 32568 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_348
timestamp 1666464484
transform 1 0 33120 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_355
timestamp 1666464484
transform 1 0 33764 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_367
timestamp 1666464484
transform 1 0 34868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_379
timestamp 1666464484
transform 1 0 35972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_417
timestamp 1666464484
transform 1 0 39468 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_425
timestamp 1666464484
transform 1 0 40204 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666464484
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_441
timestamp 1666464484
transform 1 0 41676 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1666464484
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_455
timestamp 1666464484
transform 1 0 42964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_472
timestamp 1666464484
transform 1 0 44528 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_496
timestamp 1666464484
transform 1 0 46736 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1666464484
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1666464484
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1666464484
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_219
timestamp 1666464484
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_231
timestamp 1666464484
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1666464484
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_271
timestamp 1666464484
transform 1 0 26036 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_286
timestamp 1666464484
transform 1 0 27416 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1666464484
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_335
timestamp 1666464484
transform 1 0 31924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1666464484
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_405
timestamp 1666464484
transform 1 0 38364 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_412
timestamp 1666464484
transform 1 0 39008 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_461
timestamp 1666464484
transform 1 0 43516 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666464484
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666464484
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1666464484
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_187
timestamp 1666464484
transform 1 0 18308 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1666464484
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1666464484
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1666464484
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_251
timestamp 1666464484
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_271
timestamp 1666464484
transform 1 0 26036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1666464484
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_288
timestamp 1666464484
transform 1 0 27600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_308
timestamp 1666464484
transform 1 0 29440 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_316
timestamp 1666464484
transform 1 0 30176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1666464484
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_355
timestamp 1666464484
transform 1 0 33764 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1666464484
transform 1 0 34868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_371
timestamp 1666464484
transform 1 0 35236 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1666464484
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_397
timestamp 1666464484
transform 1 0 37628 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_401
timestamp 1666464484
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_421
timestamp 1666464484
transform 1 0 39836 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_431
timestamp 1666464484
transform 1 0 40756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_443
timestamp 1666464484
transform 1 0 41860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_460
timestamp 1666464484
transform 1 0 43424 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_471
timestamp 1666464484
transform 1 0 44436 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_483
timestamp 1666464484
transform 1 0 45540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_495
timestamp 1666464484
transform 1 0 46644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1666464484
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1666464484
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1666464484
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1666464484
transform 1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_229
timestamp 1666464484
transform 1 0 22172 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_237
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_243
timestamp 1666464484
transform 1 0 23460 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1666464484
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_271
timestamp 1666464484
transform 1 0 26036 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_283
timestamp 1666464484
transform 1 0 27140 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1666464484
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_328
timestamp 1666464484
transform 1 0 31280 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_348
timestamp 1666464484
transform 1 0 33120 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1666464484
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 1666464484
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_386
timestamp 1666464484
transform 1 0 36616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_393
timestamp 1666464484
transform 1 0 37260 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1666464484
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_439
timestamp 1666464484
transform 1 0 41492 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_447
timestamp 1666464484
transform 1 0 42228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_466
timestamp 1666464484
transform 1 0 43976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1666464484
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_482
timestamp 1666464484
transform 1 0 45448 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_494
timestamp 1666464484
transform 1 0 46552 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_506
timestamp 1666464484
transform 1 0 47656 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_518
timestamp 1666464484
transform 1 0 48760 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_530
timestamp 1666464484
transform 1 0 49864 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1666464484
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_175
timestamp 1666464484
transform 1 0 17204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_179
timestamp 1666464484
transform 1 0 17572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 1666464484
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1666464484
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_210
timestamp 1666464484
transform 1 0 20424 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_216
timestamp 1666464484
transform 1 0 20976 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1666464484
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_233
timestamp 1666464484
transform 1 0 22540 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_238
timestamp 1666464484
transform 1 0 23000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_262
timestamp 1666464484
transform 1 0 25208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1666464484
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1666464484
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_302
timestamp 1666464484
transform 1 0 28888 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_314
timestamp 1666464484
transform 1 0 29992 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_326
timestamp 1666464484
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1666464484
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_342
timestamp 1666464484
transform 1 0 32568 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_365
timestamp 1666464484
transform 1 0 34684 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_401
timestamp 1666464484
transform 1 0 37996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_421
timestamp 1666464484
transform 1 0 39836 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_428
timestamp 1666464484
transform 1 0 40480 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_440
timestamp 1666464484
transform 1 0 41584 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1666464484
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_467
timestamp 1666464484
transform 1 0 44068 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_475
timestamp 1666464484
transform 1 0 44804 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_481
timestamp 1666464484
transform 1 0 45356 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_493
timestamp 1666464484
transform 1 0 46460 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_501
timestamp 1666464484
transform 1 0 47196 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1666464484
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1666464484
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1666464484
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_258
timestamp 1666464484
transform 1 0 24840 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_270
timestamp 1666464484
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_282
timestamp 1666464484
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_294
timestamp 1666464484
transform 1 0 28152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1666464484
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1666464484
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1666464484
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1666464484
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_387
timestamp 1666464484
transform 1 0 36708 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_399
timestamp 1666464484
transform 1 0 37812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_407
timestamp 1666464484
transform 1 0 38548 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_412
timestamp 1666464484
transform 1 0 39008 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_459
timestamp 1666464484
transform 1 0 43332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_467
timestamp 1666464484
transform 1 0 44068 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_474
timestamp 1666464484
transform 1 0 44712 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_495
timestamp 1666464484
transform 1 0 46644 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_507
timestamp 1666464484
transform 1 0 47748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_519
timestamp 1666464484
transform 1 0 48852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_175
timestamp 1666464484
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_179
timestamp 1666464484
transform 1 0 17572 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_190
timestamp 1666464484
transform 1 0 18584 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_202
timestamp 1666464484
transform 1 0 19688 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1666464484
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1666464484
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_257
timestamp 1666464484
transform 1 0 24748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_269
timestamp 1666464484
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1666464484
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_313
timestamp 1666464484
transform 1 0 29900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1666464484
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_377
timestamp 1666464484
transform 1 0 35788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1666464484
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_411
timestamp 1666464484
transform 1 0 38916 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_423
timestamp 1666464484
transform 1 0 40020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_435
timestamp 1666464484
transform 1 0 41124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_453
timestamp 1666464484
transform 1 0 42780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_457
timestamp 1666464484
transform 1 0 43148 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_466
timestamp 1666464484
transform 1 0 43976 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_476
timestamp 1666464484
transform 1 0 44896 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_492
timestamp 1666464484
transform 1 0 46368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1666464484
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1666464484
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1666464484
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1666464484
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_225
timestamp 1666464484
transform 1 0 21804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1666464484
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1666464484
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_261
timestamp 1666464484
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_273
timestamp 1666464484
transform 1 0 26220 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_285
timestamp 1666464484
transform 1 0 27324 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1666464484
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1666464484
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_317
timestamp 1666464484
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_473
timestamp 1666464484
transform 1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_495
timestamp 1666464484
transform 1 0 46644 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_507
timestamp 1666464484
transform 1 0 47748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_519
timestamp 1666464484
transform 1 0 48852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1666464484
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_233
timestamp 1666464484
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1666464484
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_264
timestamp 1666464484
transform 1 0 25392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1666464484
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1666464484
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_342
timestamp 1666464484
transform 1 0 32568 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_354
timestamp 1666464484
transform 1 0 33672 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_382
timestamp 1666464484
transform 1 0 36248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1666464484
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_459
timestamp 1666464484
transform 1 0 43332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_471
timestamp 1666464484
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_483
timestamp 1666464484
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_495
timestamp 1666464484
transform 1 0 46644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_241
timestamp 1666464484
transform 1 0 23276 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1666464484
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666464484
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_317
timestamp 1666464484
transform 1 0 30268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_336
timestamp 1666464484
transform 1 0 32016 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_346
timestamp 1666464484
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1666464484
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_383
timestamp 1666464484
transform 1 0 36340 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_395
timestamp 1666464484
transform 1 0 37444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_407
timestamp 1666464484
transform 1 0 38548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_467
timestamp 1666464484
transform 1 0 44068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_473
timestamp 1666464484
transform 1 0 44620 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_237
timestamp 1666464484
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_256
timestamp 1666464484
transform 1 0 24656 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_268
timestamp 1666464484
transform 1 0 25760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_326
timestamp 1666464484
transform 1 0 31096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1666464484
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_341
timestamp 1666464484
transform 1 0 32476 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_365
timestamp 1666464484
transform 1 0 34684 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_446
timestamp 1666464484
transform 1 0 42136 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_465
timestamp 1666464484
transform 1 0 43884 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_489
timestamp 1666464484
transform 1 0 46092 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_501
timestamp 1666464484
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_285
timestamp 1666464484
transform 1 0 27324 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1666464484
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1666464484
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_383
timestamp 1666464484
transform 1 0 36340 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_390
timestamp 1666464484
transform 1 0 36984 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_402
timestamp 1666464484
transform 1 0 38088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_414
timestamp 1666464484
transform 1 0 39192 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_439
timestamp 1666464484
transform 1 0 41492 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_456
timestamp 1666464484
transform 1 0 43056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_467
timestamp 1666464484
transform 1 0 44068 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_474
timestamp 1666464484
transform 1 0 44712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_484
timestamp 1666464484
transform 1 0 45632 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_491
timestamp 1666464484
transform 1 0 46276 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_503
timestamp 1666464484
transform 1 0 47380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_515
timestamp 1666464484
transform 1 0 48484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_527
timestamp 1666464484
transform 1 0 49588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_258
timestamp 1666464484
transform 1 0 24840 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_270
timestamp 1666464484
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1666464484
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_289
timestamp 1666464484
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666464484
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_317
timestamp 1666464484
transform 1 0 30268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_325
timestamp 1666464484
transform 1 0 31004 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_365
timestamp 1666464484
transform 1 0 34684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_369
timestamp 1666464484
transform 1 0 35052 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_381
timestamp 1666464484
transform 1 0 36156 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_387
timestamp 1666464484
transform 1 0 36708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1666464484
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_415
timestamp 1666464484
transform 1 0 39284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_421
timestamp 1666464484
transform 1 0 39836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_427
timestamp 1666464484
transform 1 0 40388 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_438
timestamp 1666464484
transform 1 0 41400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1666464484
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_457
timestamp 1666464484
transform 1 0 43148 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_468
timestamp 1666464484
transform 1 0 44160 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_476
timestamp 1666464484
transform 1 0 44896 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_494
timestamp 1666464484
transform 1 0 46552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1666464484
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1666464484
transform 1 0 26036 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1666464484
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_317
timestamp 1666464484
transform 1 0 30268 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_325
timestamp 1666464484
transform 1 0 31004 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_342
timestamp 1666464484
transform 1 0 32568 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_352
timestamp 1666464484
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_370
timestamp 1666464484
transform 1 0 35144 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_382
timestamp 1666464484
transform 1 0 36248 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_394
timestamp 1666464484
transform 1 0 37352 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_406
timestamp 1666464484
transform 1 0 38456 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1666464484
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_428
timestamp 1666464484
transform 1 0 40480 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_435
timestamp 1666464484
transform 1 0 41124 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_452
timestamp 1666464484
transform 1 0 42688 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_462
timestamp 1666464484
transform 1 0 43608 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_474
timestamp 1666464484
transform 1 0 44712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_484
timestamp 1666464484
transform 1 0 45632 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_496
timestamp 1666464484
transform 1 0 46736 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_508
timestamp 1666464484
transform 1 0 47840 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_520
timestamp 1666464484
transform 1 0 48944 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_230
timestamp 1666464484
transform 1 0 22264 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_242
timestamp 1666464484
transform 1 0 23368 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_268
timestamp 1666464484
transform 1 0 25760 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1666464484
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666464484
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_287
timestamp 1666464484
transform 1 0 27508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_307
timestamp 1666464484
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_314
timestamp 1666464484
transform 1 0 29992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1666464484
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_355
timestamp 1666464484
transform 1 0 33764 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_367
timestamp 1666464484
transform 1 0 34868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1666464484
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_424
timestamp 1666464484
transform 1 0 40112 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_444
timestamp 1666464484
transform 1 0 41952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_471
timestamp 1666464484
transform 1 0 44436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_483
timestamp 1666464484
transform 1 0 45540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_495
timestamp 1666464484
transform 1 0 46644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1666464484
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666464484
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_218
timestamp 1666464484
transform 1 0 21160 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_238
timestamp 1666464484
transform 1 0 23000 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_246
timestamp 1666464484
transform 1 0 23736 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1666464484
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1666464484
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_283
timestamp 1666464484
transform 1 0 27140 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_289
timestamp 1666464484
transform 1 0 27692 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1666464484
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_320
timestamp 1666464484
transform 1 0 30544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_340
timestamp 1666464484
transform 1 0 32384 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_350
timestamp 1666464484
transform 1 0 33304 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_356
timestamp 1666464484
transform 1 0 33856 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1666464484
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_397
timestamp 1666464484
transform 1 0 37628 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_404
timestamp 1666464484
transform 1 0 38272 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_412
timestamp 1666464484
transform 1 0 39008 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1666464484
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_430
timestamp 1666464484
transform 1 0 40664 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_437
timestamp 1666464484
transform 1 0 41308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_449
timestamp 1666464484
transform 1 0 42412 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_461
timestamp 1666464484
transform 1 0 43516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_473
timestamp 1666464484
transform 1 0 44620 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1666464484
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_243
timestamp 1666464484
transform 1 0 23460 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1666464484
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_297
timestamp 1666464484
transform 1 0 28428 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_304
timestamp 1666464484
transform 1 0 29072 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_316
timestamp 1666464484
transform 1 0 30176 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_331
timestamp 1666464484
transform 1 0 31556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_349
timestamp 1666464484
transform 1 0 33212 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_369
timestamp 1666464484
transform 1 0 35052 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_381
timestamp 1666464484
transform 1 0 36156 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_387
timestamp 1666464484
transform 1 0 36708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_401
timestamp 1666464484
transform 1 0 37996 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_413
timestamp 1666464484
transform 1 0 39100 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_425
timestamp 1666464484
transform 1 0 40204 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_437
timestamp 1666464484
transform 1 0 41308 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_445
timestamp 1666464484
transform 1 0 42044 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1666464484
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666464484
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666464484
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1666464484
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_235
timestamp 1666464484
transform 1 0 22724 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666464484
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_259
timestamp 1666464484
transform 1 0 24932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_276
timestamp 1666464484
transform 1 0 26496 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_283
timestamp 1666464484
transform 1 0 27140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_295
timestamp 1666464484
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_345
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1666464484
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_373
timestamp 1666464484
transform 1 0 35420 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_381
timestamp 1666464484
transform 1 0 36156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_398
timestamp 1666464484
transform 1 0 37720 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_405
timestamp 1666464484
transform 1 0 38364 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 1666464484
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_428
timestamp 1666464484
transform 1 0 40480 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_440
timestamp 1666464484
transform 1 0 41584 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_452
timestamp 1666464484
transform 1 0 42688 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_464
timestamp 1666464484
transform 1 0 43792 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666464484
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_230
timestamp 1666464484
transform 1 0 22264 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_242
timestamp 1666464484
transform 1 0 23368 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_254
timestamp 1666464484
transform 1 0 24472 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_272
timestamp 1666464484
transform 1 0 26128 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666464484
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_313
timestamp 1666464484
transform 1 0 29900 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_320
timestamp 1666464484
transform 1 0 30544 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1666464484
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_343
timestamp 1666464484
transform 1 0 32660 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_363
timestamp 1666464484
transform 1 0 34500 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_370
timestamp 1666464484
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_382
timestamp 1666464484
transform 1 0 36248 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1666464484
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_436
timestamp 1666464484
transform 1 0 41216 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1666464484
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1666464484
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1666464484
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666464484
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_245
timestamp 1666464484
transform 1 0 23644 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1666464484
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666464484
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_277
timestamp 1666464484
transform 1 0 26588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_281
timestamp 1666464484
transform 1 0 26956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_285
timestamp 1666464484
transform 1 0 27324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_297
timestamp 1666464484
transform 1 0 28428 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1666464484
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_327
timestamp 1666464484
transform 1 0 31188 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_334
timestamp 1666464484
transform 1 0 31832 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1666464484
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_397
timestamp 1666464484
transform 1 0 37628 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_409
timestamp 1666464484
transform 1 0 38732 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_417
timestamp 1666464484
transform 1 0 39468 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_431
timestamp 1666464484
transform 1 0 40756 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_443
timestamp 1666464484
transform 1 0 41860 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_455
timestamp 1666464484
transform 1 0 42964 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_467
timestamp 1666464484
transform 1 0 44068 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_120
timestamp 1666464484
transform 1 0 12144 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_132
timestamp 1666464484
transform 1 0 13248 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_144
timestamp 1666464484
transform 1 0 14352 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_156
timestamp 1666464484
transform 1 0 15456 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_233
timestamp 1666464484
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_239
timestamp 1666464484
transform 1 0 23092 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_259
timestamp 1666464484
transform 1 0 24932 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_271
timestamp 1666464484
transform 1 0 26036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1666464484
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_299
timestamp 1666464484
transform 1 0 28612 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_311
timestamp 1666464484
transform 1 0 29716 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1666464484
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_341
timestamp 1666464484
transform 1 0 32476 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_349
timestamp 1666464484
transform 1 0 33212 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_353
timestamp 1666464484
transform 1 0 33580 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_365
timestamp 1666464484
transform 1 0 34684 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_377
timestamp 1666464484
transform 1 0 35788 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1666464484
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_398
timestamp 1666464484
transform 1 0 37720 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_410
timestamp 1666464484
transform 1 0 38824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_414
timestamp 1666464484
transform 1 0 39192 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_420
timestamp 1666464484
transform 1 0 39744 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_431
timestamp 1666464484
transform 1 0 40756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_440
timestamp 1666464484
transform 1 0 41584 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666464484
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1666464484
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1666464484
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_47
timestamp 1666464484
transform 1 0 5428 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_64
timestamp 1666464484
transform 1 0 6992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1666464484
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_113
timestamp 1666464484
transform 1 0 11500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_130
timestamp 1666464484
transform 1 0 13064 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1666464484
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666464484
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1666464484
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_261
timestamp 1666464484
transform 1 0 25116 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_269
timestamp 1666464484
transform 1 0 25852 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1666464484
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_291
timestamp 1666464484
transform 1 0 27876 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1666464484
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1666464484
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_327
timestamp 1666464484
transform 1 0 31188 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_338
timestamp 1666464484
transform 1 0 32200 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1666464484
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1666464484
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_399
timestamp 1666464484
transform 1 0 37812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_409
timestamp 1666464484
transform 1 0 38732 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1666464484
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_439
timestamp 1666464484
transform 1 0 41492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_448
timestamp 1666464484
transform 1 0 42320 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_455
timestamp 1666464484
transform 1 0 42964 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_467
timestamp 1666464484
transform 1 0 44068 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666464484
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1666464484
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1666464484
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_77
timestamp 1666464484
transform 1 0 8188 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_89
timestamp 1666464484
transform 1 0 9292 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_110
timestamp 1666464484
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_120
timestamp 1666464484
transform 1 0 12144 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_140
timestamp 1666464484
transform 1 0 13984 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_152
timestamp 1666464484
transform 1 0 15088 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1666464484
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666464484
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_237
timestamp 1666464484
transform 1 0 22908 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_257
timestamp 1666464484
transform 1 0 24748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_269
timestamp 1666464484
transform 1 0 25852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 1666464484
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_288
timestamp 1666464484
transform 1 0 27600 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_297
timestamp 1666464484
transform 1 0 28428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_305
timestamp 1666464484
transform 1 0 29164 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_311
timestamp 1666464484
transform 1 0 29716 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_322
timestamp 1666464484
transform 1 0 30728 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1666464484
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_355
timestamp 1666464484
transform 1 0 33764 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_367
timestamp 1666464484
transform 1 0 34868 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1666464484
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_411
timestamp 1666464484
transform 1 0 38916 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_415
timestamp 1666464484
transform 1 0 39284 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_436
timestamp 1666464484
transform 1 0 41216 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_446
timestamp 1666464484
transform 1 0 42136 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1666464484
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1666464484
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1666464484
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_61
timestamp 1666464484
transform 1 0 6716 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 1666464484
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_106
timestamp 1666464484
transform 1 0 10856 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_126
timestamp 1666464484
transform 1 0 12696 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1666464484
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666464484
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666464484
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666464484
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_233
timestamp 1666464484
transform 1 0 22540 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_240
timestamp 1666464484
transform 1 0 23184 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1666464484
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666464484
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_265
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_274
timestamp 1666464484
transform 1 0 26312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_285
timestamp 1666464484
transform 1 0 27324 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_295
timestamp 1666464484
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1666464484
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1666464484
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_321
timestamp 1666464484
transform 1 0 30636 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_327
timestamp 1666464484
transform 1 0 31188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_331
timestamp 1666464484
transform 1 0 31556 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_335
timestamp 1666464484
transform 1 0 31924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_347
timestamp 1666464484
transform 1 0 33028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_359
timestamp 1666464484
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666464484
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_377
timestamp 1666464484
transform 1 0 35788 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_381
timestamp 1666464484
transform 1 0 36156 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666464484
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1666464484
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_426
timestamp 1666464484
transform 1 0 40296 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_446
timestamp 1666464484
transform 1 0 42136 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_450
timestamp 1666464484
transform 1 0 42504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_453
timestamp 1666464484
transform 1 0 42780 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_461
timestamp 1666464484
transform 1 0 43516 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_473
timestamp 1666464484
transform 1 0 44620 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1666464484
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_47
timestamp 1666464484
transform 1 0 5428 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1666464484
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_62
timestamp 1666464484
transform 1 0 6808 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_66
timestamp 1666464484
transform 1 0 7176 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_87
timestamp 1666464484
transform 1 0 9108 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_118
timestamp 1666464484
transform 1 0 11960 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_130
timestamp 1666464484
transform 1 0 13064 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_142
timestamp 1666464484
transform 1 0 14168 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_154
timestamp 1666464484
transform 1 0 15272 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1666464484
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666464484
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666464484
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_237
timestamp 1666464484
transform 1 0 22908 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_256
timestamp 1666464484
transform 1 0 24656 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_268
timestamp 1666464484
transform 1 0 25760 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_290
timestamp 1666464484
transform 1 0 27784 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_302
timestamp 1666464484
transform 1 0 28888 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_314
timestamp 1666464484
transform 1 0 29992 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_323
timestamp 1666464484
transform 1 0 30820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666464484
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666464484
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1666464484
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_436
timestamp 1666464484
transform 1 0 41216 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1666464484
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1666464484
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1666464484
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_61
timestamp 1666464484
transform 1 0 6716 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_72
timestamp 1666464484
transform 1 0 7728 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_79
timestamp 1666464484
transform 1 0 8372 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1666464484
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_112
timestamp 1666464484
transform 1 0 11408 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_124
timestamp 1666464484
transform 1 0 12512 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1666464484
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_146
timestamp 1666464484
transform 1 0 14536 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_150
timestamp 1666464484
transform 1 0 14904 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_167
timestamp 1666464484
transform 1 0 16468 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_179
timestamp 1666464484
transform 1 0 17572 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_191
timestamp 1666464484
transform 1 0 18676 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666464484
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666464484
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666464484
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666464484
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666464484
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666464484
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666464484
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666464484
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666464484
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_398
timestamp 1666464484
transform 1 0 37720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_410
timestamp 1666464484
transform 1 0 38824 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1666464484
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_429
timestamp 1666464484
transform 1 0 40572 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_440
timestamp 1666464484
transform 1 0 41584 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_452
timestamp 1666464484
transform 1 0 42688 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_464
timestamp 1666464484
transform 1 0 43792 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1666464484
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_47
timestamp 1666464484
transform 1 0 5428 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1666464484
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_61
timestamp 1666464484
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_67
timestamp 1666464484
transform 1 0 7268 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_75
timestamp 1666464484
transform 1 0 8004 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_79
timestamp 1666464484
transform 1 0 8372 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_103
timestamp 1666464484
transform 1 0 10580 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_109
timestamp 1666464484
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_132
timestamp 1666464484
transform 1 0 13248 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_156
timestamp 1666464484
transform 1 0 15456 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 1666464484
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_243
timestamp 1666464484
transform 1 0 23460 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_252
timestamp 1666464484
transform 1 0 24288 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_260
timestamp 1666464484
transform 1 0 25024 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1666464484
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_291
timestamp 1666464484
transform 1 0 27876 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_301
timestamp 1666464484
transform 1 0 28796 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_319
timestamp 1666464484
transform 1 0 30452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_331
timestamp 1666464484
transform 1 0 31556 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666464484
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_390
timestamp 1666464484
transform 1 0 36984 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_411
timestamp 1666464484
transform 1 0 38916 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_423
timestamp 1666464484
transform 1 0 40020 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_443
timestamp 1666464484
transform 1 0 41860 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1666464484
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1666464484
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1666464484
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_61
timestamp 1666464484
transform 1 0 6716 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_73
timestamp 1666464484
transform 1 0 7820 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_82
timestamp 1666464484
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_103
timestamp 1666464484
transform 1 0 10580 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_115
timestamp 1666464484
transform 1 0 11684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_132
timestamp 1666464484
transform 1 0 13248 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_146
timestamp 1666464484
transform 1 0 14536 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_166
timestamp 1666464484
transform 1 0 16376 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_176
timestamp 1666464484
transform 1 0 17296 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_188
timestamp 1666464484
transform 1 0 18400 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_225
timestamp 1666464484
transform 1 0 21804 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_229
timestamp 1666464484
transform 1 0 22172 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1666464484
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_258
timestamp 1666464484
transform 1 0 24840 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_264
timestamp 1666464484
transform 1 0 25392 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_270
timestamp 1666464484
transform 1 0 25944 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_279
timestamp 1666464484
transform 1 0 26772 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1666464484
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_328
timestamp 1666464484
transform 1 0 31280 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_340
timestamp 1666464484
transform 1 0 32384 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_355
timestamp 1666464484
transform 1 0 33764 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_377
timestamp 1666464484
transform 1 0 35788 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_381
timestamp 1666464484
transform 1 0 36156 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_385
timestamp 1666464484
transform 1 0 36524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_405
timestamp 1666464484
transform 1 0 38364 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_415
timestamp 1666464484
transform 1 0 39284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_425
timestamp 1666464484
transform 1 0 40204 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_442
timestamp 1666464484
transform 1 0 41768 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_452
timestamp 1666464484
transform 1 0 42688 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_464
timestamp 1666464484
transform 1 0 43792 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_47
timestamp 1666464484
transform 1 0 5428 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_103
timestamp 1666464484
transform 1 0 10580 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1666464484
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_119
timestamp 1666464484
transform 1 0 12052 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_136
timestamp 1666464484
transform 1 0 13616 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_143
timestamp 1666464484
transform 1 0 14260 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 1666464484
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1666464484
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_230
timestamp 1666464484
transform 1 0 22264 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_234
timestamp 1666464484
transform 1 0 22632 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_241
timestamp 1666464484
transform 1 0 23276 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_261
timestamp 1666464484
transform 1 0 25116 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_271
timestamp 1666464484
transform 1 0 26036 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666464484
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_303
timestamp 1666464484
transform 1 0 28980 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_318
timestamp 1666464484
transform 1 0 30360 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_330
timestamp 1666464484
transform 1 0 31464 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_365
timestamp 1666464484
transform 1 0 34684 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_372
timestamp 1666464484
transform 1 0 35328 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_384
timestamp 1666464484
transform 1 0 36432 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_411
timestamp 1666464484
transform 1 0 38916 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_419
timestamp 1666464484
transform 1 0 39652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_425
timestamp 1666464484
transform 1 0 40204 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_445
timestamp 1666464484
transform 1 0 42044 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_478
timestamp 1666464484
transform 1 0 45080 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_490
timestamp 1666464484
transform 1 0 46184 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1666464484
transform 1 0 47288 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1666464484
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1666464484
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_72
timestamp 1666464484
transform 1 0 7728 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_92
timestamp 1666464484
transform 1 0 9568 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_104
timestamp 1666464484
transform 1 0 10672 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_108
timestamp 1666464484
transform 1 0 11040 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_125
timestamp 1666464484
transform 1 0 12604 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_135
timestamp 1666464484
transform 1 0 13524 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_149
timestamp 1666464484
transform 1 0 14812 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_166
timestamp 1666464484
transform 1 0 16376 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_173
timestamp 1666464484
transform 1 0 17020 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_185
timestamp 1666464484
transform 1 0 18124 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_193
timestamp 1666464484
transform 1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_209
timestamp 1666464484
transform 1 0 20332 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_229
timestamp 1666464484
transform 1 0 22172 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_241
timestamp 1666464484
transform 1 0 23276 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1666464484
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_271
timestamp 1666464484
transform 1 0 26036 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_279
timestamp 1666464484
transform 1 0 26772 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_286
timestamp 1666464484
transform 1 0 27416 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_298
timestamp 1666464484
transform 1 0 28520 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_306
timestamp 1666464484
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1666464484
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_345
timestamp 1666464484
transform 1 0 32844 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_362
timestamp 1666464484
transform 1 0 34408 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_375
timestamp 1666464484
transform 1 0 35604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1666464484
transform 1 0 36708 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_407
timestamp 1666464484
transform 1 0 38548 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_411
timestamp 1666464484
transform 1 0 38916 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_418
timestamp 1666464484
transform 1 0 39560 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_443
timestamp 1666464484
transform 1 0 41860 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_455
timestamp 1666464484
transform 1 0 42964 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_474
timestamp 1666464484
transform 1 0 44712 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_47
timestamp 1666464484
transform 1 0 5428 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1666464484
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_67
timestamp 1666464484
transform 1 0 7268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_79
timestamp 1666464484
transform 1 0 8372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_88
timestamp 1666464484
transform 1 0 9200 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_99
timestamp 1666464484
transform 1 0 10212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_122
timestamp 1666464484
transform 1 0 12328 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_134
timestamp 1666464484
transform 1 0 13432 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_146
timestamp 1666464484
transform 1 0 14536 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_157
timestamp 1666464484
transform 1 0 15548 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_165
timestamp 1666464484
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1666464484
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_243
timestamp 1666464484
transform 1 0 23460 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_247
timestamp 1666464484
transform 1 0 23828 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_264
timestamp 1666464484
transform 1 0 25392 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1666464484
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_293
timestamp 1666464484
transform 1 0 28060 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_321
timestamp 1666464484
transform 1 0 30636 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_327
timestamp 1666464484
transform 1 0 31188 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_349
timestamp 1666464484
transform 1 0 33212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_369
timestamp 1666464484
transform 1 0 35052 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1666464484
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_415
timestamp 1666464484
transform 1 0 39284 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_427
timestamp 1666464484
transform 1 0 40388 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_433
timestamp 1666464484
transform 1 0 40940 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_445
timestamp 1666464484
transform 1 0 42044 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_457
timestamp 1666464484
transform 1 0 43148 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_463
timestamp 1666464484
transform 1 0 43700 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_474
timestamp 1666464484
transform 1 0 44712 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_481
timestamp 1666464484
transform 1 0 45356 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_493
timestamp 1666464484
transform 1 0 46460 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_501
timestamp 1666464484
transform 1 0 47196 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1666464484
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1666464484
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_58
timestamp 1666464484
transform 1 0 6440 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_69
timestamp 1666464484
transform 1 0 7452 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_79
timestamp 1666464484
transform 1 0 8372 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_103
timestamp 1666464484
transform 1 0 10580 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_115
timestamp 1666464484
transform 1 0 11684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_127
timestamp 1666464484
transform 1 0 12788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666464484
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1666464484
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1666464484
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666464484
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_258
timestamp 1666464484
transform 1 0 24840 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_270
timestamp 1666464484
transform 1 0 25944 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_282
timestamp 1666464484
transform 1 0 27048 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_294
timestamp 1666464484
transform 1 0 28152 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1666464484
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1666464484
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1666464484
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_345
timestamp 1666464484
transform 1 0 32844 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_353
timestamp 1666464484
transform 1 0 33580 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1666464484
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666464484
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_370
timestamp 1666464484
transform 1 0 35144 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_382
timestamp 1666464484
transform 1 0 36248 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_394
timestamp 1666464484
transform 1 0 37352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_398
timestamp 1666464484
transform 1 0 37720 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_404
timestamp 1666464484
transform 1 0 38272 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_416
timestamp 1666464484
transform 1 0 39376 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_465
timestamp 1666464484
transform 1 0 43884 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_472
timestamp 1666464484
transform 1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_47
timestamp 1666464484
transform 1 0 5428 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1666464484
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_66
timestamp 1666464484
transform 1 0 7176 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_78
timestamp 1666464484
transform 1 0 8280 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_82
timestamp 1666464484
transform 1 0 8648 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_103
timestamp 1666464484
transform 1 0 10580 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1666464484
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1666464484
transform 1 0 12236 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666464484
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1666464484
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1666464484
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1666464484
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666464484
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1666464484
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1666464484
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_411
timestamp 1666464484
transform 1 0 38916 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_423
timestamp 1666464484
transform 1 0 40020 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_431
timestamp 1666464484
transform 1 0 40756 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_438
timestamp 1666464484
transform 1 0 41400 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_446
timestamp 1666464484
transform 1 0 42136 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_455
timestamp 1666464484
transform 1 0 42964 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_459
timestamp 1666464484
transform 1 0 43332 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_479
timestamp 1666464484
transform 1 0 45172 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_491
timestamp 1666464484
transform 1 0 46276 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1666464484
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1666464484
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_61
timestamp 1666464484
transform 1 0 6716 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_73
timestamp 1666464484
transform 1 0 7820 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_81
timestamp 1666464484
transform 1 0 8556 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_91
timestamp 1666464484
transform 1 0 9476 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_111
timestamp 1666464484
transform 1 0 11316 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_135
timestamp 1666464484
transform 1 0 13524 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666464484
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1666464484
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1666464484
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_271
timestamp 1666464484
transform 1 0 26036 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_283
timestamp 1666464484
transform 1 0 27140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_295
timestamp 1666464484
transform 1 0 28244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1666464484
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1666464484
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1666464484
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1666464484
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_377
timestamp 1666464484
transform 1 0 35788 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_382
timestamp 1666464484
transform 1 0 36248 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_402
timestamp 1666464484
transform 1 0 38088 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_412
timestamp 1666464484
transform 1 0 39008 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_439
timestamp 1666464484
transform 1 0 41492 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_449
timestamp 1666464484
transform 1 0 42412 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_474
timestamp 1666464484
transform 1 0 44712 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_484
timestamp 1666464484
transform 1 0 45632 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_496
timestamp 1666464484
transform 1 0 46736 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_508
timestamp 1666464484
transform 1 0 47840 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_520
timestamp 1666464484
transform 1 0 48944 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_47
timestamp 1666464484
transform 1 0 5428 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1666464484
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_66
timestamp 1666464484
transform 1 0 7176 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_75
timestamp 1666464484
transform 1 0 8004 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_90
timestamp 1666464484
transform 1 0 9384 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1666464484
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1666464484
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_256
timestamp 1666464484
transform 1 0 24656 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_268
timestamp 1666464484
transform 1 0 25760 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1666464484
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1666464484
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1666464484
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1666464484
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_373
timestamp 1666464484
transform 1 0 35420 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_379
timestamp 1666464484
transform 1 0 35972 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_383
timestamp 1666464484
transform 1 0 36340 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1666464484
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_411
timestamp 1666464484
transform 1 0 38916 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_415
timestamp 1666464484
transform 1 0 39284 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_419
timestamp 1666464484
transform 1 0 39652 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_439
timestamp 1666464484
transform 1 0 41492 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_446
timestamp 1666464484
transform 1 0 42136 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_483
timestamp 1666464484
transform 1 0 45540 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_495
timestamp 1666464484
transform 1 0 46644 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1666464484
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1666464484
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_45
timestamp 1666464484
transform 1 0 5244 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_62
timestamp 1666464484
transform 1 0 6808 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_66
timestamp 1666464484
transform 1 0 7176 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_74
timestamp 1666464484
transform 1 0 7912 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_81
timestamp 1666464484
transform 1 0 8556 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_98
timestamp 1666464484
transform 1 0 10120 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_106
timestamp 1666464484
transform 1 0 10856 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_118
timestamp 1666464484
transform 1 0 11960 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_130
timestamp 1666464484
transform 1 0 13064 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1666464484
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1666464484
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1666464484
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1666464484
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1666464484
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1666464484
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666464484
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1666464484
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1666464484
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_405
timestamp 1666464484
transform 1 0 38364 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1666464484
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_441
timestamp 1666464484
transform 1 0 41676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_448
timestamp 1666464484
transform 1 0 42320 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_454
timestamp 1666464484
transform 1 0 42872 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_458
timestamp 1666464484
transform 1 0 43240 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_468
timestamp 1666464484
transform 1 0 44160 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_482
timestamp 1666464484
transform 1 0 45448 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1666464484
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_62
timestamp 1666464484
transform 1 0 6808 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_68
timestamp 1666464484
transform 1 0 7360 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_85
timestamp 1666464484
transform 1 0 8924 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_94
timestamp 1666464484
transform 1 0 9752 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_106
timestamp 1666464484
transform 1 0 10856 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1666464484
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_299
timestamp 1666464484
transform 1 0 28612 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_311
timestamp 1666464484
transform 1 0 29716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_323
timestamp 1666464484
transform 1 0 30820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1666464484
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1666464484
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_398
timestamp 1666464484
transform 1 0 37720 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_410
timestamp 1666464484
transform 1 0 38824 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_422
timestamp 1666464484
transform 1 0 39928 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1666464484
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_467
timestamp 1666464484
transform 1 0 44068 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_484
timestamp 1666464484
transform 1 0 45632 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_496
timestamp 1666464484
transform 1 0 46736 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1666464484
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1666464484
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_61
timestamp 1666464484
transform 1 0 6716 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_73
timestamp 1666464484
transform 1 0 7820 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1666464484
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1666464484
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1666464484
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1666464484
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1666464484
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1666464484
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1666464484
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1666464484
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1666464484
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1666464484
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666464484
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_427
timestamp 1666464484
transform 1 0 40388 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_431
timestamp 1666464484
transform 1 0 40756 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_443
timestamp 1666464484
transform 1 0 41860 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_455
timestamp 1666464484
transform 1 0 42964 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_467
timestamp 1666464484
transform 1 0 44068 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_495
timestamp 1666464484
transform 1 0 46644 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_507
timestamp 1666464484
transform 1 0 47748 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_519
timestamp 1666464484
transform 1 0 48852 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1666464484
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1666464484
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1666464484
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1666464484
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1666464484
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1666464484
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1666464484
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1666464484
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1666464484
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1666464484
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1666464484
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1666464484
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1666464484
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1666464484
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1666464484
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1666464484
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1666464484
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1666464484
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1666464484
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1666464484
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1666464484
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1666464484
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1666464484
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1666464484
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1666464484
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1666464484
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1666464484
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1666464484
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1666464484
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1666464484
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1666464484
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1666464484
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1666464484
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1666464484
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1666464484
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1666464484
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1666464484
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1666464484
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1666464484
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1666464484
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1666464484
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1666464484
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1666464484
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1666464484
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1666464484
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1666464484
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1666464484
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1666464484
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1666464484
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1666464484
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1666464484
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1666464484
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1666464484
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1666464484
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1666464484
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1666464484
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1666464484
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1666464484
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1666464484
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1666464484
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1666464484
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1666464484
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1666464484
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1666464484
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1666464484
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1666464484
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1666464484
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1666464484
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1666464484
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1666464484
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1666464484
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1666464484
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1666464484
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1666464484
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1666464484
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1666464484
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1666464484
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1666464484
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1666464484
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1666464484
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1666464484
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1666464484
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1666464484
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1666464484
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1666464484
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1666464484
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1666464484
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1666464484
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1666464484
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1666464484
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1666464484
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1666464484
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1666464484
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1666464484
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1666464484
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1666464484
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1666464484
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1666464484
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1666464484
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1666464484
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1666464484
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1666464484
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1666464484
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1666464484
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1666464484
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1666464484
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1666464484
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1666464484
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1666464484
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1666464484
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1666464484
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1666464484
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1666464484
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1666464484
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1666464484
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1666464484
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1666464484
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1666464484
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1666464484
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1666464484
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1666464484
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1666464484
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1666464484
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1666464484
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1666464484
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1666464484
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1666464484
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1666464484
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1666464484
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1666464484
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1666464484
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1666464484
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1666464484
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1666464484
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1666464484
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1666464484
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1666464484
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1666464484
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1666464484
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1666464484
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1666464484
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1666464484
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1666464484
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1666464484
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1666464484
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1666464484
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1666464484
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1666464484
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1666464484
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1666464484
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1666464484
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1666464484
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1666464484
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1666464484
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1666464484
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1666464484
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1666464484
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1666464484
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1666464484
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1666464484
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1666464484
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1666464484
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1666464484
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1666464484
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1666464484
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1666464484
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1666464484
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1666464484
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1666464484
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1666464484
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1666464484
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1666464484
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1666464484
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1666464484
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1666464484
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1666464484
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1666464484
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1666464484
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1666464484
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1666464484
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1666464484
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1666464484
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1666464484
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1666464484
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1666464484
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1666464484
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1666464484
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1666464484
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1666464484
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1666464484
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1666464484
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1666464484
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1666464484
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1666464484
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1666464484
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1666464484
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1666464484
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1666464484
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1666464484
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1666464484
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1666464484
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1666464484
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1666464484
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1666464484
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1666464484
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1666464484
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1666464484
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1666464484
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1666464484
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1666464484
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1666464484
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1666464484
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1666464484
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1666464484
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1666464484
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1666464484
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1666464484
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1666464484
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1666464484
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1666464484
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1666464484
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1666464484
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1666464484
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1666464484
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1666464484
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1666464484
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1666464484
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1666464484
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1666464484
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1666464484
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1666464484
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1666464484
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1666464484
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1666464484
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1666464484
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1666464484
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1666464484
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1666464484
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1666464484
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1666464484
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1666464484
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1666464484
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1666464484
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1666464484
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1666464484
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1666464484
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1666464484
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1666464484
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1666464484
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1666464484
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1666464484
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1666464484
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1666464484
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1666464484
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1666464484
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1666464484
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1666464484
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1666464484
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1666464484
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1666464484
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1666464484
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1666464484
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1666464484
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1666464484
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1666464484
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1666464484
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1666464484
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1666464484
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_41
timestamp 1666464484
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1666464484
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_63
timestamp 1666464484
transform 1 0 6900 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_75
timestamp 1666464484
transform 1 0 8004 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_83
timestamp 1666464484
transform 1 0 8740 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1666464484
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1666464484
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1666464484
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1666464484
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1666464484
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_153
timestamp 1666464484
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1666464484
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1666464484
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1666464484
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1666464484
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1666464484
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1666464484
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_265
timestamp 1666464484
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1666464484
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_293
timestamp 1666464484
transform 1 0 28060 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_301
timestamp 1666464484
transform 1 0 28796 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1666464484
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_309
timestamp 1666464484
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_321
timestamp 1666464484
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1666464484
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1666464484
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1666464484
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_365
timestamp 1666464484
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_377
timestamp 1666464484
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1666464484
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1666464484
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1666464484
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1666464484
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1666464484
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1666464484
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1666464484
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_477
timestamp 1666464484
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_489
timestamp 1666464484
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1666464484
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1666464484
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1666464484
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_539
timestamp 1666464484
transform 1 0 50692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_551
timestamp 1666464484
transform 1 0 51796 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1666464484
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1666464484
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1666464484
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_601
timestamp 1666464484
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_613
timestamp 1666464484
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0501_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45264 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0502_
timestamp 1666464484
transform 1 0 40848 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0503_
timestamp 1666464484
transform 1 0 43976 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0504_
timestamp 1666464484
transform 1 0 46276 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0505_
timestamp 1666464484
transform 1 0 42596 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0506_
timestamp 1666464484
transform 1 0 41860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0507_
timestamp 1666464484
transform 1 0 38640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0508_
timestamp 1666464484
transform 1 0 43332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0509_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0510_
timestamp 1666464484
transform 1 0 38456 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0511_
timestamp 1666464484
transform 1 0 41860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0512_
timestamp 1666464484
transform 1 0 42136 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0513_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44068 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0514_
timestamp 1666464484
transform 1 0 35052 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0515_
timestamp 1666464484
transform 1 0 38180 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0516_
timestamp 1666464484
transform 1 0 38732 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0517_
timestamp 1666464484
transform 1 0 39008 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0518_
timestamp 1666464484
transform -1 0 41400 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44988 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0520_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0521_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34868 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0522_
timestamp 1666464484
transform -1 0 33764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0523_
timestamp 1666464484
transform 1 0 31740 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0524_
timestamp 1666464484
transform 1 0 29716 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0525_
timestamp 1666464484
transform 1 0 33028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0526_
timestamp 1666464484
transform -1 0 35788 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0527_
timestamp 1666464484
transform 1 0 30728 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0528_
timestamp 1666464484
transform 1 0 33212 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0530_
timestamp 1666464484
transform 1 0 39100 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1666464484
transform -1 0 40388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0532_
timestamp 1666464484
transform 1 0 19872 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0533_
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0534_
timestamp 1666464484
transform 1 0 25024 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0535_
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0536_
timestamp 1666464484
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0537_
timestamp 1666464484
transform 1 0 25576 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0538_
timestamp 1666464484
transform -1 0 24656 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _0539_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0540_
timestamp 1666464484
transform -1 0 12880 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0541_
timestamp 1666464484
transform 1 0 2852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0542_
timestamp 1666464484
transform 1 0 34868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0543_
timestamp 1666464484
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0544_
timestamp 1666464484
transform -1 0 36156 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0545_
timestamp 1666464484
transform 1 0 32752 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0546_
timestamp 1666464484
transform 1 0 32384 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0547_
timestamp 1666464484
transform 1 0 29716 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0548_
timestamp 1666464484
transform 1 0 32936 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1666464484
transform -1 0 38272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0550_
timestamp 1666464484
transform 1 0 41584 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1666464484
transform -1 0 43516 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0553_
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0554_
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0555_
timestamp 1666464484
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0556_
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0557_
timestamp 1666464484
transform 1 0 18768 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0558_
timestamp 1666464484
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0559_
timestamp 1666464484
transform 1 0 18768 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1666464484
transform -1 0 18952 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0561_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21068 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1666464484
transform 1 0 20148 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0563_
timestamp 1666464484
transform 1 0 7176 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0564_
timestamp 1666464484
transform 1 0 6808 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0565_
timestamp 1666464484
transform 1 0 16744 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0566_
timestamp 1666464484
transform 1 0 12972 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0567_
timestamp 1666464484
transform 1 0 13064 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0568_
timestamp 1666464484
transform 1 0 10948 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0569_
timestamp 1666464484
transform -1 0 13248 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0570_
timestamp 1666464484
transform -1 0 7728 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0571_
timestamp 1666464484
transform -1 0 8372 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0573_
timestamp 1666464484
transform 1 0 25484 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0574_
timestamp 1666464484
transform 1 0 22724 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0575_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0576_
timestamp 1666464484
transform 1 0 26588 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0577_
timestamp 1666464484
transform 1 0 24564 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1666464484
transform 1 0 23092 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0580_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27048 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1666464484
transform 1 0 43148 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0582_
timestamp 1666464484
transform 1 0 40848 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0583_
timestamp 1666464484
transform 1 0 42596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0584_
timestamp 1666464484
transform 1 0 37444 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0585_
timestamp 1666464484
transform 1 0 40204 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0586_
timestamp 1666464484
transform 1 0 37444 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0587_
timestamp 1666464484
transform 1 0 38456 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0588_
timestamp 1666464484
transform 1 0 43884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0589_
timestamp 1666464484
transform 1 0 4048 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0590_
timestamp 1666464484
transform -1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0591_
timestamp 1666464484
transform -1 0 7452 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0592_
timestamp 1666464484
transform 1 0 3956 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0593_
timestamp 1666464484
transform 1 0 3956 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0594_
timestamp 1666464484
transform 1 0 4600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0595_
timestamp 1666464484
transform -1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0596_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9384 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0597_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6256 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0598_
timestamp 1666464484
transform 1 0 6808 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0599_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9568 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0600_
timestamp 1666464484
transform 1 0 10948 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0601_
timestamp 1666464484
transform -1 0 10120 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0602_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10856 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0603_
timestamp 1666464484
transform -1 0 9476 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0604_
timestamp 1666464484
transform -1 0 9752 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0605_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7268 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1666464484
transform 1 0 8280 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1666464484
transform -1 0 6072 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1666464484
transform -1 0 8004 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0609_
timestamp 1666464484
transform 1 0 6532 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1666464484
transform 1 0 6532 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1666464484
transform 1 0 5612 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0612_
timestamp 1666464484
transform -1 0 7176 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1666464484
transform 1 0 5704 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0614_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1666464484
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0616_
timestamp 1666464484
transform -1 0 22264 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0618_
timestamp 1666464484
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0619_
timestamp 1666464484
transform -1 0 21436 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0620_
timestamp 1666464484
transform -1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0621_
timestamp 1666464484
transform -1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0622_
timestamp 1666464484
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0623_
timestamp 1666464484
transform -1 0 22356 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0624_
timestamp 1666464484
transform 1 0 20884 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1666464484
transform 1 0 22632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0626_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0627_
timestamp 1666464484
transform -1 0 20976 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0628_
timestamp 1666464484
transform 1 0 19780 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1666464484
transform 1 0 21252 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0630_
timestamp 1666464484
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0632_
timestamp 1666464484
transform -1 0 39744 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0633_
timestamp 1666464484
transform 1 0 39284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0634_
timestamp 1666464484
transform -1 0 40756 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1666464484
transform 1 0 40204 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0636_
timestamp 1666464484
transform 1 0 41032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1666464484
transform 1 0 39928 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1666464484
transform 1 0 40020 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1666464484
transform 1 0 40848 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0640_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 40204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0641_
timestamp 1666464484
transform -1 0 40664 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1666464484
transform 1 0 39192 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0643_
timestamp 1666464484
transform 1 0 41124 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0644_
timestamp 1666464484
transform -1 0 40756 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1666464484
transform -1 0 40296 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0646_
timestamp 1666464484
transform 1 0 40756 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0647_
timestamp 1666464484
transform 1 0 41860 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1666464484
transform 1 0 42688 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0649_
timestamp 1666464484
transform -1 0 13800 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0651_
timestamp 1666464484
transform -1 0 15732 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1666464484
transform 1 0 14260 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0653_
timestamp 1666464484
transform 1 0 14352 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1666464484
transform -1 0 15456 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0655_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0656_
timestamp 1666464484
transform 1 0 13248 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0657_
timestamp 1666464484
transform -1 0 13616 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1666464484
transform -1 0 13064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1666464484
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0660_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14904 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0661_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1666464484
transform -1 0 36984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1666464484
transform 1 0 36616 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0664_
timestamp 1666464484
transform 1 0 37996 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 1666464484
transform 1 0 37812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0666_
timestamp 1666464484
transform 1 0 37352 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1666464484
transform 1 0 37720 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0668_
timestamp 1666464484
transform 1 0 38180 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp 1666464484
transform 1 0 38824 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1666464484
transform -1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0671_
timestamp 1666464484
transform -1 0 44160 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1666464484
transform -1 0 43240 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0673_
timestamp 1666464484
transform 1 0 43056 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1666464484
transform 1 0 44068 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0675_
timestamp 1666464484
transform 1 0 45172 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1666464484
transform 1 0 45172 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0677_
timestamp 1666464484
transform -1 0 43424 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0678_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0679_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0680_
timestamp 1666464484
transform -1 0 8740 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_4  _0681_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4692 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0682_
timestamp 1666464484
transform -1 0 12236 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1666464484
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1666464484
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0685_
timestamp 1666464484
transform -1 0 13064 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0686_
timestamp 1666464484
transform 1 0 11684 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1666464484
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0688_
timestamp 1666464484
transform 1 0 10856 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1666464484
transform 1 0 10764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0690_
timestamp 1666464484
transform 1 0 11684 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1666464484
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0692_
timestamp 1666464484
transform 1 0 11684 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0693_
timestamp 1666464484
transform 1 0 10488 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1666464484
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1666464484
transform 1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1666464484
transform -1 0 10304 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0697_
timestamp 1666464484
transform -1 0 9568 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0698_
timestamp 1666464484
transform -1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 1666464484
transform -1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0700_
timestamp 1666464484
transform 1 0 8924 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0701_
timestamp 1666464484
transform -1 0 8096 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1666464484
transform 1 0 7544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0703_
timestamp 1666464484
transform 1 0 7176 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0704_
timestamp 1666464484
transform -1 0 8464 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0705_
timestamp 1666464484
transform -1 0 9752 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1666464484
transform -1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0707_
timestamp 1666464484
transform 1 0 9108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0708_
timestamp 1666464484
transform 1 0 7728 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1666464484
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0710_
timestamp 1666464484
transform 1 0 4600 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0711_
timestamp 1666464484
transform 1 0 4232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp 1666464484
transform -1 0 5796 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1666464484
transform -1 0 5796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 1666464484
transform -1 0 3496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0715_
timestamp 1666464484
transform -1 0 44160 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0716_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 43884 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1666464484
transform -1 0 44712 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0718_
timestamp 1666464484
transform 1 0 43792 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _0719_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 44528 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _0720_
timestamp 1666464484
transform 1 0 43056 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0721_
timestamp 1666464484
transform 1 0 43240 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0722_
timestamp 1666464484
transform 1 0 44436 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1666464484
transform 1 0 45172 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0724_
timestamp 1666464484
transform 1 0 45172 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0725_
timestamp 1666464484
transform -1 0 46276 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0726_
timestamp 1666464484
transform 1 0 41768 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0727_
timestamp 1666464484
transform 1 0 42596 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0728_
timestamp 1666464484
transform -1 0 42688 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1666464484
transform -1 0 41400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0730_
timestamp 1666464484
transform 1 0 43424 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0731_
timestamp 1666464484
transform -1 0 43332 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0732_
timestamp 1666464484
transform -1 0 42136 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1666464484
transform 1 0 45172 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1666464484
transform 1 0 44896 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0735_
timestamp 1666464484
transform 1 0 45264 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0736_
timestamp 1666464484
transform -1 0 46368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1666464484
transform 1 0 42872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0738_
timestamp 1666464484
transform 1 0 44344 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0739_
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0740_
timestamp 1666464484
transform -1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0741_
timestamp 1666464484
transform -1 0 43976 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0742_
timestamp 1666464484
transform 1 0 42780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0743_
timestamp 1666464484
transform -1 0 43148 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0744_
timestamp 1666464484
transform -1 0 42136 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0745_
timestamp 1666464484
transform -1 0 43424 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0746_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 43424 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0747_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 42136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0748_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43792 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0749_
timestamp 1666464484
transform -1 0 30728 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0750_
timestamp 1666464484
transform -1 0 27784 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _0751_
timestamp 1666464484
transform -1 0 28612 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _0752_
timestamp 1666464484
transform 1 0 29900 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1666464484
transform 1 0 30084 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1666464484
transform 1 0 30544 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1666464484
transform -1 0 31556 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0756_
timestamp 1666464484
transform 1 0 30728 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1666464484
transform -1 0 31924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0758_
timestamp 1666464484
transform 1 0 29348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0759_
timestamp 1666464484
transform 1 0 29992 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0760_
timestamp 1666464484
transform 1 0 29808 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 1666464484
transform 1 0 31556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0762_
timestamp 1666464484
transform 1 0 31556 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0763_
timestamp 1666464484
transform -1 0 29256 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1666464484
transform -1 0 28244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0765_
timestamp 1666464484
transform 1 0 26404 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0766_
timestamp 1666464484
transform -1 0 28428 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0767_
timestamp 1666464484
transform -1 0 27600 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 1666464484
transform -1 0 27324 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0769_
timestamp 1666464484
transform -1 0 29072 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0770_
timestamp 1666464484
transform 1 0 27692 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0771_
timestamp 1666464484
transform -1 0 27324 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1666464484
transform -1 0 26312 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0773_
timestamp 1666464484
transform 1 0 26312 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0774_
timestamp 1666464484
transform 1 0 27140 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0775_
timestamp 1666464484
transform 1 0 28244 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1666464484
transform -1 0 9200 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0777_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11316 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0778_
timestamp 1666464484
transform 1 0 9752 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0779_
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0780_
timestamp 1666464484
transform -1 0 6808 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0781_
timestamp 1666464484
transform 1 0 4968 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0782_
timestamp 1666464484
transform 1 0 5612 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0783__235 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0783_
timestamp 1666464484
transform 1 0 6716 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0784__234
timestamp 1666464484
transform -1 0 6072 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0784_
timestamp 1666464484
transform 1 0 5520 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0785__233
timestamp 1666464484
transform -1 0 14260 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0785_
timestamp 1666464484
transform -1 0 13616 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0786_
timestamp 1666464484
transform 1 0 12052 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0786__232
timestamp 1666464484
transform -1 0 12604 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0787__231
timestamp 1666464484
transform -1 0 12328 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0787_
timestamp 1666464484
transform 1 0 11776 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0788_
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0788__230
timestamp 1666464484
transform 1 0 10948 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0789__229
timestamp 1666464484
transform 1 0 14260 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0789_
timestamp 1666464484
transform 1 0 14904 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0790__228
timestamp 1666464484
transform -1 0 17020 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0790_
timestamp 1666464484
transform 1 0 14904 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0791_
timestamp 1666464484
transform 1 0 14904 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0791__227
timestamp 1666464484
transform 1 0 14260 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0792__226
timestamp 1666464484
transform -1 0 15548 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0792_
timestamp 1666464484
transform 1 0 14996 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0793__225
timestamp 1666464484
transform 1 0 11868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0793_
timestamp 1666464484
transform 1 0 12512 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0794__224
timestamp 1666464484
transform -1 0 11960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0794_
timestamp 1666464484
transform 1 0 11224 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0795_
timestamp 1666464484
transform 1 0 11592 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0795__223
timestamp 1666464484
transform -1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0796__222
timestamp 1666464484
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0796_
timestamp 1666464484
transform 1 0 9752 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0797__221
timestamp 1666464484
transform -1 0 9568 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0797_
timestamp 1666464484
transform 1 0 9108 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0798_
timestamp 1666464484
transform 1 0 9108 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0798__220
timestamp 1666464484
transform 1 0 8372 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0799__219
timestamp 1666464484
transform 1 0 8096 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0799_
timestamp 1666464484
transform 1 0 9108 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0800__218
timestamp 1666464484
transform -1 0 5796 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0800_
timestamp 1666464484
transform 1 0 5244 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0801__217
timestamp 1666464484
transform -1 0 5888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0801_
timestamp 1666464484
transform 1 0 5244 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0802_
timestamp 1666464484
transform 1 0 5244 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0802__216
timestamp 1666464484
transform -1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0803__215
timestamp 1666464484
transform 1 0 8096 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0803_
timestamp 1666464484
transform -1 0 8556 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0804_
timestamp 1666464484
transform 1 0 44160 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0805_
timestamp 1666464484
transform 1 0 20056 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0806_
timestamp 1666464484
transform 1 0 19688 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0807_
timestamp 1666464484
transform 1 0 21528 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0808_
timestamp 1666464484
transform 1 0 21988 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0809_
timestamp 1666464484
transform -1 0 20884 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0810_
timestamp 1666464484
transform -1 0 20148 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0811__214
timestamp 1666464484
transform -1 0 12972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0811_
timestamp 1666464484
transform 1 0 12328 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0812__213
timestamp 1666464484
transform -1 0 13800 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0812_
timestamp 1666464484
transform 1 0 13340 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0813__212
timestamp 1666464484
transform -1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0813_
timestamp 1666464484
transform 1 0 13340 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0814_
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0814__211
timestamp 1666464484
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0815__210
timestamp 1666464484
transform -1 0 17664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0815_
timestamp 1666464484
transform 1 0 17020 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0816_
timestamp 1666464484
transform 1 0 16744 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0816__209
timestamp 1666464484
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0817_
timestamp 1666464484
transform 1 0 16928 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0817__208
timestamp 1666464484
transform 1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0818__207
timestamp 1666464484
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0818_
timestamp 1666464484
transform 1 0 17480 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0819__206
timestamp 1666464484
transform -1 0 21252 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0819_
timestamp 1666464484
transform 1 0 20240 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0820__205
timestamp 1666464484
transform -1 0 22264 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0820_
timestamp 1666464484
transform 1 0 20148 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0821__204
timestamp 1666464484
transform -1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0821_
timestamp 1666464484
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0822__203
timestamp 1666464484
transform 1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0822_
timestamp 1666464484
transform 1 0 20056 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0823__202
timestamp 1666464484
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0823_
timestamp 1666464484
transform 1 0 16836 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0824__201
timestamp 1666464484
transform -1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0824_
timestamp 1666464484
transform 1 0 16560 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0825__200
timestamp 1666464484
transform -1 0 17204 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0825_
timestamp 1666464484
transform 1 0 16652 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0826__199
timestamp 1666464484
transform -1 0 17848 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0826_
timestamp 1666464484
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0827_
timestamp 1666464484
transform 1 0 14260 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0827__198
timestamp 1666464484
transform 1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0828__197
timestamp 1666464484
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0828_
timestamp 1666464484
transform 1 0 14536 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0829__196
timestamp 1666464484
transform -1 0 14904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0829_
timestamp 1666464484
transform 1 0 14352 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0830__195
timestamp 1666464484
transform -1 0 17112 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0830_
timestamp 1666464484
transform 1 0 15088 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0831__194
timestamp 1666464484
transform -1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0831_
timestamp 1666464484
transform 1 0 15732 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0832__193
timestamp 1666464484
transform 1 0 15272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0832_
timestamp 1666464484
transform 1 0 15916 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0833_
timestamp 1666464484
transform -1 0 3036 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0834_
timestamp 1666464484
transform 1 0 39744 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0835_
timestamp 1666464484
transform 1 0 40480 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0836_
timestamp 1666464484
transform 1 0 38640 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0837_
timestamp 1666464484
transform 1 0 40020 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0838_
timestamp 1666464484
transform 1 0 40664 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0839__192
timestamp 1666464484
transform -1 0 36708 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0839_
timestamp 1666464484
transform 1 0 36156 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0840__191
timestamp 1666464484
transform 1 0 27232 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0840_
timestamp 1666464484
transform 1 0 27784 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0841__190
timestamp 1666464484
transform -1 0 29072 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0841_
timestamp 1666464484
transform 1 0 27784 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0842_
timestamp 1666464484
transform 1 0 36156 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0842__189
timestamp 1666464484
transform -1 0 38364 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0843__188
timestamp 1666464484
transform -1 0 36800 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0843_
timestamp 1666464484
transform 1 0 36248 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0844__187
timestamp 1666464484
transform -1 0 28428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0844_
timestamp 1666464484
transform 1 0 27876 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0845__186
timestamp 1666464484
transform -1 0 30636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0845_
timestamp 1666464484
transform 1 0 29992 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0846__185
timestamp 1666464484
transform 1 0 32384 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0846_
timestamp 1666464484
transform 1 0 33028 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0847__184
timestamp 1666464484
transform -1 0 35144 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0847_
timestamp 1666464484
transform 1 0 32936 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0848__183
timestamp 1666464484
transform -1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0848_
timestamp 1666464484
transform 1 0 30360 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0849__182
timestamp 1666464484
transform -1 0 33580 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0849_
timestamp 1666464484
transform 1 0 32936 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0850__181
timestamp 1666464484
transform -1 0 31096 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0850_
timestamp 1666464484
transform 1 0 30544 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0851__180
timestamp 1666464484
transform -1 0 32568 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0851_
timestamp 1666464484
transform 1 0 31372 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0852_
timestamp 1666464484
transform 1 0 33580 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0852__179
timestamp 1666464484
transform -1 0 34224 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0853__178
timestamp 1666464484
transform 1 0 34132 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0853_
timestamp 1666464484
transform 1 0 35052 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0854__177
timestamp 1666464484
transform 1 0 34776 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0854_
timestamp 1666464484
transform 1 0 34868 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0855__176
timestamp 1666464484
transform 1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0855_
timestamp 1666464484
transform 1 0 34868 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0856__175
timestamp 1666464484
transform -1 0 36984 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0856_
timestamp 1666464484
transform -1 0 36248 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0857_
timestamp 1666464484
transform 1 0 30360 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0857__174
timestamp 1666464484
transform -1 0 31372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0858__173
timestamp 1666464484
transform -1 0 31556 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0858_
timestamp 1666464484
transform 1 0 30912 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0859__172
timestamp 1666464484
transform 1 0 30268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0859_
timestamp 1666464484
transform 1 0 32292 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0860__171
timestamp 1666464484
transform 1 0 29716 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1666464484
transform 1 0 31096 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0861__170
timestamp 1666464484
transform -1 0 28060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0861_
timestamp 1666464484
transform 1 0 27508 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1666464484
transform 1 0 40480 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1666464484
transform 1 0 12880 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1666464484
transform -1 0 16100 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1666464484
transform -1 0 13616 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1666464484
transform -1 0 13800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0867__169
timestamp 1666464484
transform -1 0 23276 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1666464484
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0868__168
timestamp 1666464484
transform 1 0 23092 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0869__167
timestamp 1666464484
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1666464484
transform 1 0 23736 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0870__166
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0871__165
timestamp 1666464484
transform 1 0 20148 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1666464484
transform 1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0872__164
timestamp 1666464484
transform 1 0 20516 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1666464484
transform 1 0 20700 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0873__163
timestamp 1666464484
transform -1 0 21344 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1666464484
transform 1 0 20700 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0874__162
timestamp 1666464484
transform -1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1666464484
transform 1 0 20792 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0875__161
timestamp 1666464484
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1666464484
transform 1 0 24564 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0876__160
timestamp 1666464484
transform -1 0 23460 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1666464484
transform 1 0 22724 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0877__159
timestamp 1666464484
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1666464484
transform 1 0 24564 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0878__158
timestamp 1666464484
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1666464484
transform -1 0 26036 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0879__157
timestamp 1666464484
transform 1 0 21896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1666464484
transform 1 0 23184 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0880__156
timestamp 1666464484
transform -1 0 25392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0881__155
timestamp 1666464484
transform 1 0 22632 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1666464484
transform 1 0 23276 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0882__154
timestamp 1666464484
transform -1 0 23828 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1666464484
transform 1 0 23276 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0883__153
timestamp 1666464484
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1666464484
transform 1 0 16836 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0884__152
timestamp 1666464484
transform -1 0 17572 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1666464484
transform 1 0 17020 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0885__151
timestamp 1666464484
transform -1 0 18584 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1666464484
transform 1 0 18032 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0886__150
timestamp 1666464484
transform -1 0 17572 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1666464484
transform 1 0 17020 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0887__149
timestamp 1666464484
transform 1 0 16928 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1666464484
transform 1 0 17296 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0888__148
timestamp 1666464484
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1666464484
transform 1 0 17020 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0889__147
timestamp 1666464484
transform -1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1666464484
transform 1 0 17020 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0890__146
timestamp 1666464484
transform -1 0 19688 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1666464484
transform 1 0 17572 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1666464484
transform 1 0 45172 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1666464484
transform 1 0 36156 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1666464484
transform 1 0 37444 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1666464484
transform -1 0 40756 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0895__145
timestamp 1666464484
transform -1 0 34224 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1666464484
transform 1 0 32936 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1666464484
transform 1 0 33396 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0896__144
timestamp 1666464484
transform 1 0 32752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0897__143
timestamp 1666464484
transform -1 0 33120 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1666464484
transform 1 0 32568 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1666464484
transform 1 0 32292 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0898__142
timestamp 1666464484
transform 1 0 32292 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1666464484
transform 1 0 34868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0899__141
timestamp 1666464484
transform 1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0900__140
timestamp 1666464484
transform 1 0 31004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1666464484
transform 1 0 32292 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1666464484
transform 1 0 31648 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0901__139
timestamp 1666464484
transform -1 0 32568 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1666464484
transform 1 0 33396 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0902__138
timestamp 1666464484
transform -1 0 34408 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0903__137
timestamp 1666464484
transform -1 0 36984 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1666464484
transform -1 0 36064 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0904__136
timestamp 1666464484
transform -1 0 33212 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1666464484
transform 1 0 30360 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0905__135
timestamp 1666464484
transform 1 0 27140 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1666464484
transform 1 0 27968 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0906__134
timestamp 1666464484
transform -1 0 28520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1666464484
transform 1 0 27784 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0907__133
timestamp 1666464484
transform -1 0 30728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0908__132
timestamp 1666464484
transform 1 0 27324 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1666464484
transform 1 0 27968 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0909__131
timestamp 1666464484
transform 1 0 28244 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1666464484
transform 1 0 28888 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0910__130
timestamp 1666464484
transform 1 0 26404 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1666464484
transform 1 0 27784 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0911__129
timestamp 1666464484
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1666464484
transform 1 0 27784 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1666464484
transform 1 0 29900 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0912__128
timestamp 1666464484
transform 1 0 29808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0913__127
timestamp 1666464484
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1666464484
transform 1 0 29716 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0914__126
timestamp 1666464484
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1666464484
transform 1 0 32292 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0915__125
timestamp 1666464484
transform 1 0 31924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1666464484
transform 1 0 32292 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1666464484
transform 1 0 30084 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0916__124
timestamp 1666464484
transform 1 0 29624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0917__123
timestamp 1666464484
transform -1 0 30912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1666464484
transform 1 0 30268 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0918__122
timestamp 1666464484
transform 1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1666464484
transform 1 0 29900 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0919__121
timestamp 1666464484
transform -1 0 33856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1666464484
transform 1 0 45172 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1666464484
transform 1 0 43240 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1666464484
transform -1 0 45172 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0923__120
timestamp 1666464484
transform 1 0 35972 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1666464484
transform 1 0 36616 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0924__119
timestamp 1666464484
transform 1 0 36708 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1666464484
transform 1 0 37444 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0925__118
timestamp 1666464484
transform 1 0 36064 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0926__117
timestamp 1666464484
transform 1 0 37444 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1666464484
transform 1 0 37444 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0927__116
timestamp 1666464484
transform 1 0 39376 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1666464484
transform 1 0 40020 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0928__115
timestamp 1666464484
transform -1 0 42136 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1666464484
transform 1 0 40020 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0929__114
timestamp 1666464484
transform -1 0 40756 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1666464484
transform 1 0 40112 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0930__113
timestamp 1666464484
transform -1 0 42320 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1666464484
transform 1 0 40204 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1666464484
transform 1 0 40296 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0931__112
timestamp 1666464484
transform -1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0932__111
timestamp 1666464484
transform 1 0 39928 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1666464484
transform 1 0 40388 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0933__110
timestamp 1666464484
transform -1 0 40940 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1666464484
transform 1 0 40388 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0934__109
timestamp 1666464484
transform -1 0 41584 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1666464484
transform 1 0 37444 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0935__108
timestamp 1666464484
transform 1 0 36708 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0936__107
timestamp 1666464484
transform 1 0 36248 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1666464484
transform 1 0 36892 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0937__106
timestamp 1666464484
transform -1 0 37720 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1666464484
transform 1 0 37076 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1666464484
transform 1 0 37444 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0938__105
timestamp 1666464484
transform 1 0 37444 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1666464484
transform 1 0 36340 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0939__104
timestamp 1666464484
transform -1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1666464484
transform 1 0 36524 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0940__103
timestamp 1666464484
transform 1 0 35880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0941__102
timestamp 1666464484
transform -1 0 36984 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1666464484
transform -1 0 36984 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1666464484
transform 1 0 37444 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0942__101
timestamp 1666464484
transform 1 0 37444 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1666464484
transform 1 0 33212 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0943__100
timestamp 1666464484
transform -1 0 33764 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0944__99
timestamp 1666464484
transform -1 0 34132 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1666464484
transform 1 0 33580 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0945__98
timestamp 1666464484
transform 1 0 34868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1666464484
transform -1 0 36892 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1666464484
transform 1 0 32936 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0946__97
timestamp 1666464484
transform -1 0 35328 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0947__96
timestamp 1666464484
transform -1 0 45356 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1666464484
transform -1 0 45080 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0948__95
timestamp 1666464484
transform -1 0 43700 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1666464484
transform 1 0 43240 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1666464484
transform -1 0 3036 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1666464484
transform 1 0 42964 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0951__94
timestamp 1666464484
transform -1 0 43976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1666464484
transform 1 0 43240 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1666464484
transform 1 0 43792 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0952__93
timestamp 1666464484
transform -1 0 46092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0953__92
timestamp 1666464484
transform -1 0 38640 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1666464484
transform 1 0 38088 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0954__91
timestamp 1666464484
transform -1 0 39560 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1666464484
transform 1 0 39008 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0955__90
timestamp 1666464484
transform -1 0 40296 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1666464484
transform 1 0 39100 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0956__89
timestamp 1666464484
transform 1 0 38640 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1666464484
transform 1 0 40020 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0957__88
timestamp 1666464484
transform 1 0 41860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1666464484
transform 1 0 42596 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0958__87
timestamp 1666464484
transform -1 0 43056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1666464484
transform 1 0 42504 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0959__86
timestamp 1666464484
transform 1 0 43240 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1666464484
transform 1 0 44436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0960__85
timestamp 1666464484
transform -1 0 42872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1666464484
transform 1 0 42136 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0961__84
timestamp 1666464484
transform 1 0 39284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1666464484
transform 1 0 39284 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0962__83
timestamp 1666464484
transform 1 0 39928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1666464484
transform 1 0 40020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0963__82
timestamp 1666464484
transform -1 0 41400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1666464484
transform 1 0 40020 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0964__81
timestamp 1666464484
transform -1 0 40848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1666464484
transform 1 0 40020 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0965__80
timestamp 1666464484
transform 1 0 36708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1666464484
transform 1 0 36616 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0966__79
timestamp 1666464484
transform -1 0 39560 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1666464484
transform 1 0 37444 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0967__78
timestamp 1666464484
transform 1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1666464484
transform 1 0 37444 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0968__77
timestamp 1666464484
transform -1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1666464484
transform 1 0 37536 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0969__76
timestamp 1666464484
transform -1 0 44712 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1666464484
transform 1 0 44068 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0970__75
timestamp 1666464484
transform -1 0 45448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1666464484
transform 1 0 44436 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0971__74
timestamp 1666464484
transform -1 0 44712 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1666464484
transform 1 0 44160 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0972__73
timestamp 1666464484
transform 1 0 44436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1666464484
transform 1 0 45172 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0973__72
timestamp 1666464484
transform 1 0 40020 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1666464484
transform 1 0 40204 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1666464484
transform 1 0 40664 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0974__71
timestamp 1666464484
transform 1 0 40756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0975__70
timestamp 1666464484
transform -1 0 41216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1666464484
transform 1 0 40664 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0976__69
timestamp 1666464484
transform 1 0 41584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1666464484
transform 1 0 42596 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0977__68
timestamp 1666464484
transform -1 0 45448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1666464484
transform 1 0 43424 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1666464484
transform 1 0 45264 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1666464484
transform 1 0 11316 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1666464484
transform -1 0 13984 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1666464484
transform -1 0 13156 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1666464484
transform 1 0 10488 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1666464484
transform -1 0 10580 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1666464484
transform 1 0 7084 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1666464484
transform 1 0 7176 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1666464484
transform 1 0 7728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1666464484
transform 1 0 3404 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1666464484
transform 1 0 3496 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0989__67
timestamp 1666464484
transform -1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1666464484
transform 1 0 4600 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0990__66
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1666464484
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0991__65
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1666464484
transform 1 0 6532 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0992__64
timestamp 1666464484
transform -1 0 8648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1666464484
transform -1 0 8004 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1666464484
transform 1 0 2116 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0993__63
timestamp 1666464484
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0994__62
timestamp 1666464484
transform -1 0 4232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1666464484
transform 1 0 2024 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0995__61
timestamp 1666464484
transform -1 0 2760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1666464484
transform 1 0 2024 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0996__60
timestamp 1666464484
transform -1 0 4232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1666464484
transform 1 0 2576 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0997__59
timestamp 1666464484
transform 1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1666464484
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0998__58
timestamp 1666464484
transform 1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1666464484
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0999__57
timestamp 1666464484
transform -1 0 3128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1666464484
transform 1 0 2576 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1000__56
timestamp 1666464484
transform 1 0 4784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1666464484
transform -1 0 5888 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1001__55
timestamp 1666464484
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1666464484
transform 1 0 1932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1002__54
timestamp 1666464484
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1666464484
transform 1 0 2668 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1666464484
transform 1 0 1564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1003__53
timestamp 1666464484
transform -1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1004__52
timestamp 1666464484
transform -1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1666464484
transform 1 0 3404 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1005__51
timestamp 1666464484
transform -1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1666464484
transform 1 0 5428 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1666464484
transform 1 0 6532 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1006__50
timestamp 1666464484
transform 1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1666464484
transform 1 0 27140 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1666464484
transform 1 0 42964 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1666464484
transform -1 0 46552 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1666464484
transform 1 0 41584 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1666464484
transform 1 0 42596 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1666464484
transform -1 0 46644 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1666464484
transform -1 0 46644 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1666464484
transform 1 0 42596 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1666464484
transform 1 0 42688 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1017__49
timestamp 1666464484
transform -1 0 36524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1666464484
transform 1 0 35512 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1666464484
transform 1 0 37812 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1018__48
timestamp 1666464484
transform 1 0 36340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1019__47
timestamp 1666464484
transform -1 0 40480 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1666464484
transform 1 0 38088 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1020__46
timestamp 1666464484
transform -1 0 38916 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1021__45
timestamp 1666464484
transform -1 0 39008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1666464484
transform 1 0 40020 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1022__44
timestamp 1666464484
transform 1 0 37720 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1023__43
timestamp 1666464484
transform 1 0 34408 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1666464484
transform 1 0 35052 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1024__42
timestamp 1666464484
transform -1 0 36432 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1666464484
transform 1 0 35236 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1025__41
timestamp 1666464484
transform -1 0 35788 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1666464484
transform 1 0 35144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1026__40
timestamp 1666464484
transform -1 0 37260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1666464484
transform 1 0 35328 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1027__39
timestamp 1666464484
transform -1 0 41400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1666464484
transform 1 0 40480 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1028__38
timestamp 1666464484
transform 1 0 40664 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1666464484
transform 1 0 42596 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1029__37
timestamp 1666464484
transform -1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1666464484
transform 1 0 41308 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1030__36
timestamp 1666464484
transform -1 0 42872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1666464484
transform 1 0 42320 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1031__35
timestamp 1666464484
transform 1 0 39284 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1666464484
transform 1 0 40112 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1032__34
timestamp 1666464484
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1666464484
transform 1 0 38272 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1666464484
transform 1 0 40020 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1033__33
timestamp 1666464484
transform 1 0 40020 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1034__32
timestamp 1666464484
transform -1 0 40572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1666464484
transform 1 0 40020 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1035__31
timestamp 1666464484
transform -1 0 37168 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1666464484
transform 1 0 35512 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1666464484
transform 1 0 5244 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1666464484
transform 1 0 29808 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1666464484
transform 1 0 32292 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1666464484
transform -1 0 31188 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1666464484
transform 1 0 29716 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1666464484
transform 1 0 27140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1666464484
transform 1 0 26036 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1666464484
transform 1 0 25208 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1666464484
transform -1 0 28980 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1666464484
transform 1 0 24564 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1045__30
timestamp 1666464484
transform 1 0 24564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1666464484
transform 1 0 24564 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1046__29
timestamp 1666464484
transform 1 0 23828 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1666464484
transform 1 0 24748 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1047__28
timestamp 1666464484
transform -1 0 26404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1048__27
timestamp 1666464484
transform -1 0 27140 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1666464484
transform 1 0 25024 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1666464484
transform 1 0 23460 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1049__26
timestamp 1666464484
transform -1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1050__25
timestamp 1666464484
transform 1 0 22908 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1666464484
transform 1 0 23184 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1051__24
timestamp 1666464484
transform -1 0 23828 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1666464484
transform 1 0 23276 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1666464484
transform 1 0 22632 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1052__23
timestamp 1666464484
transform -1 0 23092 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1666464484
transform 1 0 21252 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1053__22
timestamp 1666464484
transform 1 0 20608 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1666464484
transform 1 0 21988 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1054__21
timestamp 1666464484
transform 1 0 20884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1666464484
transform 1 0 21528 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1055__20
timestamp 1666464484
transform -1 0 22264 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1056__19
timestamp 1666464484
transform -1 0 22264 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1666464484
transform -1 0 21528 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1057__18
timestamp 1666464484
transform 1 0 23828 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1666464484
transform 1 0 24564 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1058__17
timestamp 1666464484
transform 1 0 24380 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1666464484
transform 1 0 24564 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1666464484
transform 1 0 23644 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1059__16
timestamp 1666464484
transform -1 0 24840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1060__15
timestamp 1666464484
transform -1 0 24840 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1666464484
transform 1 0 23920 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1061__14
timestamp 1666464484
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1666464484
transform 1 0 21988 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1666464484
transform 1 0 20700 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1062__13
timestamp 1666464484
transform -1 0 21344 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1063__12
timestamp 1666464484
transform 1 0 21252 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1666464484
transform 1 0 21988 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1064__11
timestamp 1666464484
transform 1 0 21528 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1666464484
transform 1 0 22172 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1666464484
transform 1 0 19964 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1666464484
transform 1 0 9108 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23368 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1666464484
transform -1 0 14812 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1666464484
transform 1 0 31188 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1666464484
transform 1 0 4140 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1666464484
transform -1 0 4416 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1666464484
transform 1 0 13984 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1666464484
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1666464484
transform 1 0 7268 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1666464484
transform 1 0 8740 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1666464484
transform -1 0 15456 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1666464484
transform -1 0 24104 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1666464484
transform 1 0 23920 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1666464484
transform 1 0 29992 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1666464484
transform 1 0 28796 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1666464484
transform 1 0 37444 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1666464484
transform -1 0 44620 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1666464484
transform 1 0 39376 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1666464484
transform 1 0 44252 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1666464484
transform 1 0 37444 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1666464484
transform 1 0 32844 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1666464484
transform 1 0 30084 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1666464484
transform 1 0 36064 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1666464484
transform 1 0 41492 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1666464484
transform 1 0 41400 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1666464484
transform -1 0 42964 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1666464484
transform 1 0 30084 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1666464484
transform 1 0 23644 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1666464484
transform 1 0 18492 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1666464484
transform 1 0 18124 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1666464484
transform 1 0 12512 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1666464484
transform -1 0 6164 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_opt_1_0_clk
timestamp 1666464484
transform -1 0 10580 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_opt_2_0_clk
timestamp 1666464484
transform 1 0 42780 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_opt_3_0_clk
timestamp 1666464484
transform 1 0 41124 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 58052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1666464484
transform 1 0 50324 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 58052 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 6900 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 28796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform 1 0 58052 0 -1 27200
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 44888 800 45008 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 59200 3408 59800 3528 0 FreeSans 480 0 0 0 cout1
port 1 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 cout10
port 2 nsew signal tristate
flabel metal2 s 49606 59200 49662 59800 0 FreeSans 224 90 0 0 cout2
port 3 nsew signal tristate
flabel metal2 s 42522 200 42578 800 0 FreeSans 224 90 0 0 cout3
port 4 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 cout4
port 5 nsew signal tristate
flabel metal3 s 59200 48968 59800 49088 0 FreeSans 480 0 0 0 cout5
port 6 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 cout6
port 7 nsew signal tristate
flabel metal2 s 6458 59200 6514 59800 0 FreeSans 224 90 0 0 cout7
port 8 nsew signal tristate
flabel metal2 s 28354 59200 28410 59800 0 FreeSans 224 90 0 0 cout8
port 9 nsew signal tristate
flabel metal3 s 59200 26528 59800 26648 0 FreeSans 480 0 0 0 cout9
port 10 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 4646 13158 4646 13158 0 _0000_
rlabel metal1 45392 10030 45392 10030 0 _0001_
rlabel metal1 45673 45866 45673 45866 0 _0002_
rlabel metal1 40700 9554 40700 9554 0 _0003_
rlabel metal1 2821 22678 2821 22678 0 _0004_
rlabel metal1 43976 38522 43976 38522 0 _0005_
rlabel via1 20281 10030 20281 10030 0 _0006_
rlabel metal2 5842 45730 5842 45730 0 _0007_
rlabel metal2 27278 43622 27278 43622 0 _0008_
rlabel via1 45581 25942 45581 25942 0 _0009_
rlabel metal1 11040 43418 11040 43418 0 _0010_
rlabel metal1 9568 43962 9568 43962 0 _0011_
rlabel metal2 8326 45254 8326 45254 0 _0012_
rlabel via1 6490 44846 6490 44846 0 _0013_
rlabel metal2 5750 42466 5750 42466 0 _0014_
rlabel via1 5929 41582 5929 41582 0 _0015_
rlabel metal2 20746 17510 20746 17510 0 _0037_
rlabel viali 20005 17578 20005 17578 0 _0038_
rlabel metal1 21620 16762 21620 16762 0 _0039_
rlabel metal1 22489 15062 22489 15062 0 _0040_
rlabel metal1 20945 14314 20945 14314 0 _0041_
rlabel metal1 19646 15062 19646 15062 0 _0042_
rlabel metal2 40250 35496 40250 35496 0 _0065_
rlabel metal1 40848 33082 40848 33082 0 _0066_
rlabel metal2 39238 33286 39238 33286 0 _0067_
rlabel via1 40337 37230 40337 37230 0 _0068_
rlabel metal2 42734 37842 42734 37842 0 _0069_
rlabel metal2 13386 26078 13386 26078 0 _0093_
rlabel metal1 15598 24106 15598 24106 0 _0094_
rlabel metal1 13160 22678 13160 22678 0 _0095_
rlabel metal1 14367 23018 14367 23018 0 _0096_
rlabel metal2 36662 21250 36662 21250 0 _0121_
rlabel metal2 37766 21046 37766 21046 0 _0122_
rlabel metal2 39422 21318 39422 21318 0 _0123_
rlabel metal1 43362 43690 43362 43690 0 _0149_
rlabel metal1 45049 43350 45049 43350 0 _0150_
rlabel metal2 43286 13090 43286 13090 0 _0177_
rlabel metal2 11730 10914 11730 10914 0 _0205_
rlabel metal1 13999 13974 13999 13974 0 _0206_
rlabel metal1 13217 14314 13217 14314 0 _0207_
rlabel via1 10805 12206 10805 12206 0 _0208_
rlabel metal1 9618 15470 9618 15470 0 _0209_
rlabel metal1 7498 14586 7498 14586 0 _0210_
rlabel metal2 7314 12002 7314 12002 0 _0211_
rlabel metal1 8827 11798 8827 11798 0 _0212_
rlabel metal1 3997 13906 3997 13906 0 _0213_
rlabel metal1 3542 14586 3542 14586 0 _0214_
rlabel via1 43281 33558 43281 33558 0 _0233_
rlabel metal2 46230 32198 46230 32198 0 _0234_
rlabel viali 41901 31790 41901 31790 0 _0235_
rlabel metal1 42816 30702 42816 30702 0 _0236_
rlabel via1 46326 28526 46326 28526 0 _0237_
rlabel metal1 45452 29546 45452 29546 0 _0238_
rlabel metal1 42488 28118 42488 28118 0 _0239_
rlabel metal2 41906 26146 41906 26146 0 _0240_
rlabel metal2 43838 25058 43838 25058 0 _0241_
rlabel via1 30125 40494 30125 40494 0 _0261_
rlabel metal1 32230 37910 32230 37910 0 _0262_
rlabel metal1 31249 36074 31249 36074 0 _0263_
rlabel metal1 29936 37230 29936 37230 0 _0264_
rlabel metal2 27278 36550 27278 36550 0 _0265_
rlabel viali 26353 37230 26353 37230 0 _0266_
rlabel metal1 26353 40018 26353 40018 0 _0267_
rlabel metal2 28290 40630 28290 40630 0 _0268_
rlabel metal2 9062 42466 9062 42466 0 _0289_
rlabel metal2 43378 25772 43378 25772 0 _0290_
rlabel metal1 42412 24922 42412 24922 0 _0291_
rlabel metal2 28382 37196 28382 37196 0 _0292_
rlabel metal1 27922 40460 27922 40460 0 _0293_
rlabel metal2 28474 40188 28474 40188 0 _0294_
rlabel metal2 30406 40630 30406 40630 0 _0295_
rlabel metal2 30774 38488 30774 38488 0 _0296_
rlabel metal1 31050 37978 31050 37978 0 _0297_
rlabel metal1 31418 38318 31418 38318 0 _0298_
rlabel metal2 29670 37944 29670 37944 0 _0299_
rlabel metal2 30038 36992 30038 36992 0 _0300_
rlabel metal2 31786 37298 31786 37298 0 _0301_
rlabel metal1 30222 37094 30222 37094 0 _0302_
rlabel metal1 28336 37230 28336 37230 0 _0303_
rlabel metal1 27094 36890 27094 36890 0 _0304_
rlabel metal1 27684 37978 27684 37978 0 _0305_
rlabel metal2 27094 36890 27094 36890 0 _0306_
rlabel metal1 27968 38454 27968 38454 0 _0307_
rlabel metal1 27324 38182 27324 38182 0 _0308_
rlabel metal1 26404 38318 26404 38318 0 _0309_
rlabel metal1 27370 40052 27370 40052 0 _0310_
rlabel metal2 44206 13464 44206 13464 0 _0311_
rlabel metal2 43102 12240 43102 12240 0 _0312_
rlabel metal1 44252 12614 44252 12614 0 _0313_
rlabel metal2 43654 17476 43654 17476 0 _0314_
rlabel metal2 43378 17952 43378 17952 0 _0315_
rlabel metal1 42918 15674 42918 15674 0 _0316_
rlabel metal1 43378 17544 43378 17544 0 _0317_
rlabel metal1 43884 17510 43884 17510 0 _0318_
rlabel metal2 40986 43486 40986 43486 0 _0319_
rlabel metal1 41078 43316 41078 43316 0 _0320_
rlabel metal2 42642 41922 42642 41922 0 _0321_
rlabel metal2 39330 41820 39330 41820 0 _0322_
rlabel metal1 37306 41786 37306 41786 0 _0323_
rlabel metal2 38686 39372 38686 39372 0 _0324_
rlabel metal1 39192 40698 39192 40698 0 _0325_
rlabel metal1 40434 41786 40434 41786 0 _0326_
rlabel metal1 44114 44982 44114 44982 0 _0327_
rlabel metal2 45494 44676 45494 44676 0 _0328_
rlabel metal1 35006 24310 35006 24310 0 _0329_
rlabel metal2 33258 25568 33258 25568 0 _0330_
rlabel metal1 32706 24378 32706 24378 0 _0331_
rlabel metal1 32338 25262 32338 25262 0 _0332_
rlabel metal2 33902 23562 33902 23562 0 _0333_
rlabel metal1 33994 19890 33994 19890 0 _0334_
rlabel metal2 33258 20604 33258 20604 0 _0335_
rlabel metal1 33902 20026 33902 20026 0 _0336_
rlabel metal2 38870 21148 38870 21148 0 _0337_
rlabel metal1 39882 20230 39882 20230 0 _0338_
rlabel metal1 19826 25874 19826 25874 0 _0339_
rlabel metal2 19366 24820 19366 24820 0 _0340_
rlabel metal1 24426 25874 24426 25874 0 _0341_
rlabel metal1 24748 25670 24748 25670 0 _0342_
rlabel metal1 24426 25772 24426 25772 0 _0343_
rlabel metal1 25530 23834 25530 23834 0 _0344_
rlabel metal1 18906 25908 18906 25908 0 _0345_
rlabel metal2 15870 24752 15870 24752 0 _0346_
rlabel metal2 12374 23562 12374 23562 0 _0347_
rlabel metal2 37490 34782 37490 34782 0 _0348_
rlabel metal2 38042 34170 38042 34170 0 _0349_
rlabel metal1 34454 32538 34454 32538 0 _0350_
rlabel metal1 33166 33082 33166 33082 0 _0351_
rlabel metal1 33028 30906 33028 30906 0 _0352_
rlabel metal1 32361 32810 32361 32810 0 _0353_
rlabel metal2 38226 33524 38226 33524 0 _0354_
rlabel metal2 41906 37434 41906 37434 0 _0355_
rlabel metal2 42090 38148 42090 38148 0 _0356_
rlabel metal1 19964 16150 19964 16150 0 _0357_
rlabel metal2 17802 15402 17802 15402 0 _0358_
rlabel metal1 18722 14416 18722 14416 0 _0359_
rlabel metal2 22586 20604 22586 20604 0 _0360_
rlabel metal2 19090 20774 19090 20774 0 _0361_
rlabel metal1 19136 18394 19136 18394 0 _0362_
rlabel metal1 18814 20536 18814 20536 0 _0363_
rlabel metal1 19550 15504 19550 15504 0 _0364_
rlabel metal1 20654 13906 20654 13906 0 _0365_
rlabel metal1 20516 13838 20516 13838 0 _0366_
rlabel metal2 7682 39814 7682 39814 0 _0367_
rlabel metal1 7360 41582 7360 41582 0 _0368_
rlabel metal2 17250 40222 17250 40222 0 _0369_
rlabel metal1 13340 39814 13340 39814 0 _0370_
rlabel metal2 13570 39236 13570 39236 0 _0371_
rlabel metal1 12282 39610 12282 39610 0 _0372_
rlabel metal1 7682 41514 7682 41514 0 _0373_
rlabel metal1 7820 42806 7820 42806 0 _0374_
rlabel metal1 6026 45424 6026 45424 0 _0375_
rlabel metal2 25714 40698 25714 40698 0 _0376_
rlabel metal1 24380 40494 24380 40494 0 _0377_
rlabel metal1 27324 41582 27324 41582 0 _0378_
rlabel metal2 27094 34918 27094 34918 0 _0379_
rlabel metal2 25622 36278 25622 36278 0 _0380_
rlabel metal2 23598 35462 23598 35462 0 _0381_
rlabel metal2 26358 38250 26358 38250 0 _0382_
rlabel metal1 43240 23698 43240 23698 0 _0383_
rlabel metal2 42642 23460 42642 23460 0 _0384_
rlabel metal1 43746 25874 43746 25874 0 _0385_
rlabel metal1 38226 26418 38226 26418 0 _0386_
rlabel metal1 39652 26554 39652 26554 0 _0387_
rlabel metal1 38226 26350 38226 26350 0 _0388_
rlabel metal1 38870 26350 38870 26350 0 _0389_
rlabel metal1 4600 10234 4600 10234 0 _0390_
rlabel metal1 6624 13294 6624 13294 0 _0391_
rlabel metal2 4830 18428 4830 18428 0 _0392_
rlabel metal1 4554 18054 4554 18054 0 _0393_
rlabel metal1 4646 18292 4646 18292 0 _0394_
rlabel metal1 5060 18054 5060 18054 0 _0395_
rlabel metal1 6686 43690 6686 43690 0 _0396_
rlabel metal2 7130 43452 7130 43452 0 _0397_
rlabel metal2 6762 42534 6762 42534 0 _0398_
rlabel metal1 10580 42330 10580 42330 0 _0399_
rlabel via1 9706 44693 9706 44693 0 _0400_
rlabel metal1 9430 43724 9430 43724 0 _0401_
rlabel metal2 7682 45152 7682 45152 0 _0402_
rlabel metal1 8188 44846 8188 44846 0 _0403_
rlabel metal1 6118 44234 6118 44234 0 _0404_
rlabel metal1 6946 44200 6946 44200 0 _0405_
rlabel metal2 7130 44982 7130 44982 0 _0406_
rlabel metal1 6762 43112 6762 43112 0 _0407_
rlabel metal2 5934 42636 5934 42636 0 _0408_
rlabel metal2 22310 14960 22310 14960 0 _0409_
rlabel metal1 21390 15402 21390 15402 0 _0410_
rlabel metal1 20792 16558 20792 16558 0 _0411_
rlabel metal2 21114 18020 21114 18020 0 _0412_
rlabel metal1 22264 18054 22264 18054 0 _0413_
rlabel metal2 21942 14688 21942 14688 0 _0414_
rlabel metal2 22126 15266 22126 15266 0 _0415_
rlabel metal1 20194 15878 20194 15878 0 _0416_
rlabel metal1 20302 13226 20302 13226 0 _0417_
rlabel metal1 20838 13498 20838 13498 0 _0418_
rlabel metal1 40342 36754 40342 36754 0 _0419_
rlabel metal1 40756 36618 40756 36618 0 _0420_
rlabel metal1 40756 37434 40756 37434 0 _0421_
rlabel metal1 40296 35054 40296 35054 0 _0422_
rlabel metal1 40296 33082 40296 33082 0 _0423_
rlabel metal1 40296 32538 40296 32538 0 _0424_
rlabel metal1 40756 32878 40756 32878 0 _0425_
rlabel metal2 40250 34272 40250 34272 0 _0426_
rlabel metal1 39422 32912 39422 32912 0 _0427_
rlabel metal1 40940 36550 40940 36550 0 _0428_
rlabel metal2 40158 37604 40158 37604 0 _0429_
rlabel metal1 42052 37162 42052 37162 0 _0430_
rlabel metal1 42596 37230 42596 37230 0 _0431_
rlabel metal1 13432 25466 13432 25466 0 _0432_
rlabel metal1 15364 23698 15364 23698 0 _0433_
rlabel via1 14590 24922 14590 24922 0 _0434_
rlabel metal1 14996 24786 14996 24786 0 _0435_
rlabel metal2 13386 23392 13386 23392 0 _0436_
rlabel metal1 13321 21964 13321 21964 0 _0437_
rlabel metal1 13018 24786 13018 24786 0 _0438_
rlabel metal1 15594 23664 15594 23664 0 _0439_
rlabel metal1 15272 23290 15272 23290 0 _0440_
rlabel metal2 36846 20876 36846 20876 0 _0441_
rlabel metal1 37996 21114 37996 21114 0 _0442_
rlabel metal1 38134 20978 38134 20978 0 _0443_
rlabel metal2 37950 20604 37950 20604 0 _0444_
rlabel metal1 38870 21114 38870 21114 0 _0445_
rlabel metal2 39238 21386 39238 21386 0 _0446_
rlabel metal1 43332 44846 43332 44846 0 _0447_
rlabel metal1 43470 43418 43470 43418 0 _0448_
rlabel metal1 44666 42874 44666 42874 0 _0449_
rlabel metal1 45402 44812 45402 44812 0 _0450_
rlabel metal1 10764 12818 10764 12818 0 _0451_
rlabel metal2 8142 14076 8142 14076 0 _0452_
rlabel metal1 4830 12784 4830 12784 0 _0453_
rlabel metal1 6325 14382 6325 14382 0 _0454_
rlabel metal2 11914 11084 11914 11084 0 _0455_
rlabel metal1 11730 13940 11730 13940 0 _0456_
rlabel metal2 12650 13736 12650 13736 0 _0457_
rlabel metal2 14490 14212 14490 14212 0 _0458_
rlabel metal2 11178 14552 11178 14552 0 _0459_
rlabel metal1 11316 14586 11316 14586 0 _0460_
rlabel metal2 13754 14620 13754 14620 0 _0461_
rlabel metal1 11730 12920 11730 12920 0 _0462_
rlabel metal2 11086 13124 11086 13124 0 _0463_
rlabel metal2 8878 14314 8878 14314 0 _0464_
rlabel via1 9330 14314 9330 14314 0 _0465_
rlabel metal2 9154 15300 9154 15300 0 _0466_
rlabel metal2 8050 14722 8050 14722 0 _0467_
rlabel metal2 8970 15232 8970 15232 0 _0468_
rlabel metal1 7728 14382 7728 14382 0 _0469_
rlabel metal1 8510 12682 8510 12682 0 _0470_
rlabel metal1 8878 12138 8878 12138 0 _0471_
rlabel metal2 7130 11900 7130 11900 0 _0472_
rlabel metal1 8832 10710 8832 10710 0 _0473_
rlabel metal1 9062 10778 9062 10778 0 _0474_
rlabel metal2 4646 13379 4646 13379 0 _0475_
rlabel metal1 5658 14042 5658 14042 0 _0476_
rlabel metal1 3266 14348 3266 14348 0 _0477_
rlabel metal1 43654 31382 43654 31382 0 _0478_
rlabel metal1 43470 30226 43470 30226 0 _0479_
rlabel metal2 43286 28798 43286 28798 0 _0480_
rlabel metal2 44390 26316 44390 26316 0 _0481_
rlabel metal1 45402 33048 45402 33048 0 _0482_
rlabel metal1 43516 33082 43516 33082 0 _0483_
rlabel metal2 44574 32402 44574 32402 0 _0484_
rlabel metal2 45402 32368 45402 32368 0 _0485_
rlabel metal2 46046 32266 46046 32266 0 _0486_
rlabel metal2 42090 32674 42090 32674 0 _0487_
rlabel metal1 42596 32538 42596 32538 0 _0488_
rlabel metal2 41170 32572 41170 32572 0 _0489_
rlabel metal1 43194 31858 43194 31858 0 _0490_
rlabel metal1 42320 30362 42320 30362 0 _0491_
rlabel metal2 45310 28390 45310 28390 0 _0492_
rlabel metal1 45356 28186 45356 28186 0 _0493_
rlabel metal1 45908 29138 45908 29138 0 _0494_
rlabel metal1 43286 29206 43286 29206 0 _0495_
rlabel metal1 44084 29206 44084 29206 0 _0496_
rlabel metal2 43930 29444 43930 29444 0 _0497_
rlabel metal1 43332 27574 43332 27574 0 _0498_
rlabel metal1 42780 27370 42780 27370 0 _0499_
rlabel metal1 42228 27642 42228 27642 0 _0500_
rlabel metal3 2062 44948 2062 44948 0 clk
rlabel metal1 18906 24072 18906 24072 0 clknet_0_clk
rlabel metal1 5382 17646 5382 17646 0 clknet_1_0__leaf_clk
rlabel metal1 40940 17578 40940 17578 0 clknet_1_1__leaf_clk
rlabel metal2 2070 19312 2070 19312 0 clknet_leaf_0_clk
rlabel metal2 24610 42704 24610 42704 0 clknet_leaf_10_clk
rlabel metal1 36938 38318 36938 38318 0 clknet_leaf_11_clk
rlabel metal1 43286 41514 43286 41514 0 clknet_leaf_12_clk
rlabel metal1 36294 37230 36294 37230 0 clknet_leaf_13_clk
rlabel metal1 41676 31790 41676 31790 0 clknet_leaf_14_clk
rlabel metal1 37306 30158 37306 30158 0 clknet_leaf_15_clk
rlabel metal1 35190 28526 35190 28526 0 clknet_leaf_16_clk
rlabel metal1 33442 24650 33442 24650 0 clknet_leaf_17_clk
rlabel metal1 38226 24786 38226 24786 0 clknet_leaf_18_clk
rlabel metal1 40158 24820 40158 24820 0 clknet_leaf_19_clk
rlabel metal1 2944 21658 2944 21658 0 clknet_leaf_1_clk
rlabel metal1 44528 17170 44528 17170 0 clknet_leaf_20_clk
rlabel metal2 44482 10336 44482 10336 0 clknet_leaf_21_clk
rlabel metal1 32476 20366 32476 20366 0 clknet_leaf_22_clk
rlabel metal1 24794 24650 24794 24650 0 clknet_leaf_23_clk
rlabel metal1 20654 17646 20654 17646 0 clknet_leaf_24_clk
rlabel metal1 20838 14518 20838 14518 0 clknet_leaf_25_clk
rlabel metal1 11477 14314 11477 14314 0 clknet_leaf_26_clk
rlabel metal2 2714 10438 2714 10438 0 clknet_leaf_27_clk
rlabel metal1 13800 23154 13800 23154 0 clknet_leaf_2_clk
rlabel metal1 20746 25330 20746 25330 0 clknet_leaf_3_clk
rlabel metal2 5290 41072 5290 41072 0 clknet_leaf_4_clk
rlabel metal2 6762 45118 6762 45118 0 clknet_leaf_5_clk
rlabel metal2 12558 38080 12558 38080 0 clknet_leaf_6_clk
rlabel metal1 23690 42126 23690 42126 0 clknet_leaf_7_clk
rlabel metal2 23322 29376 23322 29376 0 clknet_leaf_8_clk
rlabel metal2 32338 37332 32338 37332 0 clknet_leaf_9_clk
rlabel metal2 8786 41650 8786 41650 0 clknet_opt_1_0_clk
rlabel metal2 44574 41140 44574 41140 0 clknet_opt_2_0_clk
rlabel metal2 42918 14892 42918 14892 0 clknet_opt_3_0_clk
rlabel metal1 12006 12716 12006 12716 0 counter10\[0\]
rlabel metal2 7406 17850 7406 17850 0 counter10\[10\]
rlabel metal2 7958 18564 7958 18564 0 counter10\[11\]
rlabel metal1 7682 18938 7682 18938 0 counter10\[12\]
rlabel metal2 7038 18292 7038 18292 0 counter10\[13\]
rlabel metal2 3542 18530 3542 18530 0 counter10\[14\]
rlabel metal1 3680 17850 3680 17850 0 counter10\[15\]
rlabel metal1 3726 18938 3726 18938 0 counter10\[16\]
rlabel metal1 4094 17306 4094 17306 0 counter10\[17\]
rlabel metal2 3450 20434 3450 20434 0 counter10\[18\]
rlabel metal1 4094 21012 4094 21012 0 counter10\[19\]
rlabel metal1 11224 13906 11224 13906 0 counter10\[1\]
rlabel metal2 4002 20842 4002 20842 0 counter10\[20\]
rlabel metal1 4370 20570 4370 20570 0 counter10\[21\]
rlabel metal1 3726 10030 3726 10030 0 counter10\[22\]
rlabel metal1 4508 10098 4508 10098 0 counter10\[23\]
rlabel metal2 4094 10336 4094 10336 0 counter10\[24\]
rlabel metal1 4600 10030 4600 10030 0 counter10\[25\]
rlabel metal2 6854 10336 6854 10336 0 counter10\[26\]
rlabel metal2 6946 10812 6946 10812 0 counter10\[27\]
rlabel metal2 11822 12954 11822 12954 0 counter10\[2\]
rlabel metal1 12052 12818 12052 12818 0 counter10\[3\]
rlabel metal1 9706 15062 9706 15062 0 counter10\[4\]
rlabel metal1 8510 14926 8510 14926 0 counter10\[5\]
rlabel metal1 8556 12818 8556 12818 0 counter10\[6\]
rlabel metal1 9016 12886 9016 12886 0 counter10\[7\]
rlabel metal1 4876 14042 4876 14042 0 counter10\[8\]
rlabel metal1 5658 13328 5658 13328 0 counter10\[9\]
rlabel metal1 44344 43962 44344 43962 0 counter2\[0\]
rlabel metal1 42182 40392 42182 40392 0 counter2\[10\]
rlabel metal2 41814 40324 41814 40324 0 counter2\[11\]
rlabel metal2 42182 41072 42182 41072 0 counter2\[12\]
rlabel metal2 42458 40698 42458 40698 0 counter2\[13\]
rlabel metal2 38870 40290 38870 40290 0 counter2\[14\]
rlabel metal1 38870 40596 38870 40596 0 counter2\[15\]
rlabel metal2 38778 41072 38778 41072 0 counter2\[16\]
rlabel metal2 39054 40698 39054 40698 0 counter2\[17\]
rlabel metal1 38226 37128 38226 37128 0 counter2\[18\]
rlabel metal2 38318 37740 38318 37740 0 counter2\[19\]
rlabel metal1 43976 43418 43976 43418 0 counter2\[1\]
rlabel metal2 38226 37536 38226 37536 0 counter2\[20\]
rlabel metal1 38686 37230 38686 37230 0 counter2\[21\]
rlabel metal1 34868 41242 34868 41242 0 counter2\[22\]
rlabel metal1 35006 41650 35006 41650 0 counter2\[23\]
rlabel metal2 35374 41888 35374 41888 0 counter2\[24\]
rlabel metal1 34868 41582 34868 41582 0 counter2\[25\]
rlabel metal1 43930 41242 43930 41242 0 counter2\[26\]
rlabel metal2 44666 41922 44666 41922 0 counter2\[27\]
rlabel metal1 38502 43656 38502 43656 0 counter2\[2\]
rlabel metal2 38686 43622 38686 43622 0 counter2\[3\]
rlabel metal2 38502 44336 38502 44336 0 counter2\[4\]
rlabel metal2 38778 43962 38778 43962 0 counter2\[5\]
rlabel metal1 41906 43656 41906 43656 0 counter2\[6\]
rlabel metal2 41998 43996 41998 43996 0 counter2\[7\]
rlabel metal2 41538 44608 41538 44608 0 counter2\[8\]
rlabel metal2 42182 44234 42182 44234 0 counter2\[9\]
rlabel metal2 37582 21726 37582 21726 0 counter3\[0\]
rlabel metal1 35466 21352 35466 21352 0 counter3\[10\]
rlabel metal1 35052 20570 35052 20570 0 counter3\[11\]
rlabel metal1 33396 25874 33396 25874 0 counter3\[12\]
rlabel metal1 29440 25874 29440 25874 0 counter3\[13\]
rlabel metal1 30084 20570 30084 20570 0 counter3\[14\]
rlabel metal1 30038 21114 30038 21114 0 counter3\[15\]
rlabel metal1 29624 26758 29624 26758 0 counter3\[16\]
rlabel metal1 30544 21318 30544 21318 0 counter3\[17\]
rlabel metal1 29486 25670 29486 25670 0 counter3\[18\]
rlabel metal1 29624 26214 29624 26214 0 counter3\[19\]
rlabel metal2 38226 21794 38226 21794 0 counter3\[1\]
rlabel metal1 31188 20570 31188 20570 0 counter3\[20\]
rlabel metal1 31510 23290 31510 23290 0 counter3\[21\]
rlabel metal2 33534 20400 33534 20400 0 counter3\[22\]
rlabel metal2 33718 19652 33718 19652 0 counter3\[23\]
rlabel metal2 31878 24412 31878 24412 0 counter3\[24\]
rlabel metal2 31694 24004 31694 24004 0 counter3\[25\]
rlabel metal1 31556 24378 31556 24378 0 counter3\[26\]
rlabel metal2 34638 24004 34638 24004 0 counter3\[27\]
rlabel metal2 39146 20910 39146 20910 0 counter3\[2\]
rlabel metal1 34638 24378 34638 24378 0 counter3\[3\]
rlabel metal1 34914 24242 34914 24242 0 counter3\[4\]
rlabel metal1 33994 20536 33994 20536 0 counter3\[5\]
rlabel metal2 33718 26078 33718 26078 0 counter3\[6\]
rlabel metal2 36294 21284 36294 21284 0 counter3\[7\]
rlabel metal1 33672 26758 33672 26758 0 counter3\[8\]
rlabel metal1 33258 27302 33258 27302 0 counter3\[9\]
rlabel metal1 15042 23086 15042 23086 0 counter4\[0\]
rlabel metal1 22218 27302 22218 27302 0 counter4\[10\]
rlabel metal2 22218 25670 22218 25670 0 counter4\[11\]
rlabel metal2 25254 26010 25254 26010 0 counter4\[12\]
rlabel metal1 25024 25942 25024 25942 0 counter4\[13\]
rlabel metal1 25668 26758 25668 26758 0 counter4\[14\]
rlabel metal1 24840 27302 24840 27302 0 counter4\[15\]
rlabel metal1 24288 29546 24288 29546 0 counter4\[16\]
rlabel metal1 24656 29682 24656 29682 0 counter4\[17\]
rlabel metal1 24794 29274 24794 29274 0 counter4\[18\]
rlabel metal2 24702 29920 24702 29920 0 counter4\[19\]
rlabel metal1 15180 23154 15180 23154 0 counter4\[1\]
rlabel metal1 18814 27098 18814 27098 0 counter4\[20\]
rlabel metal2 20102 28220 20102 28220 0 counter4\[21\]
rlabel metal1 20194 28084 20194 28084 0 counter4\[22\]
rlabel metal1 19182 27574 19182 27574 0 counter4\[23\]
rlabel metal1 18860 23630 18860 23630 0 counter4\[24\]
rlabel metal1 18676 23766 18676 23766 0 counter4\[25\]
rlabel metal2 18906 24310 18906 24310 0 counter4\[26\]
rlabel metal2 19182 24140 19182 24140 0 counter4\[27\]
rlabel metal2 12098 23222 12098 23222 0 counter4\[2\]
rlabel metal1 13386 23290 13386 23290 0 counter4\[3\]
rlabel metal1 24840 23290 24840 23290 0 counter4\[4\]
rlabel metal2 25806 23834 25806 23834 0 counter4\[5\]
rlabel metal1 25392 23494 25392 23494 0 counter4\[6\]
rlabel metal1 25944 23290 25944 23290 0 counter4\[7\]
rlabel metal1 21758 24922 21758 24922 0 counter4\[8\]
rlabel metal2 22126 25092 22126 25092 0 counter4\[9\]
rlabel metal1 40940 36142 40940 36142 0 counter5\[0\]
rlabel metal1 29670 32878 29670 32878 0 counter5\[10\]
rlabel metal1 31924 29274 31924 29274 0 counter5\[11\]
rlabel metal1 34684 35054 34684 35054 0 counter5\[12\]
rlabel metal1 35006 35156 35006 35156 0 counter5\[13\]
rlabel metal2 31786 30430 31786 30430 0 counter5\[14\]
rlabel metal1 34592 36006 34592 36006 0 counter5\[15\]
rlabel metal1 32200 30906 32200 30906 0 counter5\[16\]
rlabel metal1 32752 29818 32752 29818 0 counter5\[17\]
rlabel metal1 35098 34714 35098 34714 0 counter5\[18\]
rlabel metal2 36478 31926 36478 31926 0 counter5\[19\]
rlabel metal2 41262 33796 41262 33796 0 counter5\[1\]
rlabel metal1 36156 30906 36156 30906 0 counter5\[20\]
rlabel metal2 36110 32096 36110 32096 0 counter5\[21\]
rlabel metal1 35328 30022 35328 30022 0 counter5\[22\]
rlabel metal2 31786 33762 31786 33762 0 counter5\[23\]
rlabel metal1 32890 34068 32890 34068 0 counter5\[24\]
rlabel metal2 33074 33898 33074 33898 0 counter5\[25\]
rlabel metal2 32522 33524 32522 33524 0 counter5\[26\]
rlabel metal2 28934 32402 28934 32402 0 counter5\[27\]
rlabel via1 39338 33830 39338 33830 0 counter5\[2\]
rlabel metal1 41354 36720 41354 36720 0 counter5\[3\]
rlabel metal2 41630 37468 41630 37468 0 counter5\[4\]
rlabel metal2 37582 34340 37582 34340 0 counter5\[5\]
rlabel metal1 29854 32980 29854 32980 0 counter5\[6\]
rlabel metal2 29762 33456 29762 33456 0 counter5\[7\]
rlabel metal1 37628 36006 37628 36006 0 counter5\[8\]
rlabel metal2 37766 34748 37766 34748 0 counter5\[9\]
rlabel metal2 21114 16864 21114 16864 0 counter6\[0\]
rlabel metal1 18676 17306 18676 17306 0 counter6\[10\]
rlabel metal2 18814 18462 18814 18462 0 counter6\[11\]
rlabel metal1 18584 18054 18584 18054 0 counter6\[12\]
rlabel metal1 18998 17850 18998 17850 0 counter6\[13\]
rlabel metal1 22218 21012 22218 21012 0 counter6\[14\]
rlabel metal2 22126 20434 22126 20434 0 counter6\[15\]
rlabel metal2 21482 21216 21482 21216 0 counter6\[16\]
rlabel metal2 22402 20740 22402 20740 0 counter6\[17\]
rlabel metal1 18538 20298 18538 20298 0 counter6\[18\]
rlabel metal1 18032 20026 18032 20026 0 counter6\[19\]
rlabel metal2 22126 17748 22126 17748 0 counter6\[1\]
rlabel metal1 18400 21114 18400 21114 0 counter6\[20\]
rlabel metal1 18998 21454 18998 21454 0 counter6\[21\]
rlabel metal1 16146 16456 16146 16456 0 counter6\[22\]
rlabel metal1 16100 16218 16100 16218 0 counter6\[23\]
rlabel metal2 16146 16864 16146 16864 0 counter6\[24\]
rlabel metal2 16514 16116 16514 16116 0 counter6\[25\]
rlabel metal2 17158 14042 17158 14042 0 counter6\[26\]
rlabel metal1 17894 14484 17894 14484 0 counter6\[27\]
rlabel metal2 22954 18020 22954 18020 0 counter6\[2\]
rlabel metal2 22218 15300 22218 15300 0 counter6\[3\]
rlabel metal1 19918 15402 19918 15402 0 counter6\[4\]
rlabel metal1 19044 15130 19044 15130 0 counter6\[5\]
rlabel metal1 14490 20026 14490 20026 0 counter6\[6\]
rlabel metal2 14766 19924 14766 19924 0 counter6\[7\]
rlabel metal1 14996 20230 14996 20230 0 counter6\[8\]
rlabel metal2 15686 20230 15686 20230 0 counter6\[9\]
rlabel metal1 9798 42228 9798 42228 0 counter7\[0\]
rlabel metal2 13294 42704 13294 42704 0 counter7\[10\]
rlabel metal2 13202 41140 13202 41140 0 counter7\[11\]
rlabel metal1 12788 41514 12788 41514 0 counter7\[12\]
rlabel metal1 16813 40494 16813 40494 0 counter7\[13\]
rlabel metal2 16790 41072 16790 41072 0 counter7\[14\]
rlabel metal2 16882 40732 16882 40732 0 counter7\[15\]
rlabel metal2 16790 40018 16790 40018 0 counter7\[16\]
rlabel metal2 13938 38148 13938 38148 0 counter7\[17\]
rlabel metal1 12880 38522 12880 38522 0 counter7\[18\]
rlabel metal1 13110 37434 13110 37434 0 counter7\[19\]
rlabel metal2 9890 42874 9890 42874 0 counter7\[1\]
rlabel metal1 12144 37978 12144 37978 0 counter7\[20\]
rlabel metal1 11224 39406 11224 39406 0 counter7\[21\]
rlabel metal2 11178 40256 11178 40256 0 counter7\[22\]
rlabel metal1 10764 39406 10764 39406 0 counter7\[23\]
rlabel metal2 6946 40086 6946 40086 0 counter7\[24\]
rlabel metal2 6670 39780 6670 39780 0 counter7\[25\]
rlabel metal2 7314 39032 7314 39032 0 counter7\[26\]
rlabel metal1 7314 38522 7314 38522 0 counter7\[27\]
rlabel metal1 9476 45050 9476 45050 0 counter7\[2\]
rlabel metal1 9200 45526 9200 45526 0 counter7\[3\]
rlabel metal2 5934 44540 5934 44540 0 counter7\[4\]
rlabel via1 6302 43282 6302 43282 0 counter7\[5\]
rlabel metal1 7774 42194 7774 42194 0 counter7\[6\]
rlabel metal2 7406 38726 7406 38726 0 counter7\[7\]
rlabel metal1 7084 37094 7084 37094 0 counter7\[8\]
rlabel metal1 12742 41242 12742 41242 0 counter7\[9\]
rlabel metal1 31786 37298 31786 37298 0 counter8\[0\]
rlabel metal1 26542 33966 26542 33966 0 counter8\[10\]
rlabel metal2 26634 34544 26634 34544 0 counter8\[11\]
rlabel metal2 24886 37060 24886 37060 0 counter8\[12\]
rlabel metal2 24610 38080 24610 38080 0 counter8\[13\]
rlabel metal2 24702 37468 24702 37468 0 counter8\[14\]
rlabel metal1 24610 37128 24610 37128 0 counter8\[15\]
rlabel metal1 22908 34986 22908 34986 0 counter8\[16\]
rlabel metal2 23322 34884 23322 34884 0 counter8\[17\]
rlabel metal1 23184 34170 23184 34170 0 counter8\[18\]
rlabel metal2 20102 34986 20102 34986 0 counter8\[19\]
rlabel metal2 31878 37468 31878 37468 0 counter8\[1\]
rlabel metal1 25898 41446 25898 41446 0 counter8\[20\]
rlabel metal1 25760 43622 25760 43622 0 counter8\[21\]
rlabel metal1 25530 41208 25530 41208 0 counter8\[22\]
rlabel metal1 25484 41990 25484 41990 0 counter8\[23\]
rlabel metal2 22954 40596 22954 40596 0 counter8\[24\]
rlabel metal1 22448 41446 22448 41446 0 counter8\[25\]
rlabel metal1 23230 41990 23230 41990 0 counter8\[26\]
rlabel metal2 23598 40324 23598 40324 0 counter8\[27\]
rlabel metal1 31970 37196 31970 37196 0 counter8\[2\]
rlabel metal1 32062 37332 32062 37332 0 counter8\[3\]
rlabel metal1 28566 36856 28566 36856 0 counter8\[4\]
rlabel metal1 27692 38318 27692 38318 0 counter8\[5\]
rlabel metal1 27830 40086 27830 40086 0 counter8\[6\]
rlabel metal1 27462 41242 27462 41242 0 counter8\[7\]
rlabel metal1 26128 33082 26128 33082 0 counter8\[8\]
rlabel metal2 26726 34374 26726 34374 0 counter8\[9\]
rlabel metal1 44528 31790 44528 31790 0 counter9\[0\]
rlabel metal1 38732 23834 38732 23834 0 counter9\[10\]
rlabel metal1 39882 27030 39882 27030 0 counter9\[11\]
rlabel metal1 40342 26860 40342 26860 0 counter9\[12\]
rlabel metal1 40158 26758 40158 26758 0 counter9\[13\]
rlabel metal2 40526 27132 40526 27132 0 counter9\[14\]
rlabel metal1 37490 28152 37490 28152 0 counter9\[15\]
rlabel metal2 37674 28220 37674 28220 0 counter9\[16\]
rlabel metal1 37030 27574 37030 27574 0 counter9\[17\]
rlabel metal1 37260 27098 37260 27098 0 counter9\[18\]
rlabel metal2 41906 21522 41906 21522 0 counter9\[19\]
rlabel metal1 42872 32538 42872 32538 0 counter9\[1\]
rlabel metal2 43378 21828 43378 21828 0 counter9\[20\]
rlabel metal1 42964 22202 42964 22202 0 counter9\[21\]
rlabel metal2 43746 21556 43746 21556 0 counter9\[22\]
rlabel metal2 41630 23868 41630 23868 0 counter9\[23\]
rlabel metal2 40894 23834 40894 23834 0 counter9\[24\]
rlabel metal2 41538 23392 41538 23392 0 counter9\[25\]
rlabel metal2 41722 24106 41722 24106 0 counter9\[26\]
rlabel metal2 36938 24310 36938 24310 0 counter9\[27\]
rlabel metal1 42458 32402 42458 32402 0 counter9\[2\]
rlabel metal1 44022 31858 44022 31858 0 counter9\[3\]
rlabel metal1 45264 28050 45264 28050 0 counter9\[4\]
rlabel via1 44574 29155 44574 29155 0 counter9\[5\]
rlabel metal1 43516 28186 43516 28186 0 counter9\[6\]
rlabel metal2 43470 26690 43470 26690 0 counter9\[7\]
rlabel metal1 44160 25874 44160 25874 0 counter9\[8\]
rlabel metal1 37214 24582 37214 24582 0 counter9\[9\]
rlabel metal1 44436 13498 44436 13498 0 counter\[0\]
rlabel metal1 43792 11322 43792 11322 0 counter\[10\]
rlabel metal1 41308 15130 41308 15130 0 counter\[11\]
rlabel metal1 41722 14586 41722 14586 0 counter\[12\]
rlabel metal1 41814 14042 41814 14042 0 counter\[13\]
rlabel metal1 41676 15674 41676 15674 0 counter\[14\]
rlabel metal1 38686 17544 38686 17544 0 counter\[15\]
rlabel metal2 38870 17884 38870 17884 0 counter\[16\]
rlabel metal1 38824 17306 38824 17306 0 counter\[17\]
rlabel metal2 38962 18122 38962 18122 0 counter\[18\]
rlabel metal1 45954 17170 45954 17170 0 counter\[19\]
rlabel metal2 45310 13974 45310 13974 0 counter\[1\]
rlabel metal1 46414 17068 46414 17068 0 counter\[20\]
rlabel metal2 46322 17510 46322 17510 0 counter\[21\]
rlabel metal2 46598 16966 46598 16966 0 counter\[22\]
rlabel metal1 41814 17306 41814 17306 0 counter\[23\]
rlabel metal1 42734 18156 42734 18156 0 counter\[24\]
rlabel metal2 42642 18326 42642 18326 0 counter\[25\]
rlabel metal2 44022 17646 44022 17646 0 counter\[26\]
rlabel metal1 45126 13838 45126 13838 0 counter\[27\]
rlabel metal2 45586 14348 45586 14348 0 counter\[2\]
rlabel metal1 39560 11322 39560 11322 0 counter\[3\]
rlabel metal1 40986 11628 40986 11628 0 counter\[4\]
rlabel metal2 40894 12070 40894 12070 0 counter\[5\]
rlabel metal2 41446 11526 41446 11526 0 counter\[6\]
rlabel metal2 44022 10914 44022 10914 0 counter\[7\]
rlabel metal1 44068 10234 44068 10234 0 counter\[8\]
rlabel metal2 45862 10948 45862 10948 0 counter\[9\]
rlabel metal2 58282 3417 58282 3417 0 cout1
rlabel metal2 46 1520 46 1520 0 cout10
rlabel metal1 50140 57562 50140 57562 0 cout2
rlabel metal2 42550 1520 42550 1520 0 cout3
rlabel metal2 1794 22355 1794 22355 0 cout4
rlabel via2 58282 49045 58282 49045 0 cout5
rlabel metal2 21298 1520 21298 1520 0 cout6
rlabel metal1 6578 57562 6578 57562 0 cout7
rlabel metal1 28474 57562 28474 57562 0 cout8
rlabel metal2 58282 26673 58282 26673 0 cout9
rlabel metal1 57822 3502 57822 3502 0 net1
rlabel metal2 58098 26316 58098 26316 0 net10
rlabel metal2 33534 40902 33534 40902 0 net100
rlabel metal1 37720 36754 37720 36754 0 net101
rlabel via1 36666 37842 36666 37842 0 net102
rlabel metal1 36462 38250 36462 38250 0 net103
rlabel metal2 36662 36958 36662 36958 0 net104
rlabel metal1 37720 39610 37720 39610 0 net105
rlabel via1 37393 41582 37393 41582 0 net106
rlabel metal1 36830 40426 36830 40426 0 net107
rlabel metal1 37342 40018 37342 40018 0 net108
rlabel metal2 41354 40358 41354 40358 0 net109
rlabel metal2 22494 39950 22494 39950 0 net11
rlabel via1 40705 41582 40705 41582 0 net110
rlabel metal1 40418 40086 40418 40086 0 net111
rlabel metal1 40664 39610 40664 39610 0 net112
rlabel metal1 41303 44778 41303 44778 0 net113
rlabel metal1 40475 45526 40475 45526 0 net114
rlabel metal1 41119 44370 41119 44370 0 net115
rlabel via1 40337 43758 40337 43758 0 net116
rlabel via1 37761 44370 37761 44370 0 net117
rlabel metal2 36294 44574 36294 44574 0 net118
rlabel via1 37761 43350 37761 43350 0 net119
rlabel metal1 21804 42126 21804 42126 0 net12
rlabel metal1 36554 43690 36554 43690 0 net120
rlabel metal1 33580 23290 33580 23290 0 net121
rlabel metal1 29936 24174 29936 24174 0 net122
rlabel metal1 30631 23766 30631 23766 0 net123
rlabel metal2 29854 24242 29854 24242 0 net124
rlabel metal1 32368 19414 32368 19414 0 net125
rlabel via1 32609 20910 32609 20910 0 net126
rlabel metal1 29608 23018 29608 23018 0 net127
rlabel metal2 30038 20230 30038 20230 0 net128
rlabel metal1 28377 26350 28377 26350 0 net129
rlabel metal2 21114 41310 21114 41310 0 net13
rlabel metal1 28004 25874 28004 25874 0 net130
rlabel metal1 28832 21522 28832 21522 0 net131
rlabel metal1 27554 26996 27554 26996 0 net132
rlabel metal2 30498 20400 30498 20400 0 net133
rlabel metal2 28290 20230 28290 20230 0 net134
rlabel metal2 27370 26962 27370 26962 0 net135
rlabel metal1 31827 26962 31827 26962 0 net136
rlabel metal2 36754 20706 36754 20706 0 net137
rlabel metal2 34178 21318 34178 21318 0 net138
rlabel via1 31965 27370 31965 27370 0 net139
rlabel via1 22305 40018 22305 40018 0 net14
rlabel metal1 32506 27030 32506 27030 0 net140
rlabel metal1 35236 20026 35236 20026 0 net141
rlabel metal1 32568 25874 32568 25874 0 net142
rlabel via1 32885 20502 32885 20502 0 net143
rlabel metal1 33340 24786 33340 24786 0 net144
rlabel metal1 33621 24174 33621 24174 0 net145
rlabel metal1 18671 24786 18671 24786 0 net146
rlabel via1 17337 25262 17337 25262 0 net147
rlabel metal1 17096 23766 17096 23766 0 net148
rlabel metal1 17378 24174 17378 24174 0 net149
rlabel via1 24237 42262 24237 42262 0 net15
rlabel via1 17337 27438 17337 27438 0 net150
rlabel via1 18349 28118 18349 28118 0 net151
rlabel via1 17337 28526 17337 28526 0 net152
rlabel metal2 16790 27438 16790 27438 0 net153
rlabel via1 23593 30294 23593 30294 0 net154
rlabel metal1 23214 29206 23214 29206 0 net155
rlabel metal2 25162 30770 25162 30770 0 net156
rlabel metal1 22478 29546 22478 29546 0 net157
rlabel metal1 24890 27438 24890 27438 0 net158
rlabel metal1 25249 27030 25249 27030 0 net159
rlabel metal1 24564 40698 24564 40698 0 net16
rlabel metal1 23133 27030 23133 27030 0 net160
rlabel via1 24881 26350 24881 26350 0 net161
rlabel via1 21109 25262 21109 25262 0 net162
rlabel via1 21017 27438 21017 27438 0 net163
rlabel via1 21017 24106 21017 24106 0 net164
rlabel via1 20373 24786 20373 24786 0 net165
rlabel via1 24881 23086 24881 23086 0 net166
rlabel via1 24053 23698 24053 23698 0 net167
rlabel metal2 23322 23868 23322 23868 0 net168
rlabel metal1 22995 23018 22995 23018 0 net169
rlabel via1 24881 43758 24881 43758 0 net17
rlabel metal1 27728 31790 27728 31790 0 net170
rlabel via1 31413 32810 31413 32810 0 net171
rlabel metal1 31142 33592 31142 33592 0 net172
rlabel via1 31229 33966 31229 33966 0 net173
rlabel metal1 31050 32402 31050 32402 0 net174
rlabel metal1 36355 30294 36355 30294 0 net175
rlabel metal1 35323 31790 35323 31790 0 net176
rlabel metal1 35277 30634 35277 30634 0 net177
rlabel metal1 35042 31314 35042 31314 0 net178
rlabel metal1 33948 34170 33948 34170 0 net179
rlabel metal1 24456 41514 24456 41514 0 net18
rlabel metal1 31827 29614 31827 29614 0 net180
rlabel via1 30861 30634 30861 30634 0 net181
rlabel via1 33253 36142 33253 36142 0 net182
rlabel metal1 31091 30294 31091 30294 0 net183
rlabel metal1 33667 35054 33667 35054 0 net184
rlabel metal1 32614 35700 32614 35700 0 net185
rlabel via1 30309 29138 30309 29138 0 net186
rlabel via1 28193 33558 28193 33558 0 net187
rlabel via1 36565 35054 36565 35054 0 net188
rlabel metal1 37301 36074 37301 36074 0 net189
rlabel metal1 21635 34646 21635 34646 0 net19
rlabel metal1 28469 33966 28469 33966 0 net190
rlabel metal1 28004 32878 28004 32878 0 net191
rlabel via1 36473 33898 36473 33898 0 net192
rlabel metal1 15854 14314 15854 14314 0 net193
rlabel via1 16049 13294 16049 13294 0 net194
rlabel metal1 16141 15470 16141 15470 0 net195
rlabel via1 14669 17238 14669 17238 0 net196
rlabel metal1 14520 16150 14520 16150 0 net197
rlabel metal2 14122 16286 14122 16286 0 net198
rlabel metal1 17383 21590 17383 21590 0 net199
rlabel metal1 1748 9894 1748 9894 0 net2
rlabel metal2 22034 33694 22034 33694 0 net20
rlabel metal1 17015 20842 17015 20842 0 net200
rlabel metal1 16790 22406 16790 22406 0 net201
rlabel metal1 16866 20502 16866 20502 0 net202
rlabel metal1 20184 20434 20184 20434 0 net203
rlabel via1 20373 21590 20373 21590 0 net204
rlabel metal1 21247 19822 21247 19822 0 net205
rlabel metal1 20787 20910 20787 20910 0 net206
rlabel metal1 18211 17578 18211 17578 0 net207
rlabel metal2 17066 18054 17066 18054 0 net208
rlabel metal2 16330 18462 16330 18462 0 net209
rlabel metal2 22310 34374 22310 34374 0 net21
rlabel metal1 17383 17238 17383 17238 0 net210
rlabel metal1 14536 18938 14536 18938 0 net211
rlabel metal1 13795 20434 13795 20434 0 net212
rlabel via1 13657 19346 13657 19346 0 net213
rlabel metal1 12691 19754 12691 19754 0 net214
rlabel metal1 8336 38318 8336 38318 0 net215
rlabel via1 5561 38318 5561 38318 0 net216
rlabel via1 5561 39406 5561 39406 0 net217
rlabel via1 5561 40494 5561 40494 0 net218
rlabel metal1 9328 39406 9328 39406 0 net219
rlabel metal1 21190 34986 21190 34986 0 net22
rlabel metal2 8602 40868 8602 40868 0 net220
rlabel via1 9425 40494 9425 40494 0 net221
rlabel metal1 10345 37910 10345 37910 0 net222
rlabel metal2 11914 36958 11914 36958 0 net223
rlabel metal1 11633 38250 11633 38250 0 net224
rlabel metal1 12098 37876 12098 37876 0 net225
rlabel via1 15313 39406 15313 39406 0 net226
rlabel metal1 14858 39610 14858 39610 0 net227
rlabel metal1 16003 41582 16003 41582 0 net228
rlabel metal1 14848 40494 14848 40494 0 net229
rlabel metal1 22908 36754 22908 36754 0 net23
rlabel metal2 11178 41310 11178 41310 0 net230
rlabel via1 12093 40494 12093 40494 0 net231
rlabel metal2 12374 43486 12374 43486 0 net232
rlabel metal1 13672 41106 13672 41106 0 net233
rlabel via1 5837 37230 5837 37230 0 net234
rlabel metal2 7038 38284 7038 38284 0 net235
rlabel via1 23593 37910 23593 37910 0 net24
rlabel metal1 23322 38522 23322 38522 0 net25
rlabel metal2 23782 36550 23782 36550 0 net26
rlabel metal1 26123 35054 26123 35054 0 net27
rlabel metal2 26174 33660 26174 33660 0 net28
rlabel metal1 24472 33966 24472 33966 0 net29
rlabel metal1 48484 57426 48484 57426 0 net3
rlabel metal1 24840 32402 24840 32402 0 net30
rlabel metal2 36386 24480 36386 24480 0 net31
rlabel via1 40337 25262 40337 25262 0 net32
rlabel metal1 40296 23290 40296 23290 0 net33
rlabel via1 38589 24854 38589 24854 0 net34
rlabel metal1 40332 24786 40332 24786 0 net35
rlabel via1 42637 20910 42637 20910 0 net36
rlabel via1 41625 21998 41625 21998 0 net37
rlabel via1 42913 21522 42913 21522 0 net38
rlabel via1 40797 20910 40797 20910 0 net39
rlabel metal1 42274 9350 42274 9350 0 net4
rlabel metal2 37030 27200 37030 27200 0 net40
rlabel via1 35461 27438 35461 27438 0 net41
rlabel metal2 36202 28696 36202 28696 0 net42
rlabel metal1 34638 28084 34638 28084 0 net43
rlabel metal1 38226 26894 38226 26894 0 net44
rlabel metal1 38727 28118 38727 28118 0 net45
rlabel via1 38681 27030 38681 27030 0 net46
rlabel metal1 39279 27370 39279 27370 0 net47
rlabel metal1 37260 23290 37260 23290 0 net48
rlabel metal2 36294 25024 36294 25024 0 net49
rlabel metal2 1610 22202 1610 22202 0 net5
rlabel metal1 5796 9554 5796 9554 0 net50
rlabel via1 5745 10030 5745 10030 0 net51
rlabel metal1 3859 10642 3859 10642 0 net52
rlabel metal1 2622 10608 2622 10608 0 net53
rlabel metal1 3813 11730 3813 11730 0 net54
rlabel via1 2249 11050 2249 11050 0 net55
rlabel via1 5570 20502 5570 20502 0 net56
rlabel via1 2893 20502 2893 20502 0 net57
rlabel metal2 2162 20638 2162 20638 0 net58
rlabel via1 2341 19822 2341 19822 0 net59
rlabel metal2 45586 47260 45586 47260 0 net6
rlabel metal2 4002 16966 4002 16966 0 net60
rlabel via1 2341 18734 2341 18734 0 net61
rlabel metal1 3169 17646 3169 17646 0 net62
rlabel metal1 2208 17102 2208 17102 0 net63
rlabel metal1 8065 17578 8065 17578 0 net64
rlabel metal1 6348 19278 6348 19278 0 net65
rlabel metal1 6348 18190 6348 18190 0 net66
rlabel metal1 5285 17238 5285 17238 0 net67
rlabel metal1 44477 13974 44477 13974 0 net68
rlabel viali 42913 17238 42913 17238 0 net69
rlabel metal1 21712 9894 21712 9894 0 net7
rlabel via1 40981 18734 40981 18734 0 net70
rlabel metal2 40986 17510 40986 17510 0 net71
rlabel metal1 40424 17170 40424 17170 0 net72
rlabel metal1 45070 16558 45070 16558 0 net73
rlabel via1 44477 18326 44477 18326 0 net74
rlabel metal1 44983 17238 44983 17238 0 net75
rlabel metal1 44431 16150 44431 16150 0 net76
rlabel via1 37853 18666 37853 18666 0 net77
rlabel metal1 37566 17238 37566 17238 0 net78
rlabel metal1 38543 18258 38543 18258 0 net79
rlabel metal1 6762 57426 6762 57426 0 net8
rlabel via1 36933 17578 36933 17578 0 net80
rlabel metal1 40475 15470 40475 15470 0 net81
rlabel metal1 40751 13974 40751 13974 0 net82
rlabel via1 40337 14382 40337 14382 0 net83
rlabel via1 39601 14994 39601 14994 0 net84
rlabel via1 42453 11050 42453 11050 0 net85
rlabel via1 44753 10710 44753 10710 0 net86
rlabel metal2 42826 9758 42826 9758 0 net87
rlabel metal1 42412 10574 42412 10574 0 net88
rlabel metal1 39590 11050 39590 11050 0 net89
rlabel metal1 28658 57426 28658 57426 0 net9
rlabel metal1 39739 12886 39739 12886 0 net90
rlabel via1 39325 11798 39325 11798 0 net91
rlabel via1 38405 11050 38405 11050 0 net92
rlabel metal2 45862 14790 45862 14790 0 net93
rlabel metal1 43649 14314 43649 14314 0 net94
rlabel viali 43557 41582 43557 41582 0 net95
rlabel metal1 44957 41174 44957 41174 0 net96
rlabel metal1 35052 41106 35052 41106 0 net97
rlabel metal2 35098 42432 35098 42432 0 net98
rlabel via1 33897 42194 33897 42194 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
