VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO posoco2000
  CLASS BLOCK ;
  FOREIGN posoco2000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.840 299.000 7.440 ;
    END
  END clk
  PIN segm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.440 299.000 72.040 ;
    END
  END segm[0]
  PIN segm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1.000 183.910 4.000 ;
    END
  END segm[1]
  PIN segm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 299.000 204.640 ;
    END
  END segm[2]
  PIN segm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 299.000 269.240 ;
    END
  END segm[3]
  PIN segm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 261.840 4.000 262.440 ;
    END
  END segm[4]
  PIN segm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 296.000 209.670 299.000 ;
    END
  END segm[5]
  PIN segm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END segm[6]
  PIN segm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 296.000 84.090 299.000 ;
    END
  END segm[7]
  PIN sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1.000 248.310 4.000 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1.000 61.550 4.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 296.000 145.270 299.000 ;
    END
  END sel[2]
  PIN sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 64.640 4.000 65.240 ;
    END
  END sel[3]
  PIN sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 129.240 4.000 129.840 ;
    END
  END sel[4]
  PIN sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 296.000 270.850 299.000 ;
    END
  END sel[5]
  PIN sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1.000 122.730 4.000 ;
    END
  END sel[6]
  PIN sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 193.840 4.000 194.440 ;
    END
  END sel[7]
  PIN sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 296.000 22.910 299.000 ;
    END
  END sel[8]
  PIN sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 299.000 136.640 ;
    END
  END sel[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 294.400 288.560 ;
      LAYER met2 ;
        RECT 0.100 295.720 22.350 296.000 ;
        RECT 23.190 295.720 83.530 296.000 ;
        RECT 84.370 295.720 144.710 296.000 ;
        RECT 145.550 295.720 209.110 296.000 ;
        RECT 209.950 295.720 270.290 296.000 ;
        RECT 271.130 295.720 292.010 296.000 ;
        RECT 0.100 4.280 292.010 295.720 ;
        RECT 0.650 4.000 60.990 4.280 ;
        RECT 61.830 4.000 122.170 4.280 ;
        RECT 123.010 4.000 183.350 4.280 ;
        RECT 184.190 4.000 247.750 4.280 ;
        RECT 248.590 4.000 292.010 4.280 ;
      LAYER met3 ;
        RECT 4.000 269.640 296.000 288.485 ;
        RECT 4.000 268.240 295.600 269.640 ;
        RECT 4.000 262.840 296.000 268.240 ;
        RECT 4.400 261.440 296.000 262.840 ;
        RECT 4.000 205.040 296.000 261.440 ;
        RECT 4.000 203.640 295.600 205.040 ;
        RECT 4.000 194.840 296.000 203.640 ;
        RECT 4.400 193.440 296.000 194.840 ;
        RECT 4.000 137.040 296.000 193.440 ;
        RECT 4.000 135.640 295.600 137.040 ;
        RECT 4.000 130.240 296.000 135.640 ;
        RECT 4.400 128.840 296.000 130.240 ;
        RECT 4.000 72.440 296.000 128.840 ;
        RECT 4.000 71.040 295.600 72.440 ;
        RECT 4.000 65.640 296.000 71.040 ;
        RECT 4.400 64.240 296.000 65.640 ;
        RECT 4.000 7.840 296.000 64.240 ;
        RECT 4.000 6.975 295.600 7.840 ;
  END
END posoco2000
END LIBRARY

