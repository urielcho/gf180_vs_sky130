magic
tech sky130A
magscale 1 2
timestamp 1671750178
<< viali >>
rect 1685 57545 1719 57579
rect 9229 57545 9263 57579
rect 14473 57545 14507 57579
rect 19533 57545 19567 57579
rect 24685 57545 24719 57579
rect 35725 57545 35759 57579
rect 41521 57545 41555 57579
rect 46673 57545 46707 57579
rect 53113 57545 53147 57579
rect 58265 57545 58299 57579
rect 2789 57477 2823 57511
rect 29929 57477 29963 57511
rect 30481 57477 30515 57511
rect 1869 57409 1903 57443
rect 9413 57409 9447 57443
rect 13737 57409 13771 57443
rect 14289 57409 14323 57443
rect 19717 57409 19751 57443
rect 24869 57409 24903 57443
rect 35541 57409 35575 57443
rect 40877 57409 40911 57443
rect 41337 57409 41371 57443
rect 46029 57409 46063 57443
rect 46489 57409 46523 57443
rect 52929 57409 52963 57443
rect 58081 57409 58115 57443
rect 20269 57341 20303 57375
rect 2881 57205 2915 57239
rect 9873 57205 9907 57239
rect 25329 57205 25363 57239
rect 30573 57205 30607 57239
rect 52285 57205 52319 57239
rect 57437 57205 57471 57239
rect 2605 57001 2639 57035
rect 35265 57001 35299 57035
rect 58265 57001 58299 57035
rect 35081 56797 35115 56831
rect 58081 56797 58115 56831
rect 1961 56661 1995 56695
rect 35725 56661 35759 56695
rect 57621 56661 57655 56695
rect 1869 51969 1903 52003
rect 58081 51969 58115 52003
rect 1685 51765 1719 51799
rect 2329 51765 2363 51799
rect 57437 51765 57471 51799
rect 58265 51765 58299 51799
rect 29745 47957 29779 47991
rect 25053 47685 25087 47719
rect 28273 47617 28307 47651
rect 28457 47617 28491 47651
rect 28733 47617 28767 47651
rect 33425 47617 33459 47651
rect 25605 47549 25639 47583
rect 29285 47549 29319 47583
rect 33241 47549 33275 47583
rect 22385 47413 22419 47447
rect 23029 47413 23063 47447
rect 23673 47413 23707 47447
rect 24961 47413 24995 47447
rect 30297 47413 30331 47447
rect 31309 47413 31343 47447
rect 33977 47413 34011 47447
rect 28733 47209 28767 47243
rect 32597 47209 32631 47243
rect 26709 47141 26743 47175
rect 27905 47141 27939 47175
rect 23213 47073 23247 47107
rect 31769 47073 31803 47107
rect 22017 47005 22051 47039
rect 22201 47005 22235 47039
rect 23029 47005 23063 47039
rect 23489 47005 23523 47039
rect 24869 47005 24903 47039
rect 25145 47005 25179 47039
rect 26525 47005 26559 47039
rect 26801 47005 26835 47039
rect 27721 47005 27755 47039
rect 27905 47005 27939 47039
rect 29101 47005 29135 47039
rect 30849 47005 30883 47039
rect 31033 47005 31067 47039
rect 22109 46937 22143 46971
rect 23397 46937 23431 46971
rect 24961 46937 24995 46971
rect 27537 46937 27571 46971
rect 30297 46937 30331 46971
rect 33425 46937 33459 46971
rect 23949 46869 23983 46903
rect 25329 46869 25363 46903
rect 25881 46869 25915 46903
rect 26341 46869 26375 46903
rect 28549 46869 28583 46903
rect 28733 46869 28767 46903
rect 33333 46869 33367 46903
rect 33977 46869 34011 46903
rect 30113 46665 30147 46699
rect 24869 46597 24903 46631
rect 33517 46597 33551 46631
rect 1869 46529 1903 46563
rect 21281 46529 21315 46563
rect 21465 46529 21499 46563
rect 22293 46529 22327 46563
rect 23305 46529 23339 46563
rect 25053 46529 25087 46563
rect 25237 46529 25271 46563
rect 26157 46529 26191 46563
rect 26341 46529 26375 46563
rect 26617 46529 26651 46563
rect 28089 46529 28123 46563
rect 28457 46529 28491 46563
rect 29929 46529 29963 46563
rect 30205 46529 30239 46563
rect 31125 46529 31159 46563
rect 32413 46529 32447 46563
rect 33241 46529 33275 46563
rect 24317 46461 24351 46495
rect 22477 46393 22511 46427
rect 24041 46393 24075 46427
rect 25145 46393 25179 46427
rect 26433 46393 26467 46427
rect 31585 46393 31619 46427
rect 1685 46325 1719 46359
rect 2329 46325 2363 46359
rect 21465 46325 21499 46359
rect 23121 46325 23155 46359
rect 23857 46325 23891 46359
rect 25881 46325 25915 46359
rect 26249 46325 26283 46359
rect 27537 46325 27571 46359
rect 28457 46325 28491 46359
rect 28641 46325 28675 46359
rect 29285 46325 29319 46359
rect 29745 46325 29779 46359
rect 30941 46325 30975 46359
rect 32689 46325 32723 46359
rect 34161 46325 34195 46359
rect 34713 46325 34747 46359
rect 30757 46053 30791 46087
rect 25881 45985 25915 46019
rect 28825 45985 28859 46019
rect 30665 45985 30699 46019
rect 31861 45985 31895 46019
rect 22569 45917 22603 45951
rect 22845 45917 22879 45951
rect 23765 45917 23799 45951
rect 23949 45917 23983 45951
rect 24777 45917 24811 45951
rect 24961 45917 24995 45951
rect 25053 45917 25087 45951
rect 26525 45917 26559 45951
rect 26985 45917 27019 45951
rect 27629 45917 27663 45951
rect 27721 45917 27755 45951
rect 27905 45917 27939 45951
rect 27997 45917 28031 45951
rect 29009 45917 29043 45951
rect 29929 45917 29963 45951
rect 30205 45917 30239 45951
rect 30573 45917 30607 45951
rect 32137 45917 32171 45951
rect 32597 45917 32631 45951
rect 32965 45917 32999 45951
rect 33701 45917 33735 45951
rect 33885 45917 33919 45951
rect 58081 45917 58115 45951
rect 21557 45849 21591 45883
rect 21925 45849 21959 45883
rect 24593 45849 24627 45883
rect 27445 45849 27479 45883
rect 29193 45849 29227 45883
rect 20453 45781 20487 45815
rect 21005 45781 21039 45815
rect 22385 45781 22419 45815
rect 22753 45781 22787 45815
rect 23857 45781 23891 45815
rect 26525 45781 26559 45815
rect 33885 45781 33919 45815
rect 34897 45781 34931 45815
rect 57529 45781 57563 45815
rect 58265 45781 58299 45815
rect 22293 45577 22327 45611
rect 30941 45577 30975 45611
rect 31033 45577 31067 45611
rect 25697 45509 25731 45543
rect 27261 45509 27295 45543
rect 20821 45441 20855 45475
rect 21005 45441 21039 45475
rect 21281 45441 21315 45475
rect 22201 45441 22235 45475
rect 22477 45441 22511 45475
rect 23305 45441 23339 45475
rect 24593 45441 24627 45475
rect 25053 45441 25087 45475
rect 25513 45441 25547 45475
rect 25789 45441 25823 45475
rect 26433 45441 26467 45475
rect 26617 45441 26651 45475
rect 28549 45441 28583 45475
rect 28825 45441 28859 45475
rect 29009 45441 29043 45475
rect 30205 45441 30239 45475
rect 30849 45441 30883 45475
rect 31217 45441 31251 45475
rect 32598 45441 32632 45475
rect 32965 45441 32999 45475
rect 33609 45441 33643 45475
rect 34437 45441 34471 45475
rect 21097 45373 21131 45407
rect 21189 45373 21223 45407
rect 23581 45373 23615 45407
rect 24777 45373 24811 45407
rect 24869 45373 24903 45407
rect 33057 45373 33091 45407
rect 24685 45305 24719 45339
rect 27629 45305 27663 45339
rect 30665 45305 30699 45339
rect 32413 45305 32447 45339
rect 21465 45237 21499 45271
rect 22661 45237 22695 45271
rect 23121 45237 23155 45271
rect 23489 45237 23523 45271
rect 24409 45237 24443 45271
rect 25789 45237 25823 45271
rect 26525 45237 26559 45271
rect 27721 45237 27755 45271
rect 28365 45237 28399 45271
rect 29745 45237 29779 45271
rect 30113 45237 30147 45271
rect 31677 45237 31711 45271
rect 35909 45237 35943 45271
rect 21465 45033 21499 45067
rect 23305 45033 23339 45067
rect 34161 45033 34195 45067
rect 34897 45033 34931 45067
rect 28273 44965 28307 44999
rect 32137 44965 32171 44999
rect 20085 44897 20119 44931
rect 23664 44897 23698 44931
rect 23765 44897 23799 44931
rect 27261 44897 27295 44931
rect 32873 44897 32907 44931
rect 20637 44829 20671 44863
rect 21373 44829 21407 44863
rect 21465 44829 21499 44863
rect 22477 44829 22511 44863
rect 22569 44829 22603 44863
rect 22753 44829 22787 44863
rect 22845 44829 22879 44863
rect 23489 44829 23523 44863
rect 23581 44829 23615 44863
rect 25605 44829 25639 44863
rect 25697 44829 25731 44863
rect 25789 44829 25823 44863
rect 25973 44829 26007 44863
rect 26709 44829 26743 44863
rect 27629 44829 27663 44863
rect 28089 44829 28123 44863
rect 29009 44829 29043 44863
rect 29193 44829 29227 44863
rect 29929 44829 29963 44863
rect 30113 44829 30147 44863
rect 32045 44829 32079 44863
rect 32229 44829 32263 44863
rect 32965 44829 32999 44863
rect 33609 44829 33643 44863
rect 24869 44761 24903 44795
rect 27445 44761 27479 44795
rect 29745 44761 29779 44795
rect 31033 44761 31067 44795
rect 19533 44693 19567 44727
rect 21097 44693 21131 44727
rect 22293 44693 22327 44727
rect 25329 44693 25363 44727
rect 29101 44693 29135 44727
rect 31309 44693 31343 44727
rect 25329 44489 25363 44523
rect 20453 44421 20487 44455
rect 21189 44421 21223 44455
rect 34621 44421 34655 44455
rect 34821 44421 34855 44455
rect 19257 44353 19291 44387
rect 20913 44353 20947 44387
rect 21005 44353 21039 44387
rect 22017 44353 22051 44387
rect 22201 44353 22235 44387
rect 22753 44353 22787 44387
rect 22937 44353 22971 44387
rect 24133 44353 24167 44387
rect 24317 44353 24351 44387
rect 25145 44353 25179 44387
rect 25421 44353 25455 44387
rect 26249 44353 26283 44387
rect 27261 44353 27295 44387
rect 27445 44353 27479 44387
rect 27905 44353 27939 44387
rect 28089 44353 28123 44387
rect 28917 44353 28951 44387
rect 29101 44353 29135 44387
rect 29561 44353 29595 44387
rect 29745 44353 29779 44387
rect 30297 44353 30331 44387
rect 30481 44353 30515 44387
rect 31309 44353 31343 44387
rect 32505 44353 32539 44387
rect 33425 44353 33459 44387
rect 33977 44353 34011 44387
rect 19441 44285 19475 44319
rect 24501 44285 24535 44319
rect 26525 44285 26559 44319
rect 30389 44285 30423 44319
rect 33241 44285 33275 44319
rect 22845 44217 22879 44251
rect 33885 44217 33919 44251
rect 19073 44149 19107 44183
rect 21189 44149 21223 44183
rect 22201 44149 22235 44183
rect 23581 44149 23615 44183
rect 24961 44149 24995 44183
rect 26341 44149 26375 44183
rect 26433 44149 26467 44183
rect 27261 44149 27295 44183
rect 28089 44149 28123 44183
rect 29101 44149 29135 44183
rect 29653 44149 29687 44183
rect 31033 44149 31067 44183
rect 32413 44149 32447 44183
rect 34805 44149 34839 44183
rect 34989 44149 35023 44183
rect 21373 43945 21407 43979
rect 23857 43945 23891 43979
rect 30849 43945 30883 43979
rect 32689 43945 32723 43979
rect 33517 43945 33551 43979
rect 18429 43877 18463 43911
rect 25973 43877 26007 43911
rect 30113 43877 30147 43911
rect 31861 43877 31895 43911
rect 25881 43809 25915 43843
rect 26157 43809 26191 43843
rect 27721 43809 27755 43843
rect 30757 43809 30791 43843
rect 34989 43809 35023 43843
rect 18705 43741 18739 43775
rect 18889 43741 18923 43775
rect 20085 43741 20119 43775
rect 20361 43741 20395 43775
rect 20545 43741 20579 43775
rect 21005 43741 21039 43775
rect 21189 43741 21223 43775
rect 21465 43741 21499 43775
rect 23673 43741 23707 43775
rect 24041 43741 24075 43775
rect 25605 43741 25639 43775
rect 26433 43741 26467 43775
rect 27169 43741 27203 43775
rect 27261 43741 27295 43775
rect 27445 43741 27479 43775
rect 27537 43741 27571 43775
rect 28181 43741 28215 43775
rect 28365 43741 28399 43775
rect 28825 43741 28859 43775
rect 29009 43741 29043 43775
rect 29929 43741 29963 43775
rect 30021 43741 30055 43775
rect 30205 43741 30239 43775
rect 31033 43741 31067 43775
rect 31677 43741 31711 43775
rect 34897 43741 34931 43775
rect 35081 43741 35115 43775
rect 20177 43673 20211 43707
rect 20269 43673 20303 43707
rect 22109 43673 22143 43707
rect 22477 43673 22511 43707
rect 32597 43673 32631 43707
rect 33793 43673 33827 43707
rect 18613 43605 18647 43639
rect 19901 43605 19935 43639
rect 23489 43605 23523 43639
rect 24777 43605 24811 43639
rect 28273 43605 28307 43639
rect 28917 43605 28951 43639
rect 29745 43605 29779 43639
rect 31217 43605 31251 43639
rect 35633 43605 35667 43639
rect 23397 43401 23431 43435
rect 25421 43401 25455 43435
rect 20913 43333 20947 43367
rect 23673 43333 23707 43367
rect 27321 43333 27355 43367
rect 27537 43333 27571 43367
rect 28181 43333 28215 43367
rect 31217 43333 31251 43367
rect 32413 43333 32447 43367
rect 18521 43265 18555 43299
rect 18889 43265 18923 43299
rect 19073 43265 19107 43299
rect 20085 43265 20119 43299
rect 20177 43265 20211 43299
rect 20269 43265 20303 43299
rect 20453 43265 20487 43299
rect 21097 43265 21131 43299
rect 21189 43265 21223 43299
rect 22477 43265 22511 43299
rect 22569 43265 22603 43299
rect 22753 43265 22787 43299
rect 22845 43265 22879 43299
rect 23535 43265 23569 43299
rect 23765 43265 23799 43299
rect 23948 43265 23982 43299
rect 24041 43265 24075 43299
rect 24501 43265 24535 43299
rect 24685 43265 24719 43299
rect 25605 43265 25639 43299
rect 25697 43265 25731 43299
rect 25881 43265 25915 43299
rect 28273 43265 28307 43299
rect 28549 43265 28583 43299
rect 29009 43265 29043 43299
rect 29377 43265 29411 43299
rect 29745 43265 29779 43299
rect 30481 43265 30515 43299
rect 33701 43265 33735 43299
rect 35173 43265 35207 43299
rect 33885 43197 33919 43231
rect 19349 43129 19383 43163
rect 20913 43129 20947 43163
rect 25789 43129 25823 43163
rect 26525 43129 26559 43163
rect 27169 43129 27203 43163
rect 34713 43129 34747 43163
rect 19257 43061 19291 43095
rect 19809 43061 19843 43095
rect 22293 43061 22327 43095
rect 24685 43061 24719 43095
rect 27353 43061 27387 43095
rect 30573 43061 30607 43095
rect 31309 43061 31343 43095
rect 32689 43061 32723 43095
rect 25053 42857 25087 42891
rect 30021 42857 30055 42891
rect 31217 42857 31251 42891
rect 31401 42857 31435 42891
rect 28089 42789 28123 42823
rect 33701 42789 33735 42823
rect 23305 42721 23339 42755
rect 25513 42721 25547 42755
rect 25697 42721 25731 42755
rect 25973 42721 26007 42755
rect 27169 42721 27203 42755
rect 28273 42721 28307 42755
rect 28733 42721 28767 42755
rect 31493 42721 31527 42755
rect 20453 42653 20487 42687
rect 20545 42653 20579 42687
rect 20729 42653 20763 42687
rect 20821 42653 20855 42687
rect 21465 42653 21499 42687
rect 21741 42653 21775 42687
rect 22201 42653 22235 42687
rect 22477 42653 22511 42687
rect 25789 42653 25823 42687
rect 25881 42653 25915 42687
rect 27077 42653 27111 42687
rect 27261 42653 27295 42687
rect 27353 42653 27387 42687
rect 27997 42653 28031 42687
rect 28917 42653 28951 42687
rect 29929 42653 29963 42687
rect 30113 42653 30147 42687
rect 31585 42653 31619 42687
rect 32505 42653 32539 42687
rect 32689 42653 32723 42687
rect 33425 42653 33459 42687
rect 34161 42653 34195 42687
rect 34897 42653 34931 42687
rect 19809 42585 19843 42619
rect 21373 42585 21407 42619
rect 22661 42585 22695 42619
rect 29101 42585 29135 42619
rect 35081 42585 35115 42619
rect 20269 42517 20303 42551
rect 22293 42517 22327 42551
rect 24041 42517 24075 42551
rect 27537 42517 27571 42551
rect 28273 42517 28307 42551
rect 32597 42517 32631 42551
rect 35265 42517 35299 42551
rect 35817 42517 35851 42551
rect 20453 42313 20487 42347
rect 27721 42313 27755 42347
rect 28641 42245 28675 42279
rect 19717 42177 19751 42211
rect 20361 42177 20395 42211
rect 20637 42177 20671 42211
rect 21373 42177 21407 42211
rect 22293 42177 22327 42211
rect 22385 42177 22419 42211
rect 22477 42177 22511 42211
rect 22661 42177 22695 42211
rect 23673 42177 23707 42211
rect 24409 42177 24443 42211
rect 24593 42177 24627 42211
rect 25053 42177 25087 42211
rect 25237 42177 25271 42211
rect 25881 42177 25915 42211
rect 26065 42177 26099 42211
rect 27718 42177 27752 42211
rect 28917 42177 28951 42211
rect 29009 42177 29043 42211
rect 29101 42177 29135 42211
rect 29285 42177 29319 42211
rect 30389 42177 30423 42211
rect 30481 42177 30515 42211
rect 30665 42177 30699 42211
rect 31401 42177 31435 42211
rect 31566 42177 31600 42211
rect 31677 42177 31711 42211
rect 31769 42177 31803 42211
rect 32505 42177 32539 42211
rect 32781 42177 32815 42211
rect 33885 42177 33919 42211
rect 33977 42177 34011 42211
rect 34069 42177 34103 42211
rect 34265 42177 34299 42211
rect 19625 42109 19659 42143
rect 19809 42109 19843 42143
rect 23397 42109 23431 42143
rect 23581 42109 23615 42143
rect 23765 42109 23799 42143
rect 23857 42109 23891 42143
rect 28181 42109 28215 42143
rect 22017 42041 22051 42075
rect 28089 42041 28123 42075
rect 30573 42041 30607 42075
rect 33609 42041 33643 42075
rect 19441 41973 19475 42007
rect 20821 41973 20855 42007
rect 24593 41973 24627 42007
rect 25145 41973 25179 42007
rect 25697 41973 25731 42007
rect 26065 41973 26099 42007
rect 26617 41973 26651 42007
rect 27537 41973 27571 42007
rect 30205 41973 30239 42007
rect 31217 41973 31251 42007
rect 32321 41973 32355 42007
rect 32689 41973 32723 42007
rect 34805 41973 34839 42007
rect 23673 41769 23707 41803
rect 23857 41769 23891 41803
rect 26801 41769 26835 41803
rect 30665 41769 30699 41803
rect 34989 41769 35023 41803
rect 21833 41701 21867 41735
rect 24685 41701 24719 41735
rect 32505 41701 32539 41735
rect 20085 41633 20119 41667
rect 35173 41633 35207 41667
rect 21925 41565 21959 41599
rect 22385 41565 22419 41599
rect 25329 41565 25363 41599
rect 25421 41565 25455 41599
rect 25605 41565 25639 41599
rect 25697 41565 25731 41599
rect 27077 41565 27111 41599
rect 27169 41565 27203 41599
rect 27261 41565 27295 41599
rect 27445 41565 27479 41599
rect 28549 41565 28583 41599
rect 28641 41565 28675 41599
rect 29009 41565 29043 41599
rect 29745 41565 29779 41599
rect 29929 41565 29963 41599
rect 30757 41565 30791 41599
rect 30849 41565 30883 41599
rect 31585 41565 31619 41599
rect 32689 41565 32723 41599
rect 32965 41565 32999 41599
rect 33609 41565 33643 41599
rect 34897 41565 34931 41599
rect 35633 41565 35667 41599
rect 21649 41497 21683 41531
rect 23489 41497 23523 41531
rect 23705 41497 23739 41531
rect 28825 41497 28859 41531
rect 28917 41497 28951 41531
rect 30573 41497 30607 41531
rect 33425 41497 33459 41531
rect 33793 41497 33827 41531
rect 20545 41429 20579 41463
rect 21097 41429 21131 41463
rect 21925 41429 21959 41463
rect 22569 41429 22603 41463
rect 25145 41429 25179 41463
rect 26341 41429 26375 41463
rect 27905 41429 27939 41463
rect 29193 41429 29227 41463
rect 29837 41429 29871 41463
rect 32873 41429 32907 41463
rect 35173 41429 35207 41463
rect 35725 41429 35759 41463
rect 36369 41429 36403 41463
rect 23029 41225 23063 41259
rect 23197 41225 23231 41259
rect 26249 41225 26283 41259
rect 31493 41225 31527 41259
rect 32521 41225 32555 41259
rect 23397 41157 23431 41191
rect 26401 41157 26435 41191
rect 26617 41157 26651 41191
rect 29561 41157 29595 41191
rect 32321 41157 32355 41191
rect 19349 41089 19383 41123
rect 20085 41089 20119 41123
rect 20177 41089 20211 41123
rect 20913 41089 20947 41123
rect 21097 41089 21131 41123
rect 21373 41089 21407 41123
rect 22201 41089 22235 41123
rect 22477 41089 22511 41123
rect 24041 41089 24075 41123
rect 24225 41089 24259 41123
rect 24961 41089 24995 41123
rect 25145 41089 25179 41123
rect 25421 41089 25455 41123
rect 25697 41089 25731 41123
rect 27445 41089 27479 41123
rect 27537 41089 27571 41123
rect 29377 41089 29411 41123
rect 29745 41089 29779 41123
rect 30205 41089 30239 41123
rect 33517 41089 33551 41123
rect 33701 41089 33735 41123
rect 33793 41089 33827 41123
rect 33977 41089 34011 41123
rect 34437 41089 34471 41123
rect 20453 41021 20487 41055
rect 21189 41021 21223 41055
rect 22385 41021 22419 41055
rect 24133 41021 24167 41055
rect 24317 41021 24351 41055
rect 24501 41021 24535 41055
rect 27261 41021 27295 41055
rect 20361 40953 20395 40987
rect 21281 40953 21315 40987
rect 22293 40953 22327 40987
rect 25329 40953 25363 40987
rect 30757 40953 30791 40987
rect 33609 40953 33643 40987
rect 18705 40885 18739 40919
rect 19901 40885 19935 40919
rect 22017 40885 22051 40919
rect 23213 40885 23247 40919
rect 26433 40885 26467 40919
rect 27353 40885 27387 40919
rect 28273 40885 28307 40919
rect 28917 40885 28951 40919
rect 32505 40885 32539 40919
rect 32689 40885 32723 40919
rect 33333 40885 33367 40919
rect 20177 40681 20211 40715
rect 24685 40681 24719 40715
rect 28549 40681 28583 40715
rect 33885 40681 33919 40715
rect 25237 40613 25271 40647
rect 25881 40613 25915 40647
rect 18521 40545 18555 40579
rect 20269 40545 20303 40579
rect 23857 40545 23891 40579
rect 27077 40545 27111 40579
rect 27261 40545 27295 40579
rect 27353 40545 27387 40579
rect 30941 40545 30975 40579
rect 1869 40477 1903 40511
rect 2329 40477 2363 40511
rect 18245 40477 18279 40511
rect 18337 40477 18371 40511
rect 19807 40477 19841 40511
rect 21741 40477 21775 40511
rect 21833 40477 21867 40511
rect 22017 40477 22051 40511
rect 22109 40477 22143 40511
rect 22937 40477 22971 40511
rect 23029 40477 23063 40511
rect 23213 40477 23247 40511
rect 23305 40477 23339 40511
rect 23765 40477 23799 40511
rect 23949 40477 23983 40511
rect 24593 40477 24627 40511
rect 24777 40477 24811 40511
rect 27169 40477 27203 40511
rect 28181 40477 28215 40511
rect 29745 40477 29779 40511
rect 30665 40477 30699 40511
rect 31761 40477 31795 40511
rect 31861 40477 31895 40511
rect 32045 40477 32079 40511
rect 32137 40477 32171 40511
rect 32597 40477 32631 40511
rect 32781 40477 32815 40511
rect 33241 40477 33275 40511
rect 33425 40477 33459 40511
rect 33885 40477 33919 40511
rect 34069 40477 34103 40511
rect 58081 40477 58115 40511
rect 17785 40409 17819 40443
rect 21557 40409 21591 40443
rect 28549 40409 28583 40443
rect 32689 40409 32723 40443
rect 1685 40341 1719 40375
rect 18521 40341 18555 40375
rect 19625 40341 19659 40375
rect 19809 40341 19843 40375
rect 21097 40341 21131 40375
rect 22753 40341 22787 40375
rect 26433 40341 26467 40375
rect 27537 40341 27571 40375
rect 28733 40341 28767 40375
rect 30297 40341 30331 40375
rect 30757 40341 30791 40375
rect 31585 40341 31619 40375
rect 33333 40341 33367 40375
rect 34989 40341 35023 40375
rect 35633 40341 35667 40375
rect 36093 40341 36127 40375
rect 57621 40341 57655 40375
rect 58265 40341 58299 40375
rect 19894 40137 19928 40171
rect 22661 40137 22695 40171
rect 23305 40137 23339 40171
rect 30005 40137 30039 40171
rect 35357 40137 35391 40171
rect 17325 40069 17359 40103
rect 19809 40069 19843 40103
rect 19993 40069 20027 40103
rect 23397 40069 23431 40103
rect 28917 40069 28951 40103
rect 30205 40069 30239 40103
rect 17785 40001 17819 40035
rect 17969 40001 18003 40035
rect 18429 40001 18463 40035
rect 18613 40001 18647 40035
rect 19717 40001 19751 40035
rect 20913 40001 20947 40035
rect 22201 40001 22235 40035
rect 23489 40001 23523 40035
rect 24133 40001 24167 40035
rect 25027 40001 25061 40035
rect 25237 40001 25271 40035
rect 26341 40001 26375 40035
rect 26525 40001 26559 40035
rect 27537 40001 27571 40035
rect 28825 40001 28859 40035
rect 29009 40001 29043 40035
rect 29193 40001 29227 40035
rect 29285 40001 29319 40035
rect 31309 40001 31343 40035
rect 32321 40001 32355 40035
rect 32505 40001 32539 40035
rect 32597 40001 32631 40035
rect 32689 40001 32723 40035
rect 36001 40001 36035 40035
rect 17877 39933 17911 39967
rect 23121 39933 23155 39967
rect 24409 39933 24443 39967
rect 25145 39933 25179 39967
rect 25329 39933 25363 39967
rect 26617 39933 26651 39967
rect 27353 39933 27387 39967
rect 27445 39933 27479 39967
rect 27629 39933 27663 39967
rect 31217 39933 31251 39967
rect 33609 39933 33643 39967
rect 33885 39933 33919 39967
rect 35909 39933 35943 39967
rect 29837 39865 29871 39899
rect 18521 39797 18555 39831
rect 18797 39797 18831 39831
rect 21465 39797 21499 39831
rect 22385 39797 22419 39831
rect 23213 39797 23247 39831
rect 23949 39797 23983 39831
rect 24317 39797 24351 39831
rect 24869 39797 24903 39831
rect 26157 39797 26191 39831
rect 27169 39797 27203 39831
rect 28641 39797 28675 39831
rect 30021 39797 30055 39831
rect 30941 39797 30975 39831
rect 31309 39797 31343 39831
rect 32965 39797 32999 39831
rect 36277 39797 36311 39831
rect 18521 39593 18555 39627
rect 26157 39593 26191 39627
rect 27537 39593 27571 39627
rect 28549 39593 28583 39627
rect 32597 39593 32631 39627
rect 25145 39525 25179 39559
rect 27905 39525 27939 39559
rect 17785 39457 17819 39491
rect 21097 39457 21131 39491
rect 22661 39457 22695 39491
rect 30665 39457 30699 39491
rect 32781 39457 32815 39491
rect 32873 39457 32907 39491
rect 35725 39457 35759 39491
rect 36093 39457 36127 39491
rect 37473 39457 37507 39491
rect 20177 39389 20211 39423
rect 20269 39389 20303 39423
rect 20729 39389 20763 39423
rect 20821 39389 20855 39423
rect 21373 39389 21407 39423
rect 22385 39389 22419 39423
rect 22569 39389 22603 39423
rect 22753 39389 22787 39423
rect 22937 39389 22971 39423
rect 23581 39389 23615 39423
rect 23765 39389 23799 39423
rect 24869 39389 24903 39423
rect 25881 39389 25915 39423
rect 26157 39389 26191 39423
rect 26617 39389 26651 39423
rect 26801 39389 26835 39423
rect 27721 39389 27755 39423
rect 27813 39389 27847 39423
rect 27997 39389 28031 39423
rect 28687 39389 28721 39423
rect 28917 39389 28951 39423
rect 29100 39389 29134 39423
rect 29193 39389 29227 39423
rect 29745 39389 29779 39423
rect 29929 39389 29963 39423
rect 30573 39389 30607 39423
rect 30757 39389 30791 39423
rect 31309 39389 31343 39423
rect 32965 39389 32999 39423
rect 33057 39389 33091 39423
rect 34897 39389 34931 39423
rect 18505 39321 18539 39355
rect 18705 39321 18739 39355
rect 22201 39321 22235 39355
rect 25145 39321 25179 39355
rect 26065 39321 26099 39355
rect 28825 39321 28859 39355
rect 30113 39321 30147 39355
rect 16497 39253 16531 39287
rect 17325 39253 17359 39287
rect 18337 39253 18371 39287
rect 23397 39253 23431 39287
rect 24961 39253 24995 39287
rect 26709 39253 26743 39287
rect 32137 39253 32171 39287
rect 33701 39253 33735 39287
rect 34253 39253 34287 39287
rect 18153 39049 18187 39083
rect 18705 39049 18739 39083
rect 20269 39049 20303 39083
rect 21373 39049 21407 39083
rect 32321 39049 32355 39083
rect 33885 39049 33919 39083
rect 36277 39049 36311 39083
rect 16865 38981 16899 39015
rect 19257 38981 19291 39015
rect 22385 38981 22419 39015
rect 28181 38981 28215 39015
rect 28365 38981 28399 39015
rect 31401 38981 31435 39015
rect 31493 38981 31527 39015
rect 32689 38981 32723 39015
rect 16129 38913 16163 38947
rect 16313 38913 16347 38947
rect 17068 38913 17102 38947
rect 17233 38913 17267 38947
rect 17325 38913 17359 38947
rect 17785 38913 17819 38947
rect 17969 38913 18003 38947
rect 20453 38913 20487 38947
rect 20545 38913 20579 38947
rect 22201 38913 22235 38947
rect 22293 38913 22327 38947
rect 22569 38913 22603 38947
rect 22661 38913 22695 38947
rect 23489 38913 23523 38947
rect 23582 38913 23616 38947
rect 23765 38913 23799 38947
rect 23857 38913 23891 38947
rect 23995 38913 24029 38947
rect 25053 38913 25087 38947
rect 25237 38913 25271 38947
rect 25421 38913 25455 38947
rect 26249 38913 26283 38947
rect 26341 38913 26375 38947
rect 26617 38913 26651 38947
rect 27445 38913 27479 38947
rect 28457 38913 28491 38947
rect 30021 38913 30055 38947
rect 30205 38913 30239 38947
rect 30297 38913 30331 38947
rect 30481 38913 30515 38947
rect 31309 38913 31343 38947
rect 31677 38913 31711 38947
rect 32505 38913 32539 38947
rect 32597 38913 32631 38947
rect 32873 38913 32907 38947
rect 32965 38913 32999 38947
rect 34161 38913 34195 38947
rect 35265 38913 35299 38947
rect 20637 38845 20671 38879
rect 20729 38845 20763 38879
rect 24961 38845 24995 38879
rect 27353 38845 27387 38879
rect 27537 38845 27571 38879
rect 27629 38845 27663 38879
rect 30665 38845 30699 38879
rect 34069 38845 34103 38879
rect 34253 38845 34287 38879
rect 34345 38845 34379 38879
rect 35173 38845 35207 38879
rect 28181 38777 28215 38811
rect 29009 38777 29043 38811
rect 30389 38777 30423 38811
rect 16221 38709 16255 38743
rect 19809 38709 19843 38743
rect 22017 38709 22051 38743
rect 24133 38709 24167 38743
rect 26065 38709 26099 38743
rect 26525 38709 26559 38743
rect 27169 38709 27203 38743
rect 29469 38709 29503 38743
rect 31125 38709 31159 38743
rect 34897 38709 34931 38743
rect 35081 38709 35115 38743
rect 35817 38709 35851 38743
rect 17785 38505 17819 38539
rect 18337 38505 18371 38539
rect 18521 38505 18555 38539
rect 22017 38505 22051 38539
rect 28641 38505 28675 38539
rect 30757 38505 30791 38539
rect 24869 38437 24903 38471
rect 30297 38437 30331 38471
rect 32965 38437 32999 38471
rect 16405 38369 16439 38403
rect 16589 38369 16623 38403
rect 19993 38369 20027 38403
rect 21925 38369 21959 38403
rect 26157 38369 26191 38403
rect 26801 38369 26835 38403
rect 27261 38369 27295 38403
rect 30573 38369 30607 38403
rect 32321 38369 32355 38403
rect 33241 38369 33275 38403
rect 33358 38369 33392 38403
rect 33517 38369 33551 38403
rect 35173 38369 35207 38403
rect 16313 38301 16347 38335
rect 16497 38301 16531 38335
rect 17601 38301 17635 38335
rect 17877 38301 17911 38335
rect 19441 38301 19475 38335
rect 19901 38301 19935 38335
rect 20545 38301 20579 38335
rect 20913 38301 20947 38335
rect 21373 38301 21407 38335
rect 21833 38301 21867 38335
rect 22155 38301 22189 38335
rect 22293 38301 22327 38335
rect 22753 38301 22787 38335
rect 22937 38301 22971 38335
rect 23673 38301 23707 38335
rect 24593 38301 24627 38335
rect 26065 38301 26099 38335
rect 26985 38301 27019 38335
rect 27445 38301 27479 38335
rect 28825 38301 28859 38335
rect 28917 38301 28951 38335
rect 29101 38301 29135 38335
rect 29193 38301 29227 38335
rect 30389 38301 30423 38335
rect 30849 38301 30883 38335
rect 32505 38301 32539 38335
rect 18705 38233 18739 38267
rect 23857 38233 23891 38267
rect 35449 38233 35483 38267
rect 37197 38233 37231 38267
rect 16129 38165 16163 38199
rect 17325 38165 17359 38199
rect 18505 38165 18539 38199
rect 22753 38165 22787 38199
rect 24041 38165 24075 38199
rect 25053 38165 25087 38199
rect 25605 38165 25639 38199
rect 29745 38165 29779 38199
rect 30481 38165 30515 38199
rect 31309 38165 31343 38199
rect 34161 38165 34195 38199
rect 17877 37961 17911 37995
rect 18705 37961 18739 37995
rect 19625 37961 19659 37995
rect 21373 37961 21407 37995
rect 28549 37961 28583 37995
rect 31493 37961 31527 37995
rect 33241 37961 33275 37995
rect 34253 37961 34287 37995
rect 34713 37961 34747 37995
rect 35357 37961 35391 37995
rect 17693 37893 17727 37927
rect 23181 37893 23215 37927
rect 23397 37893 23431 37927
rect 26157 37893 26191 37927
rect 15485 37825 15519 37859
rect 15669 37825 15703 37859
rect 17969 37825 18003 37859
rect 18797 37825 18831 37859
rect 19809 37825 19843 37859
rect 19993 37825 20027 37859
rect 20453 37825 20487 37859
rect 20729 37825 20763 37859
rect 22201 37825 22235 37859
rect 22385 37825 22419 37859
rect 23857 37825 23891 37859
rect 24593 37825 24627 37859
rect 24777 37825 24811 37859
rect 25651 37825 25685 37859
rect 25789 37825 25823 37859
rect 27169 37825 27203 37859
rect 27353 37825 27387 37859
rect 27445 37825 27479 37859
rect 27721 37825 27755 37859
rect 28733 37825 28767 37859
rect 28917 37825 28951 37859
rect 29561 37825 29595 37859
rect 29699 37825 29733 37859
rect 34069 37825 34103 37859
rect 35173 37825 35207 37859
rect 22109 37757 22143 37791
rect 22293 37757 22327 37791
rect 26065 37757 26099 37791
rect 27629 37757 27663 37791
rect 29929 37757 29963 37791
rect 33885 37757 33919 37791
rect 35081 37757 35115 37791
rect 17693 37689 17727 37723
rect 25513 37689 25547 37723
rect 29837 37689 29871 37723
rect 35817 37689 35851 37723
rect 15485 37621 15519 37655
rect 17233 37621 17267 37655
rect 22569 37621 22603 37655
rect 23029 37621 23063 37655
rect 23213 37621 23247 37655
rect 24041 37621 24075 37655
rect 24685 37621 24719 37655
rect 28917 37621 28951 37655
rect 30389 37621 30423 37655
rect 31033 37621 31067 37655
rect 32781 37621 32815 37655
rect 18889 37417 18923 37451
rect 23857 37417 23891 37451
rect 28089 37417 28123 37451
rect 30757 37417 30791 37451
rect 33977 37417 34011 37451
rect 31677 37349 31711 37383
rect 35541 37349 35575 37383
rect 15761 37281 15795 37315
rect 18337 37281 18371 37315
rect 23765 37281 23799 37315
rect 25329 37281 25363 37315
rect 31861 37281 31895 37315
rect 15577 37213 15611 37247
rect 16221 37213 16255 37247
rect 16405 37213 16439 37247
rect 17049 37213 17083 37247
rect 17233 37213 17267 37247
rect 20637 37213 20671 37247
rect 20913 37213 20947 37247
rect 22385 37213 22419 37247
rect 22478 37213 22512 37247
rect 22753 37213 22787 37247
rect 22850 37213 22884 37247
rect 23673 37213 23707 37247
rect 24777 37213 24811 37247
rect 24869 37213 24903 37247
rect 25053 37213 25087 37247
rect 25145 37213 25179 37247
rect 25789 37213 25823 37247
rect 25973 37213 26007 37247
rect 26525 37213 26559 37247
rect 26709 37213 26743 37247
rect 27629 37213 27663 37247
rect 27721 37213 27755 37247
rect 27905 37213 27939 37247
rect 28549 37213 28583 37247
rect 30849 37213 30883 37247
rect 31585 37213 31619 37247
rect 31769 37213 31803 37247
rect 32045 37213 32079 37247
rect 32505 37213 32539 37247
rect 32689 37213 32723 37247
rect 32873 37213 32907 37247
rect 34897 37213 34931 37247
rect 35081 37213 35115 37247
rect 15393 37145 15427 37179
rect 21925 37145 21959 37179
rect 22661 37145 22695 37179
rect 26617 37145 26651 37179
rect 28733 37145 28767 37179
rect 28917 37145 28951 37179
rect 33793 37145 33827 37179
rect 16497 37077 16531 37111
rect 17233 37077 17267 37111
rect 17785 37077 17819 37111
rect 19717 37077 19751 37111
rect 20453 37077 20487 37111
rect 20821 37077 20855 37111
rect 23029 37077 23063 37111
rect 24041 37077 24075 37111
rect 25881 37077 25915 37111
rect 30113 37077 30147 37111
rect 30395 37077 30429 37111
rect 30481 37077 30515 37111
rect 30573 37077 30607 37111
rect 31401 37077 31435 37111
rect 33993 37077 34027 37111
rect 34161 37077 34195 37111
rect 34989 37077 35023 37111
rect 36185 37077 36219 37111
rect 24133 36873 24167 36907
rect 31677 36873 31711 36907
rect 33885 36873 33919 36907
rect 16313 36805 16347 36839
rect 22109 36805 22143 36839
rect 22293 36805 22327 36839
rect 27629 36805 27663 36839
rect 29101 36805 29135 36839
rect 15117 36737 15151 36771
rect 16129 36737 16163 36771
rect 17509 36737 17543 36771
rect 18797 36737 18831 36771
rect 19441 36737 19475 36771
rect 19625 36737 19659 36771
rect 20361 36737 20395 36771
rect 20453 36737 20487 36771
rect 20637 36737 20671 36771
rect 20729 36737 20763 36771
rect 22385 36737 22419 36771
rect 22482 36737 22516 36771
rect 23949 36737 23983 36771
rect 24225 36737 24259 36771
rect 25329 36737 25363 36771
rect 25513 36737 25547 36771
rect 25789 36737 25823 36771
rect 26249 36737 26283 36771
rect 27905 36737 27939 36771
rect 28365 36737 28399 36771
rect 28549 36737 28583 36771
rect 29837 36737 29871 36771
rect 29929 36737 29963 36771
rect 30665 36737 30699 36771
rect 30849 36737 30883 36771
rect 31493 36737 31527 36771
rect 32505 36737 32539 36771
rect 32689 36737 32723 36771
rect 32781 36737 32815 36771
rect 33793 36737 33827 36771
rect 34069 36737 34103 36771
rect 34989 36737 35023 36771
rect 15209 36669 15243 36703
rect 15485 36669 15519 36703
rect 16865 36669 16899 36703
rect 17785 36669 17819 36703
rect 18889 36669 18923 36703
rect 19533 36669 19567 36703
rect 22201 36669 22235 36703
rect 23305 36669 23339 36703
rect 25605 36669 25639 36703
rect 30021 36669 30055 36703
rect 30113 36669 30147 36703
rect 31309 36669 31343 36703
rect 34621 36669 34655 36703
rect 36369 36669 36403 36703
rect 18429 36601 18463 36635
rect 25421 36601 25455 36635
rect 32321 36601 32355 36635
rect 33241 36601 33275 36635
rect 34069 36601 34103 36635
rect 15945 36533 15979 36567
rect 20913 36533 20947 36567
rect 23765 36533 23799 36567
rect 25145 36533 25179 36567
rect 26433 36533 26467 36567
rect 28457 36533 28491 36567
rect 29653 36533 29687 36567
rect 30757 36533 30791 36567
rect 17509 36329 17543 36363
rect 18429 36329 18463 36363
rect 18659 36329 18693 36363
rect 21189 36329 21223 36363
rect 27629 36329 27663 36363
rect 31125 36329 31159 36363
rect 31769 36329 31803 36363
rect 20361 36261 20395 36295
rect 27077 36261 27111 36295
rect 33609 36261 33643 36295
rect 17693 36193 17727 36227
rect 20637 36193 20671 36227
rect 21557 36193 21591 36227
rect 22661 36193 22695 36227
rect 22753 36193 22787 36227
rect 24777 36193 24811 36227
rect 25605 36193 25639 36227
rect 27813 36193 27847 36227
rect 30021 36193 30055 36227
rect 31309 36193 31343 36227
rect 32689 36193 32723 36227
rect 17233 36125 17267 36159
rect 18337 36125 18371 36159
rect 18521 36125 18555 36159
rect 18797 36125 18831 36159
rect 19441 36125 19475 36159
rect 19625 36125 19659 36159
rect 20269 36125 20303 36159
rect 20545 36125 20579 36159
rect 21373 36125 21407 36159
rect 22569 36125 22603 36159
rect 22845 36125 22879 36159
rect 24869 36125 24903 36159
rect 24961 36125 24995 36159
rect 25053 36125 25087 36159
rect 25973 36125 26007 36159
rect 26801 36125 26835 36159
rect 26893 36125 26927 36159
rect 27537 36125 27571 36159
rect 29101 36125 29135 36159
rect 29929 36125 29963 36159
rect 31033 36125 31067 36159
rect 32781 36125 32815 36159
rect 33425 36125 33459 36159
rect 34161 36125 34195 36159
rect 34345 36125 34379 36159
rect 34897 36125 34931 36159
rect 35081 36125 35115 36159
rect 35173 36125 35207 36159
rect 35265 36125 35299 36159
rect 36553 36125 36587 36159
rect 23489 36057 23523 36091
rect 23857 36057 23891 36091
rect 25789 36057 25823 36091
rect 27077 36057 27111 36091
rect 28733 36057 28767 36091
rect 31309 36057 31343 36091
rect 19533 35989 19567 36023
rect 20729 35989 20763 36023
rect 22385 35989 22419 36023
rect 24593 35989 24627 36023
rect 27813 35989 27847 36023
rect 30297 35989 30331 36023
rect 32413 35989 32447 36023
rect 34161 35989 34195 36023
rect 35541 35989 35575 36023
rect 36093 35989 36127 36023
rect 14197 35785 14231 35819
rect 16865 35785 16899 35819
rect 20637 35785 20671 35819
rect 25053 35785 25087 35819
rect 28089 35785 28123 35819
rect 31769 35785 31803 35819
rect 32521 35785 32555 35819
rect 32689 35785 32723 35819
rect 33333 35785 33367 35819
rect 34345 35785 34379 35819
rect 14749 35717 14783 35751
rect 21465 35717 21499 35751
rect 22845 35717 22879 35751
rect 22937 35717 22971 35751
rect 24225 35717 24259 35751
rect 25421 35717 25455 35751
rect 27169 35717 27203 35751
rect 27353 35717 27387 35751
rect 30113 35717 30147 35751
rect 32321 35717 32355 35751
rect 33977 35717 34011 35751
rect 14105 35649 14139 35683
rect 14289 35649 14323 35683
rect 14933 35649 14967 35683
rect 15025 35649 15059 35683
rect 15577 35649 15611 35683
rect 15761 35649 15795 35683
rect 15853 35649 15887 35683
rect 15945 35649 15979 35683
rect 17233 35649 17267 35683
rect 19625 35649 19659 35683
rect 20269 35649 20303 35683
rect 20453 35649 20487 35683
rect 22569 35649 22603 35683
rect 22717 35649 22751 35683
rect 23034 35649 23068 35683
rect 24409 35649 24443 35683
rect 24593 35649 24627 35683
rect 25237 35649 25271 35683
rect 25329 35649 25363 35683
rect 25605 35649 25639 35683
rect 26433 35649 26467 35683
rect 26617 35649 26651 35683
rect 27997 35649 28031 35683
rect 28181 35649 28215 35683
rect 29009 35649 29043 35683
rect 29193 35649 29227 35683
rect 29929 35649 29963 35683
rect 30757 35649 30791 35683
rect 31125 35649 31159 35683
rect 33149 35649 33183 35683
rect 34161 35649 34195 35683
rect 34805 35649 34839 35683
rect 35173 35649 35207 35683
rect 17141 35581 17175 35615
rect 19349 35581 19383 35615
rect 20177 35581 20211 35615
rect 26525 35581 26559 35615
rect 28733 35581 28767 35615
rect 29561 35581 29595 35615
rect 36553 35581 36587 35615
rect 14749 35513 14783 35547
rect 19073 35513 19107 35547
rect 23765 35513 23799 35547
rect 18613 35445 18647 35479
rect 19441 35445 19475 35479
rect 23213 35445 23247 35479
rect 27537 35445 27571 35479
rect 30573 35445 30607 35479
rect 31033 35445 31067 35479
rect 32505 35445 32539 35479
rect 14565 35241 14599 35275
rect 14749 35241 14783 35275
rect 19533 35241 19567 35275
rect 25605 35241 25639 35275
rect 30849 35241 30883 35275
rect 17693 35173 17727 35207
rect 15669 35105 15703 35139
rect 16865 35105 16899 35139
rect 18153 35105 18187 35139
rect 29837 35105 29871 35139
rect 30021 35105 30055 35139
rect 30113 35105 30147 35139
rect 31861 35105 31895 35139
rect 33241 35105 33275 35139
rect 35817 35105 35851 35139
rect 1869 35037 1903 35071
rect 15577 35037 15611 35071
rect 17049 35037 17083 35071
rect 17233 35037 17267 35071
rect 18061 35037 18095 35071
rect 19441 35037 19475 35071
rect 19625 35037 19659 35071
rect 20545 35037 20579 35071
rect 20729 35037 20763 35071
rect 20821 35037 20855 35071
rect 20913 35037 20947 35071
rect 22661 35037 22695 35071
rect 22845 35037 22879 35071
rect 23029 35037 23063 35071
rect 24777 35037 24811 35071
rect 25053 35037 25087 35071
rect 26249 35037 26283 35071
rect 26617 35037 26651 35071
rect 27077 35037 27111 35071
rect 28365 35037 28399 35071
rect 28549 35037 28583 35071
rect 29929 35037 29963 35071
rect 31585 35037 31619 35071
rect 31769 35037 31803 35071
rect 31953 35037 31987 35071
rect 32137 35037 32171 35071
rect 33149 35037 33183 35071
rect 33333 35037 33367 35071
rect 33425 35037 33459 35071
rect 33977 35037 34011 35071
rect 34161 35037 34195 35071
rect 36093 35037 36127 35071
rect 14933 34969 14967 35003
rect 15393 34969 15427 35003
rect 22753 34969 22787 35003
rect 24961 34969 24995 35003
rect 26341 34969 26375 35003
rect 26433 34969 26467 35003
rect 28089 34969 28123 35003
rect 1685 34901 1719 34935
rect 2329 34901 2363 34935
rect 14733 34901 14767 34935
rect 16037 34901 16071 34935
rect 21189 34901 21223 34935
rect 21649 34901 21683 34935
rect 22477 34901 22511 34935
rect 24593 34901 24627 34935
rect 26065 34901 26099 34935
rect 27261 34901 27295 34935
rect 30297 34901 30331 34935
rect 31401 34901 31435 34935
rect 32965 34901 32999 34935
rect 34069 34901 34103 34935
rect 36645 34901 36679 34935
rect 15485 34697 15519 34731
rect 18245 34697 18279 34731
rect 22937 34697 22971 34731
rect 24869 34697 24903 34731
rect 29101 34697 29135 34731
rect 58265 34697 58299 34731
rect 18613 34629 18647 34663
rect 19809 34629 19843 34663
rect 26617 34629 26651 34663
rect 27169 34629 27203 34663
rect 27905 34629 27939 34663
rect 33057 34629 33091 34663
rect 34529 34629 34563 34663
rect 18429 34561 18463 34595
rect 21005 34561 21039 34595
rect 22477 34561 22511 34595
rect 23397 34561 23431 34595
rect 23581 34561 23615 34595
rect 23673 34561 23707 34595
rect 24777 34561 24811 34595
rect 24961 34561 24995 34595
rect 25605 34561 25639 34595
rect 27721 34561 27755 34595
rect 27997 34561 28031 34595
rect 28089 34561 28123 34595
rect 28825 34561 28859 34595
rect 29653 34561 29687 34595
rect 29745 34561 29779 34595
rect 30021 34561 30055 34595
rect 30849 34561 30883 34595
rect 31125 34561 31159 34595
rect 32321 34561 32355 34595
rect 33885 34561 33919 34595
rect 35541 34561 35575 34595
rect 35725 34561 35759 34595
rect 36553 34561 36587 34595
rect 37657 34561 37691 34595
rect 58081 34561 58115 34595
rect 15025 34493 15059 34527
rect 15117 34493 15151 34527
rect 19165 34493 19199 34527
rect 21097 34493 21131 34527
rect 22293 34493 22327 34527
rect 22569 34493 22603 34527
rect 25789 34493 25823 34527
rect 29837 34493 29871 34527
rect 30665 34493 30699 34527
rect 30941 34493 30975 34527
rect 31033 34493 31067 34527
rect 31677 34493 31711 34527
rect 32413 34493 32447 34527
rect 33977 34493 34011 34527
rect 36645 34493 36679 34527
rect 36921 34493 36955 34527
rect 37565 34493 37599 34527
rect 57437 34493 57471 34527
rect 21373 34425 21407 34459
rect 33517 34425 33551 34459
rect 38025 34425 38059 34459
rect 14841 34357 14875 34391
rect 20361 34357 20395 34391
rect 28273 34357 28307 34391
rect 30021 34357 30055 34391
rect 35633 34357 35667 34391
rect 15669 34153 15703 34187
rect 20913 34153 20947 34187
rect 23581 34153 23615 34187
rect 30665 34153 30699 34187
rect 33793 34153 33827 34187
rect 17417 34085 17451 34119
rect 23397 34085 23431 34119
rect 29193 34085 29227 34119
rect 32597 34085 32631 34119
rect 33425 34085 33459 34119
rect 38945 34085 38979 34119
rect 15393 34017 15427 34051
rect 18429 34017 18463 34051
rect 20085 34017 20119 34051
rect 20361 34017 20395 34051
rect 20821 34017 20855 34051
rect 22293 34017 22327 34051
rect 24777 34017 24811 34051
rect 25237 34017 25271 34051
rect 25789 34017 25823 34051
rect 27537 34017 27571 34051
rect 27721 34017 27755 34051
rect 28641 34017 28675 34051
rect 30021 34017 30055 34051
rect 31401 34017 31435 34051
rect 31585 34017 31619 34051
rect 32413 34017 32447 34051
rect 33517 34017 33551 34051
rect 34989 34017 35023 34051
rect 35449 34017 35483 34051
rect 15301 33949 15335 33983
rect 17601 33949 17635 33983
rect 17693 33949 17727 33983
rect 18337 33949 18371 33983
rect 18521 33949 18555 33983
rect 18613 33949 18647 33983
rect 19993 33949 20027 33983
rect 21097 33949 21131 33983
rect 21741 33949 21775 33983
rect 22753 33949 22787 33983
rect 24869 33949 24903 33983
rect 26157 33949 26191 33983
rect 26249 33949 26283 33983
rect 27445 33949 27479 33983
rect 27629 33949 27663 33983
rect 31309 33949 31343 33983
rect 31493 33949 31527 33983
rect 32689 33949 32723 33983
rect 33149 33949 33183 33983
rect 33333 33949 33367 33983
rect 33609 33949 33643 33983
rect 35081 33949 35115 33983
rect 36093 33949 36127 33983
rect 36277 33949 36311 33983
rect 38669 33949 38703 33983
rect 38945 33949 38979 33983
rect 17417 33881 17451 33915
rect 22109 33881 22143 33915
rect 23765 33881 23799 33915
rect 26433 33881 26467 33915
rect 28825 33881 28859 33915
rect 30297 33881 30331 33915
rect 32413 33881 32447 33915
rect 18153 33813 18187 33847
rect 21281 33813 21315 33847
rect 21925 33813 21959 33847
rect 22017 33813 22051 33847
rect 23565 33813 23599 33847
rect 24593 33813 24627 33847
rect 24961 33813 24995 33847
rect 25145 33813 25179 33847
rect 25881 33813 25915 33847
rect 26065 33813 26099 33847
rect 27905 33813 27939 33847
rect 28733 33813 28767 33847
rect 30205 33813 30239 33847
rect 31125 33813 31159 33847
rect 34253 33813 34287 33847
rect 35909 33813 35943 33847
rect 38761 33813 38795 33847
rect 19533 33609 19567 33643
rect 19717 33609 19751 33643
rect 22201 33609 22235 33643
rect 23029 33609 23063 33643
rect 25145 33609 25179 33643
rect 27261 33609 27295 33643
rect 28181 33609 28215 33643
rect 30389 33609 30423 33643
rect 34805 33609 34839 33643
rect 36277 33609 36311 33643
rect 37841 33609 37875 33643
rect 38393 33609 38427 33643
rect 24041 33541 24075 33575
rect 24777 33541 24811 33575
rect 26433 33541 26467 33575
rect 27445 33541 27479 33575
rect 33609 33541 33643 33575
rect 33793 33541 33827 33575
rect 25007 33507 25041 33541
rect 15025 33473 15059 33507
rect 15853 33473 15887 33507
rect 16037 33473 16071 33507
rect 17969 33473 18003 33507
rect 19349 33473 19383 33507
rect 19625 33473 19659 33507
rect 20821 33473 20855 33507
rect 21005 33473 21039 33507
rect 22845 33473 22879 33507
rect 23305 33473 23339 33507
rect 23765 33473 23799 33507
rect 23857 33473 23891 33507
rect 25605 33473 25639 33507
rect 25789 33473 25823 33507
rect 26617 33473 26651 33507
rect 27169 33473 27203 33507
rect 30297 33473 30331 33507
rect 31033 33473 31067 33507
rect 31217 33473 31251 33507
rect 31677 33473 31711 33507
rect 32321 33473 32355 33507
rect 32505 33473 32539 33507
rect 32597 33473 32631 33507
rect 32689 33473 32723 33507
rect 34253 33473 34287 33507
rect 35633 33473 35667 33507
rect 35817 33473 35851 33507
rect 36645 33473 36679 33507
rect 37473 33473 37507 33507
rect 37657 33473 37691 33507
rect 38301 33473 38335 33507
rect 38577 33473 38611 33507
rect 39681 33473 39715 33507
rect 40049 33473 40083 33507
rect 15117 33405 15151 33439
rect 15393 33405 15427 33439
rect 17877 33405 17911 33439
rect 20637 33405 20671 33439
rect 20913 33405 20947 33439
rect 21097 33405 21131 33439
rect 22661 33405 22695 33439
rect 22937 33405 22971 33439
rect 23213 33405 23247 33439
rect 33425 33405 33459 33439
rect 36737 33405 36771 33439
rect 40693 33405 40727 33439
rect 25697 33337 25731 33371
rect 27445 33337 27479 33371
rect 29193 33337 29227 33371
rect 16037 33269 16071 33303
rect 17601 33269 17635 33303
rect 19901 33269 19935 33303
rect 24041 33269 24075 33303
rect 24983 33269 25017 33303
rect 26249 33269 26283 33303
rect 31217 33269 31251 33303
rect 32965 33269 32999 33303
rect 35725 33269 35759 33303
rect 36921 33269 36955 33303
rect 38761 33269 38795 33303
rect 22109 33065 22143 33099
rect 31309 33065 31343 33099
rect 31953 33065 31987 33099
rect 32321 33065 32355 33099
rect 33241 33065 33275 33099
rect 34069 33065 34103 33099
rect 38853 33065 38887 33099
rect 40417 33065 40451 33099
rect 15945 32997 15979 33031
rect 16773 32997 16807 33031
rect 27813 32997 27847 33031
rect 29837 32997 29871 33031
rect 15669 32929 15703 32963
rect 17233 32929 17267 32963
rect 21005 32929 21039 32963
rect 22201 32929 22235 32963
rect 26248 32929 26282 32963
rect 26441 32929 26475 32963
rect 27353 32929 27387 32963
rect 28549 32929 28583 32963
rect 29009 32929 29043 32963
rect 32229 32929 32263 32963
rect 36553 32929 36587 32963
rect 37013 32929 37047 32963
rect 17141 32861 17175 32895
rect 20821 32861 20855 32895
rect 21281 32861 21315 32895
rect 21925 32861 21959 32895
rect 23029 32861 23063 32895
rect 23305 32861 23339 32895
rect 24593 32861 24627 32895
rect 24869 32861 24903 32895
rect 26157 32861 26191 32895
rect 26340 32861 26374 32895
rect 27445 32861 27479 32895
rect 28641 32861 28675 32895
rect 29745 32861 29779 32895
rect 29929 32861 29963 32895
rect 31861 32861 31895 32895
rect 32137 32861 32171 32895
rect 33241 32861 33275 32895
rect 33333 32861 33367 32895
rect 34897 32861 34931 32895
rect 35817 32861 35851 32895
rect 36001 32861 36035 32895
rect 36645 32861 36679 32895
rect 36829 32861 36863 32895
rect 37565 32861 37599 32895
rect 37657 32861 37691 32895
rect 40233 32861 40267 32895
rect 18889 32793 18923 32827
rect 19533 32793 19567 32827
rect 21189 32793 21223 32827
rect 23213 32793 23247 32827
rect 25053 32793 25087 32827
rect 38669 32793 38703 32827
rect 38885 32793 38919 32827
rect 40049 32793 40083 32827
rect 16129 32725 16163 32759
rect 19809 32725 19843 32759
rect 21741 32725 21775 32759
rect 22845 32725 22879 32759
rect 23765 32725 23799 32759
rect 24685 32725 24719 32759
rect 26617 32725 26651 32759
rect 33609 32725 33643 32759
rect 35817 32725 35851 32759
rect 37841 32725 37875 32759
rect 39037 32725 39071 32759
rect 25973 32521 26007 32555
rect 30481 32521 30515 32555
rect 31769 32521 31803 32555
rect 35265 32521 35299 32555
rect 36093 32521 36127 32555
rect 39589 32521 39623 32555
rect 20545 32453 20579 32487
rect 24869 32453 24903 32487
rect 25891 32453 25925 32487
rect 27261 32453 27295 32487
rect 27997 32453 28031 32487
rect 32781 32453 32815 32487
rect 36369 32453 36403 32487
rect 18429 32385 18463 32419
rect 19625 32385 19659 32419
rect 20453 32385 20487 32419
rect 20637 32385 20671 32419
rect 23397 32385 23431 32419
rect 23489 32385 23523 32419
rect 23673 32385 23707 32419
rect 24593 32385 24627 32419
rect 24961 32385 24995 32419
rect 25789 32385 25823 32419
rect 26157 32385 26191 32419
rect 27445 32385 27479 32419
rect 27537 32385 27571 32419
rect 28825 32385 28859 32419
rect 29009 32385 29043 32419
rect 29469 32385 29503 32419
rect 31309 32385 31343 32419
rect 32965 32385 32999 32419
rect 33057 32385 33091 32419
rect 33609 32385 33643 32419
rect 33701 32385 33735 32419
rect 33977 32385 34011 32419
rect 34345 32385 34379 32419
rect 35173 32385 35207 32419
rect 35449 32385 35483 32419
rect 36093 32385 36127 32419
rect 36185 32385 36219 32419
rect 37657 32385 37691 32419
rect 37933 32385 37967 32419
rect 38577 32385 38611 32419
rect 38853 32385 38887 32419
rect 39405 32385 39439 32419
rect 39589 32385 39623 32419
rect 15853 32317 15887 32351
rect 18245 32317 18279 32351
rect 19717 32317 19751 32351
rect 23581 32317 23615 32351
rect 24501 32317 24535 32351
rect 30205 32317 30239 32351
rect 30389 32317 30423 32351
rect 32781 32317 32815 32351
rect 34161 32317 34195 32351
rect 38669 32317 38703 32351
rect 38761 32317 38795 32351
rect 15485 32249 15519 32283
rect 25605 32249 25639 32283
rect 28825 32249 28859 32283
rect 30849 32249 30883 32283
rect 15393 32181 15427 32215
rect 18613 32181 18647 32215
rect 19901 32181 19935 32215
rect 21373 32181 21407 32215
rect 23213 32181 23247 32215
rect 27261 32181 27295 32215
rect 31401 32181 31435 32215
rect 35633 32181 35667 32215
rect 37473 32181 37507 32215
rect 37841 32181 37875 32215
rect 38393 32181 38427 32215
rect 22017 31977 22051 32011
rect 24593 31977 24627 32011
rect 24961 31977 24995 32011
rect 26985 31977 27019 32011
rect 28365 31977 28399 32011
rect 30389 31977 30423 32011
rect 36093 31977 36127 32011
rect 37657 31977 37691 32011
rect 26893 31909 26927 31943
rect 31677 31909 31711 31943
rect 16681 31841 16715 31875
rect 16957 31841 16991 31875
rect 18613 31841 18647 31875
rect 19993 31841 20027 31875
rect 20453 31841 20487 31875
rect 23121 31841 23155 31875
rect 27537 31841 27571 31875
rect 31217 31841 31251 31875
rect 33793 31841 33827 31875
rect 33885 31841 33919 31875
rect 34897 31841 34931 31875
rect 35541 31841 35575 31875
rect 36461 31841 36495 31875
rect 15301 31773 15335 31807
rect 15761 31773 15795 31807
rect 17049 31773 17083 31807
rect 18061 31773 18095 31807
rect 18245 31773 18279 31807
rect 20085 31773 20119 31807
rect 20913 31773 20947 31807
rect 21097 31773 21131 31807
rect 21281 31773 21315 31807
rect 21741 31773 21775 31807
rect 22017 31773 22051 31807
rect 23029 31773 23063 31807
rect 24777 31773 24811 31807
rect 25053 31773 25087 31807
rect 25513 31773 25547 31807
rect 25697 31773 25731 31807
rect 26985 31773 27019 31807
rect 30481 31773 30515 31807
rect 31309 31773 31343 31807
rect 32505 31773 32539 31807
rect 32689 31773 32723 31807
rect 33609 31773 33643 31807
rect 33701 31773 33735 31807
rect 35449 31773 35483 31807
rect 35633 31773 35667 31807
rect 36277 31773 36311 31807
rect 37289 31773 37323 31807
rect 37473 31773 37507 31807
rect 21833 31705 21867 31739
rect 26249 31705 26283 31739
rect 26709 31705 26743 31739
rect 27813 31705 27847 31739
rect 18521 31637 18555 31671
rect 22661 31637 22695 31671
rect 25697 31637 25731 31671
rect 32597 31637 32631 31671
rect 34069 31637 34103 31671
rect 15577 31433 15611 31467
rect 22109 31433 22143 31467
rect 24777 31433 24811 31467
rect 27261 31433 27295 31467
rect 28089 31433 28123 31467
rect 32689 31433 32723 31467
rect 34361 31433 34395 31467
rect 34529 31433 34563 31467
rect 15117 31365 15151 31399
rect 27429 31365 27463 31399
rect 27629 31365 27663 31399
rect 30849 31365 30883 31399
rect 33149 31365 33183 31399
rect 33333 31365 33367 31399
rect 34161 31365 34195 31399
rect 36737 31365 36771 31399
rect 14841 31297 14875 31331
rect 14933 31297 14967 31331
rect 15761 31297 15795 31331
rect 15945 31297 15979 31331
rect 16037 31297 16071 31331
rect 18061 31297 18095 31331
rect 22017 31297 22051 31331
rect 22293 31297 22327 31331
rect 24593 31297 24627 31331
rect 24869 31297 24903 31331
rect 25881 31297 25915 31331
rect 26065 31297 26099 31331
rect 28457 31297 28491 31331
rect 29193 31297 29227 31331
rect 31033 31297 31067 31331
rect 32505 31297 32539 31331
rect 35357 31297 35391 31331
rect 36553 31297 36587 31331
rect 17693 31229 17727 31263
rect 18153 31229 18187 31263
rect 25789 31229 25823 31263
rect 25973 31229 26007 31263
rect 26249 31229 26283 31263
rect 28549 31229 28583 31263
rect 30113 31229 30147 31263
rect 31217 31229 31251 31263
rect 32321 31229 32355 31263
rect 35173 31229 35207 31263
rect 15117 31161 15151 31195
rect 22477 31093 22511 31127
rect 24593 31093 24627 31127
rect 27445 31093 27479 31127
rect 33517 31093 33551 31127
rect 34345 31093 34379 31127
rect 35541 31093 35575 31127
rect 36921 31093 36955 31127
rect 15853 30889 15887 30923
rect 16037 30889 16071 30923
rect 20545 30889 20579 30923
rect 25973 30889 26007 30923
rect 27445 30889 27479 30923
rect 31493 30889 31527 30923
rect 34161 30889 34195 30923
rect 34345 30889 34379 30923
rect 36185 30889 36219 30923
rect 22109 30821 22143 30855
rect 24593 30821 24627 30855
rect 32781 30821 32815 30855
rect 16129 30753 16163 30787
rect 17969 30753 18003 30787
rect 21281 30753 21315 30787
rect 30665 30753 30699 30787
rect 34989 30753 35023 30787
rect 37289 30753 37323 30787
rect 38025 30753 38059 30787
rect 16221 30685 16255 30719
rect 18245 30685 18279 30719
rect 18889 30685 18923 30719
rect 19717 30685 19751 30719
rect 21833 30685 21867 30719
rect 22569 30685 22603 30719
rect 22753 30685 22787 30719
rect 23857 30685 23891 30719
rect 24041 30685 24075 30719
rect 24777 30685 24811 30719
rect 24869 30685 24903 30719
rect 25605 30685 25639 30719
rect 26433 30685 26467 30719
rect 27445 30685 27479 30719
rect 27537 30685 27571 30719
rect 28273 30685 28307 30719
rect 28457 30685 28491 30719
rect 30573 30685 30607 30719
rect 31401 30685 31435 30719
rect 31585 30685 31619 30719
rect 32689 30685 32723 30719
rect 32965 30685 32999 30719
rect 33885 30685 33919 30719
rect 34897 30685 34931 30719
rect 35081 30685 35115 30719
rect 35633 30685 35667 30719
rect 35725 30685 35759 30719
rect 35909 30685 35943 30719
rect 36001 30685 36035 30719
rect 37197 30685 37231 30719
rect 19901 30617 19935 30651
rect 20529 30617 20563 30651
rect 20729 30617 20763 30651
rect 22109 30617 22143 30651
rect 23949 30617 23983 30651
rect 24593 30617 24627 30651
rect 25789 30617 25823 30651
rect 19533 30549 19567 30583
rect 20361 30549 20395 30583
rect 21925 30549 21959 30583
rect 22569 30549 22603 30583
rect 26617 30549 26651 30583
rect 27813 30549 27847 30583
rect 28365 30549 28399 30583
rect 29009 30549 29043 30583
rect 30941 30549 30975 30583
rect 17969 30345 18003 30379
rect 23857 30345 23891 30379
rect 26249 30345 26283 30379
rect 26617 30345 26651 30379
rect 27629 30345 27663 30379
rect 20177 30277 20211 30311
rect 20361 30277 20395 30311
rect 29377 30277 29411 30311
rect 33977 30277 34011 30311
rect 34193 30277 34227 30311
rect 34897 30277 34931 30311
rect 35725 30277 35759 30311
rect 36737 30277 36771 30311
rect 18153 30209 18187 30243
rect 18429 30209 18463 30243
rect 18613 30209 18647 30243
rect 19717 30209 19751 30243
rect 20453 30209 20487 30243
rect 20913 30209 20947 30243
rect 21005 30209 21039 30243
rect 22753 30209 22787 30243
rect 24041 30209 24075 30243
rect 24685 30209 24719 30243
rect 24869 30209 24903 30243
rect 27537 30209 27571 30243
rect 28365 30209 28399 30243
rect 28457 30209 28491 30243
rect 28641 30209 28675 30243
rect 28733 30209 28767 30243
rect 31585 30209 31619 30243
rect 32781 30209 32815 30243
rect 34805 30209 34839 30243
rect 34989 30209 35023 30243
rect 35909 30209 35943 30243
rect 36093 30209 36127 30243
rect 36185 30209 36219 30243
rect 36645 30209 36679 30243
rect 36829 30209 36863 30243
rect 21189 30141 21223 30175
rect 22661 30141 22695 30175
rect 25973 30141 26007 30175
rect 26157 30141 26191 30175
rect 27721 30141 27755 30175
rect 31677 30141 31711 30175
rect 33241 30141 33275 30175
rect 20177 30073 20211 30107
rect 27169 30073 27203 30107
rect 31217 30073 31251 30107
rect 21097 30005 21131 30039
rect 22477 30005 22511 30039
rect 25053 30005 25087 30039
rect 28917 30005 28951 30039
rect 32873 30005 32907 30039
rect 34161 30005 34195 30039
rect 34345 30005 34379 30039
rect 20821 29801 20855 29835
rect 22569 29801 22603 29835
rect 27629 29801 27663 29835
rect 28641 29801 28675 29835
rect 19717 29733 19751 29767
rect 26157 29733 26191 29767
rect 32965 29733 32999 29767
rect 20729 29665 20763 29699
rect 21833 29665 21867 29699
rect 24869 29665 24903 29699
rect 25145 29665 25179 29699
rect 26617 29665 26651 29699
rect 19625 29597 19659 29631
rect 19809 29597 19843 29631
rect 19901 29597 19935 29631
rect 20821 29597 20855 29631
rect 21741 29597 21775 29631
rect 22385 29597 22419 29631
rect 22569 29597 22603 29631
rect 24777 29597 24811 29631
rect 25973 29597 26007 29631
rect 26893 29597 26927 29631
rect 28549 29597 28583 29631
rect 29837 29597 29871 29631
rect 32229 29597 32263 29631
rect 32689 29597 32723 29631
rect 32965 29597 32999 29631
rect 33517 29597 33551 29631
rect 30849 29529 30883 29563
rect 34161 29529 34195 29563
rect 19441 29461 19475 29495
rect 20453 29461 20487 29495
rect 21373 29461 21407 29495
rect 23857 29461 23891 29495
rect 31309 29461 31343 29495
rect 32781 29461 32815 29495
rect 33517 29461 33551 29495
rect 2421 29257 2455 29291
rect 27169 29257 27203 29291
rect 28457 29257 28491 29291
rect 29009 29257 29043 29291
rect 30665 29257 30699 29291
rect 31769 29257 31803 29291
rect 16957 29189 16991 29223
rect 20913 29189 20947 29223
rect 30205 29189 30239 29223
rect 30757 29189 30791 29223
rect 30941 29189 30975 29223
rect 31401 29189 31435 29223
rect 31601 29189 31635 29223
rect 34069 29189 34103 29223
rect 1869 29121 1903 29155
rect 18245 29121 18279 29155
rect 19165 29121 19199 29155
rect 19349 29121 19383 29155
rect 19993 29121 20027 29155
rect 20085 29121 20119 29155
rect 20637 29121 20671 29155
rect 23581 29121 23615 29155
rect 23765 29121 23799 29155
rect 24935 29121 24969 29155
rect 25031 29121 25065 29155
rect 25237 29121 25271 29155
rect 26065 29121 26099 29155
rect 26617 29121 26651 29155
rect 27353 29121 27387 29155
rect 28273 29121 28307 29155
rect 28549 29121 28583 29155
rect 29653 29121 29687 29155
rect 29837 29121 29871 29155
rect 30665 29121 30699 29155
rect 32504 29121 32538 29155
rect 32689 29121 32723 29155
rect 58081 29121 58115 29155
rect 17417 29053 17451 29087
rect 18153 29053 18187 29087
rect 20729 29053 20763 29087
rect 24317 29053 24351 29087
rect 25145 29053 25179 29087
rect 27537 29053 27571 29087
rect 32413 29053 32447 29087
rect 32597 29053 32631 29087
rect 33793 29053 33827 29087
rect 35817 29053 35851 29087
rect 57437 29053 57471 29087
rect 1685 28985 1719 29019
rect 17325 28985 17359 29019
rect 19257 28985 19291 29019
rect 19809 28985 19843 29019
rect 20637 28985 20671 29019
rect 32873 28985 32907 29019
rect 58265 28985 58299 29019
rect 17877 28917 17911 28951
rect 23673 28917 23707 28951
rect 24777 28917 24811 28951
rect 30113 28917 30147 28951
rect 31585 28917 31619 28951
rect 19625 28713 19659 28747
rect 20177 28713 20211 28747
rect 17877 28645 17911 28679
rect 25513 28645 25547 28679
rect 18061 28577 18095 28611
rect 19901 28577 19935 28611
rect 20637 28577 20671 28611
rect 23121 28577 23155 28611
rect 23581 28577 23615 28611
rect 26249 28577 26283 28611
rect 28273 28577 28307 28611
rect 29929 28577 29963 28611
rect 18613 28509 18647 28543
rect 18889 28509 18923 28543
rect 19993 28509 20027 28543
rect 22293 28509 22327 28543
rect 22477 28509 22511 28543
rect 23489 28509 23523 28543
rect 26801 28509 26835 28543
rect 27629 28509 27663 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 28825 28509 28859 28543
rect 29009 28509 29043 28543
rect 30941 28509 30975 28543
rect 32505 28509 32539 28543
rect 32781 28509 32815 28543
rect 35265 28509 35299 28543
rect 17601 28441 17635 28475
rect 19533 28441 19567 28475
rect 20821 28441 20855 28475
rect 21005 28441 21039 28475
rect 25145 28441 25179 28475
rect 35541 28441 35575 28475
rect 37289 28441 37323 28475
rect 18613 28373 18647 28407
rect 22385 28373 22419 28407
rect 25605 28373 25639 28407
rect 26985 28373 27019 28407
rect 29009 28373 29043 28407
rect 24869 28169 24903 28203
rect 29653 28169 29687 28203
rect 18889 28101 18923 28135
rect 23305 28101 23339 28135
rect 27169 28101 27203 28135
rect 28917 28101 28951 28135
rect 31125 28101 31159 28135
rect 20085 28033 20119 28067
rect 20913 28033 20947 28067
rect 22293 28033 22327 28067
rect 23121 28033 23155 28067
rect 24409 28033 24443 28067
rect 25421 28033 25455 28067
rect 25605 28033 25639 28067
rect 33149 28033 33183 28067
rect 33609 28033 33643 28067
rect 34805 28033 34839 28067
rect 34989 28033 35023 28067
rect 35081 28033 35115 28067
rect 35173 28033 35207 28067
rect 35909 28033 35943 28067
rect 19257 27965 19291 27999
rect 19349 27965 19383 27999
rect 19533 27965 19567 27999
rect 21005 27965 21039 27999
rect 22201 27965 22235 27999
rect 22661 27965 22695 27999
rect 23489 27965 23523 27999
rect 25329 27965 25363 27999
rect 29193 27965 29227 27999
rect 31401 27965 31435 27999
rect 22017 27829 22051 27863
rect 24685 27829 24719 27863
rect 25789 27829 25823 27863
rect 35449 27829 35483 27863
rect 36461 27829 36495 27863
rect 28365 27625 28399 27659
rect 36166 27625 36200 27659
rect 26341 27557 26375 27591
rect 30757 27557 30791 27591
rect 22293 27489 22327 27523
rect 26893 27489 26927 27523
rect 29009 27489 29043 27523
rect 20637 27421 20671 27455
rect 22385 27421 22419 27455
rect 23213 27421 23247 27455
rect 23673 27421 23707 27455
rect 25605 27421 25639 27455
rect 27077 27421 27111 27455
rect 27261 27421 27295 27455
rect 27905 27421 27939 27455
rect 30665 27421 30699 27455
rect 30849 27421 30883 27455
rect 31309 27421 31343 27455
rect 34161 27421 34195 27455
rect 34345 27421 34379 27455
rect 35909 27421 35943 27455
rect 20821 27353 20855 27387
rect 21005 27353 21039 27387
rect 24593 27353 24627 27387
rect 35081 27353 35115 27387
rect 35265 27353 35299 27387
rect 37933 27353 37967 27387
rect 38393 27353 38427 27387
rect 22017 27285 22051 27319
rect 23857 27285 23891 27319
rect 27721 27285 27755 27319
rect 30113 27285 30147 27319
rect 31493 27285 31527 27319
rect 32597 27285 32631 27319
rect 33241 27285 33275 27319
rect 34253 27285 34287 27319
rect 34897 27285 34931 27319
rect 24685 27081 24719 27115
rect 30021 27081 30055 27115
rect 35357 27081 35391 27115
rect 37473 27081 37507 27115
rect 39497 27081 39531 27115
rect 23857 27013 23891 27047
rect 27445 27013 27479 27047
rect 31493 27013 31527 27047
rect 34069 27013 34103 27047
rect 21189 26945 21223 26979
rect 21373 26945 21407 26979
rect 31769 26945 31803 26979
rect 32873 26945 32907 26979
rect 33793 26945 33827 26979
rect 33977 26945 34011 26979
rect 34713 26945 34747 26979
rect 34897 26945 34931 26979
rect 34989 26945 35023 26979
rect 35081 26945 35115 26979
rect 36277 26945 36311 26979
rect 38485 26945 38519 26979
rect 20453 26877 20487 26911
rect 24133 26877 24167 26911
rect 27169 26877 27203 26911
rect 32689 26877 32723 26911
rect 38301 26877 38335 26911
rect 22385 26741 22419 26775
rect 28917 26741 28951 26775
rect 33057 26741 33091 26775
rect 36093 26741 36127 26775
rect 36829 26741 36863 26775
rect 38945 26741 38979 26775
rect 41889 26741 41923 26775
rect 42809 26741 42843 26775
rect 23673 26537 23707 26571
rect 30021 26537 30055 26571
rect 33425 26537 33459 26571
rect 34161 26537 34195 26571
rect 35265 26537 35299 26571
rect 29193 26469 29227 26503
rect 30113 26469 30147 26503
rect 31953 26469 31987 26503
rect 39405 26469 39439 26503
rect 24593 26401 24627 26435
rect 26617 26401 26651 26435
rect 27721 26401 27755 26435
rect 30481 26401 30515 26435
rect 35817 26401 35851 26435
rect 37841 26401 37875 26435
rect 40141 26401 40175 26435
rect 23949 26333 23983 26367
rect 27445 26333 27479 26367
rect 31033 26333 31067 26367
rect 33241 26333 33275 26367
rect 34069 26333 34103 26367
rect 34253 26333 34287 26367
rect 34897 26333 34931 26367
rect 39221 26333 39255 26367
rect 41153 26333 41187 26367
rect 42533 26333 42567 26367
rect 42993 26333 43027 26367
rect 24869 26265 24903 26299
rect 31401 26265 31435 26299
rect 32689 26265 32723 26299
rect 35081 26265 35115 26299
rect 36093 26265 36127 26299
rect 38301 26265 38335 26299
rect 38669 26265 38703 26299
rect 42257 26265 42291 26299
rect 43269 26265 43303 26299
rect 40601 26197 40635 26231
rect 24133 25993 24167 26027
rect 26617 25993 26651 26027
rect 31401 25993 31435 26027
rect 33149 25993 33183 26027
rect 35725 25993 35759 26027
rect 38301 25993 38335 26027
rect 41061 25993 41095 26027
rect 29469 25925 29503 25959
rect 34345 25925 34379 25959
rect 35357 25925 35391 25959
rect 36277 25925 36311 25959
rect 42625 25925 42659 25959
rect 26249 25857 26283 25891
rect 33609 25857 33643 25891
rect 33793 25857 33827 25891
rect 34253 25857 34287 25891
rect 34437 25857 34471 25891
rect 35173 25857 35207 25891
rect 35449 25857 35483 25891
rect 35541 25857 35575 25891
rect 36185 25857 36219 25891
rect 36369 25857 36403 25891
rect 39497 25857 39531 25891
rect 40141 25857 40175 25891
rect 41153 25857 41187 25891
rect 43453 25857 43487 25891
rect 43545 25857 43579 25891
rect 46029 25857 46063 25891
rect 46489 25857 46523 25891
rect 26341 25789 26375 25823
rect 29193 25789 29227 25823
rect 36829 25789 36863 25823
rect 37841 25789 37875 25823
rect 41245 25789 41279 25823
rect 28641 25721 28675 25755
rect 38209 25721 38243 25755
rect 27261 25653 27295 25687
rect 27905 25653 27939 25687
rect 30941 25653 30975 25687
rect 33609 25653 33643 25687
rect 39865 25653 39899 25687
rect 40693 25653 40727 25687
rect 41981 25653 42015 25687
rect 27537 25449 27571 25483
rect 33885 25449 33919 25483
rect 34069 25449 34103 25483
rect 35265 25449 35299 25483
rect 39313 25449 39347 25483
rect 40049 25449 40083 25483
rect 41061 25449 41095 25483
rect 30941 25381 30975 25415
rect 39129 25381 39163 25415
rect 41705 25381 41739 25415
rect 33149 25313 33183 25347
rect 38117 25313 38151 25347
rect 40877 25313 40911 25347
rect 42349 25313 42383 25347
rect 26893 25245 26927 25279
rect 30481 25245 30515 25279
rect 33425 25245 33459 25279
rect 35081 25245 35115 25279
rect 35265 25245 35299 25279
rect 35909 25245 35943 25279
rect 40049 25245 40083 25279
rect 40233 25245 40267 25279
rect 41153 25245 41187 25279
rect 42441 25245 42475 25279
rect 43361 25245 43395 25279
rect 45201 25245 45235 25279
rect 26985 25177 27019 25211
rect 31401 25177 31435 25211
rect 34053 25177 34087 25211
rect 34253 25177 34287 25211
rect 36185 25177 36219 25211
rect 38853 25177 38887 25211
rect 42809 25177 42843 25211
rect 44097 25177 44131 25211
rect 45477 25177 45511 25211
rect 30481 25109 30515 25143
rect 35449 25109 35483 25143
rect 37657 25109 37691 25143
rect 40417 25109 40451 25143
rect 40877 25109 40911 25143
rect 42165 25109 42199 25143
rect 44189 25109 44223 25143
rect 31033 24905 31067 24939
rect 32873 24905 32907 24939
rect 41061 24905 41095 24939
rect 41153 24905 41187 24939
rect 42809 24905 42843 24939
rect 42977 24905 43011 24939
rect 43177 24837 43211 24871
rect 31769 24769 31803 24803
rect 34161 24769 34195 24803
rect 34253 24769 34287 24803
rect 34345 24769 34379 24803
rect 34529 24769 34563 24803
rect 35817 24769 35851 24803
rect 36461 24769 36495 24803
rect 37933 24769 37967 24803
rect 38117 24769 38151 24803
rect 38577 24769 38611 24803
rect 39221 24769 39255 24803
rect 39773 24769 39807 24803
rect 40969 24769 41003 24803
rect 41337 24769 41371 24803
rect 43821 24769 43855 24803
rect 44833 24769 44867 24803
rect 44925 24769 44959 24803
rect 45292 24769 45326 24803
rect 45937 24769 45971 24803
rect 24225 24701 24259 24735
rect 25053 24701 25087 24735
rect 33885 24701 33919 24735
rect 35541 24701 35575 24735
rect 38485 24701 38519 24735
rect 41429 24701 41463 24735
rect 35633 24633 35667 24667
rect 36829 24633 36863 24667
rect 41889 24633 41923 24667
rect 45477 24633 45511 24667
rect 28273 24565 28307 24599
rect 33425 24565 33459 24599
rect 34989 24565 35023 24599
rect 35725 24565 35759 24599
rect 36921 24565 36955 24599
rect 40049 24565 40083 24599
rect 40693 24565 40727 24599
rect 42993 24565 43027 24599
rect 43913 24565 43947 24599
rect 34161 24361 34195 24395
rect 35725 24361 35759 24395
rect 39405 24361 39439 24395
rect 40693 24361 40727 24395
rect 44465 24361 44499 24395
rect 38485 24293 38519 24327
rect 42809 24293 42843 24327
rect 28917 24225 28951 24259
rect 29193 24225 29227 24259
rect 30573 24225 30607 24259
rect 33057 24225 33091 24259
rect 40785 24225 40819 24259
rect 42625 24225 42659 24259
rect 25973 24157 26007 24191
rect 26617 24157 26651 24191
rect 27905 24157 27939 24191
rect 28089 24157 28123 24191
rect 28825 24157 28859 24191
rect 30481 24157 30515 24191
rect 31309 24157 31343 24191
rect 33333 24157 33367 24191
rect 34069 24157 34103 24191
rect 34253 24157 34287 24191
rect 35541 24157 35575 24191
rect 35817 24157 35851 24191
rect 36737 24157 36771 24191
rect 36921 24157 36955 24191
rect 37105 24157 37139 24191
rect 37289 24157 37323 24191
rect 38715 24157 38749 24191
rect 38945 24157 38979 24191
rect 40322 24157 40356 24191
rect 41521 24157 41555 24191
rect 41610 24151 41644 24185
rect 41705 24157 41739 24191
rect 41889 24157 41923 24191
rect 42901 24157 42935 24191
rect 43913 24157 43947 24191
rect 46213 24157 46247 24191
rect 27445 24089 27479 24123
rect 37013 24089 37047 24123
rect 38853 24089 38887 24123
rect 43545 24089 43579 24123
rect 45293 24089 45327 24123
rect 45661 24089 45695 24123
rect 27905 24021 27939 24055
rect 30113 24021 30147 24055
rect 35357 24021 35391 24055
rect 37933 24021 37967 24055
rect 40141 24021 40175 24055
rect 40325 24021 40359 24055
rect 41245 24021 41279 24055
rect 42441 24021 42475 24055
rect 46305 24021 46339 24055
rect 24961 23817 24995 23851
rect 29101 23817 29135 23851
rect 37473 23817 37507 23851
rect 43361 23817 43395 23851
rect 44532 23817 44566 23851
rect 24409 23749 24443 23783
rect 27169 23749 27203 23783
rect 28241 23749 28275 23783
rect 28457 23749 28491 23783
rect 30113 23749 30147 23783
rect 41981 23749 42015 23783
rect 1869 23681 1903 23715
rect 24317 23681 24351 23715
rect 24501 23681 24535 23715
rect 25237 23681 25271 23715
rect 26617 23681 26651 23715
rect 27353 23681 27387 23715
rect 29101 23681 29135 23715
rect 29285 23681 29319 23715
rect 31585 23681 31619 23715
rect 32505 23681 32539 23715
rect 32689 23681 32723 23715
rect 32965 23681 32999 23715
rect 33149 23681 33183 23715
rect 33977 23681 34011 23715
rect 34805 23681 34839 23715
rect 35817 23681 35851 23715
rect 36829 23681 36863 23715
rect 37657 23681 37691 23715
rect 38669 23681 38703 23715
rect 39681 23681 39715 23715
rect 40877 23681 40911 23715
rect 41153 23681 41187 23715
rect 43177 23681 43211 23715
rect 43453 23681 43487 23715
rect 44097 23681 44131 23715
rect 44833 23681 44867 23715
rect 25145 23613 25179 23647
rect 25329 23613 25363 23647
rect 25421 23613 25455 23647
rect 26341 23613 26375 23647
rect 27629 23613 27663 23647
rect 31677 23613 31711 23647
rect 33609 23613 33643 23647
rect 35909 23613 35943 23647
rect 37749 23613 37783 23647
rect 37841 23613 37875 23647
rect 37933 23613 37967 23647
rect 40693 23613 40727 23647
rect 44925 23613 44959 23647
rect 26525 23545 26559 23579
rect 27537 23545 27571 23579
rect 28089 23545 28123 23579
rect 30481 23545 30515 23579
rect 31217 23545 31251 23579
rect 41061 23545 41095 23579
rect 45753 23545 45787 23579
rect 1685 23477 1719 23511
rect 2421 23477 2455 23511
rect 26433 23477 26467 23511
rect 28273 23477 28307 23511
rect 30573 23477 30607 23511
rect 33701 23477 33735 23511
rect 33793 23477 33827 23511
rect 33977 23477 34011 23511
rect 34529 23477 34563 23511
rect 36001 23477 36035 23511
rect 36185 23477 36219 23511
rect 36737 23477 36771 23511
rect 38761 23477 38795 23511
rect 39497 23477 39531 23511
rect 41705 23477 41739 23511
rect 42993 23477 43027 23511
rect 23489 23273 23523 23307
rect 34253 23273 34287 23307
rect 35909 23273 35943 23307
rect 31125 23205 31159 23239
rect 43545 23205 43579 23239
rect 26433 23137 26467 23171
rect 27445 23137 27479 23171
rect 27905 23137 27939 23171
rect 28641 23137 28675 23171
rect 29193 23137 29227 23171
rect 30849 23137 30883 23171
rect 32413 23137 32447 23171
rect 36645 23137 36679 23171
rect 40325 23137 40359 23171
rect 41889 23137 41923 23171
rect 21925 23069 21959 23103
rect 22017 23069 22051 23103
rect 23213 23069 23247 23103
rect 25145 23069 25179 23103
rect 25421 23069 25455 23103
rect 25605 23069 25639 23103
rect 26065 23069 26099 23103
rect 26249 23069 26283 23103
rect 27813 23069 27847 23103
rect 29745 23069 29779 23103
rect 30297 23069 30331 23103
rect 30757 23069 30791 23103
rect 32321 23069 32355 23103
rect 33241 23069 33275 23103
rect 33425 23069 33459 23103
rect 34161 23069 34195 23103
rect 34345 23069 34379 23103
rect 34897 23069 34931 23103
rect 35081 23069 35115 23103
rect 36553 23069 36587 23103
rect 36737 23069 36771 23103
rect 37565 23069 37599 23103
rect 38945 23069 38979 23103
rect 39313 23069 39347 23103
rect 39405 23069 39439 23103
rect 40233 23069 40267 23103
rect 40417 23069 40451 23103
rect 40509 23069 40543 23103
rect 40693 23069 40727 23103
rect 41245 23069 41279 23103
rect 41429 23069 41463 23103
rect 42073 23069 42107 23103
rect 42165 23069 42199 23103
rect 42717 23069 42751 23103
rect 45569 23069 45603 23103
rect 46121 23069 46155 23103
rect 35725 23001 35759 23035
rect 35941 23001 35975 23035
rect 38761 23001 38795 23035
rect 43821 23001 43855 23035
rect 45201 23001 45235 23035
rect 21741 22933 21775 22967
rect 22385 22933 22419 22967
rect 23673 22933 23707 22967
rect 24961 22933 24995 22967
rect 31677 22933 31711 22967
rect 33333 22933 33367 22967
rect 34989 22933 35023 22967
rect 36093 22933 36127 22967
rect 37841 22933 37875 22967
rect 40049 22933 40083 22967
rect 41337 22933 41371 22967
rect 43361 22933 43395 22967
rect 44281 22933 44315 22967
rect 22845 22729 22879 22763
rect 24593 22729 24627 22763
rect 24961 22729 24995 22763
rect 27261 22729 27295 22763
rect 27813 22729 27847 22763
rect 32413 22729 32447 22763
rect 32781 22729 32815 22763
rect 35173 22729 35207 22763
rect 39497 22729 39531 22763
rect 41889 22729 41923 22763
rect 29009 22661 29043 22695
rect 30757 22661 30791 22695
rect 35725 22661 35759 22695
rect 41245 22661 41279 22695
rect 57437 22661 57471 22695
rect 23581 22593 23615 22627
rect 23857 22593 23891 22627
rect 24777 22593 24811 22627
rect 24869 22593 24903 22627
rect 25237 22593 25271 22627
rect 27169 22593 27203 22627
rect 27353 22593 27387 22627
rect 28181 22593 28215 22627
rect 28273 22593 28307 22627
rect 30941 22593 30975 22627
rect 32597 22593 32631 22627
rect 32873 22593 32907 22627
rect 34161 22593 34195 22627
rect 34253 22593 34287 22627
rect 34437 22593 34471 22627
rect 34529 22593 34563 22627
rect 34989 22593 35023 22627
rect 35265 22593 35299 22627
rect 35909 22593 35943 22627
rect 36139 22593 36173 22627
rect 36369 22593 36403 22627
rect 36829 22593 36863 22627
rect 38025 22593 38059 22627
rect 38301 22593 38335 22627
rect 40325 22593 40359 22627
rect 40417 22593 40451 22627
rect 41153 22593 41187 22627
rect 41337 22593 41371 22627
rect 41797 22593 41831 22627
rect 41981 22593 42015 22627
rect 42901 22593 42935 22627
rect 43637 22593 43671 22627
rect 45017 22593 45051 22627
rect 45569 22593 45603 22627
rect 46121 22593 46155 22627
rect 58081 22593 58115 22627
rect 25145 22525 25179 22559
rect 28457 22525 28491 22559
rect 29837 22525 29871 22559
rect 36001 22525 36035 22559
rect 36277 22525 36311 22559
rect 37933 22525 37967 22559
rect 38393 22525 38427 22559
rect 38853 22525 38887 22559
rect 39037 22525 39071 22559
rect 39129 22525 39163 22559
rect 40141 22525 40175 22559
rect 40233 22525 40267 22559
rect 42625 22525 42659 22559
rect 44557 22525 44591 22559
rect 46397 22525 46431 22559
rect 33977 22457 34011 22491
rect 34989 22457 35023 22491
rect 42717 22457 42751 22491
rect 45293 22457 45327 22491
rect 58265 22457 58299 22491
rect 30573 22389 30607 22423
rect 31401 22389 31435 22423
rect 33425 22389 33459 22423
rect 37749 22389 37783 22423
rect 39957 22389 39991 22423
rect 43085 22389 43119 22423
rect 43913 22389 43947 22423
rect 25053 22185 25087 22219
rect 35081 22185 35115 22219
rect 38209 22185 38243 22219
rect 42901 22185 42935 22219
rect 44189 22185 44223 22219
rect 25881 22117 25915 22151
rect 32965 22117 32999 22151
rect 26525 22049 26559 22083
rect 26985 22049 27019 22083
rect 32689 22049 32723 22083
rect 33057 22049 33091 22083
rect 35725 22049 35759 22083
rect 36737 22049 36771 22083
rect 38485 22049 38519 22083
rect 38669 22049 38703 22083
rect 39313 22049 39347 22083
rect 40693 22049 40727 22083
rect 42349 22049 42383 22083
rect 22201 21981 22235 22015
rect 25145 21981 25179 22015
rect 25605 21981 25639 22015
rect 25789 21981 25823 22015
rect 26893 21981 26927 22015
rect 30573 21981 30607 22015
rect 30849 21981 30883 22015
rect 31493 21981 31527 22015
rect 31585 21981 31619 22015
rect 31677 21981 31711 22015
rect 31769 21981 31803 22015
rect 32841 21981 32875 22015
rect 33149 21981 33183 22015
rect 33885 21981 33919 22015
rect 34069 21981 34103 22015
rect 34897 21981 34931 22015
rect 35909 21981 35943 22015
rect 36001 21981 36035 22015
rect 36129 21981 36163 22015
rect 37381 21981 37415 22015
rect 38393 21981 38427 22015
rect 38577 21981 38611 22015
rect 40049 21981 40083 22015
rect 40233 21981 40267 22015
rect 43088 21959 43122 21993
rect 43177 21981 43211 22015
rect 43361 21981 43395 22015
rect 43453 21981 43487 22015
rect 44097 21981 44131 22015
rect 44189 21981 44223 22015
rect 45385 21981 45419 22015
rect 45661 21981 45695 22015
rect 45845 21981 45879 22015
rect 21189 21913 21223 21947
rect 23397 21913 23431 21947
rect 23765 21913 23799 21947
rect 37197 21913 37231 21947
rect 37749 21913 37783 21947
rect 42073 21913 42107 21947
rect 23305 21845 23339 21879
rect 23489 21845 23523 21879
rect 23581 21845 23615 21879
rect 31309 21845 31343 21879
rect 33701 21845 33735 21879
rect 40049 21845 40083 21879
rect 41245 21845 41279 21879
rect 45201 21845 45235 21879
rect 23673 21641 23707 21675
rect 23765 21641 23799 21675
rect 25513 21641 25547 21675
rect 29009 21641 29043 21675
rect 30205 21641 30239 21675
rect 31033 21641 31067 21675
rect 32413 21641 32447 21675
rect 34529 21641 34563 21675
rect 35725 21641 35759 21675
rect 44833 21641 44867 21675
rect 45937 21641 45971 21675
rect 30297 21573 30331 21607
rect 32597 21573 32631 21607
rect 33885 21573 33919 21607
rect 34989 21573 35023 21607
rect 42073 21573 42107 21607
rect 42717 21573 42751 21607
rect 23581 21505 23615 21539
rect 25697 21505 25731 21539
rect 27905 21505 27939 21539
rect 31217 21505 31251 21539
rect 31401 21505 31435 21539
rect 32321 21505 32355 21539
rect 33793 21505 33827 21539
rect 33977 21505 34011 21539
rect 34713 21505 34747 21539
rect 34805 21505 34839 21539
rect 35541 21505 35575 21539
rect 35725 21505 35759 21539
rect 36185 21505 36219 21539
rect 36277 21505 36311 21539
rect 37565 21505 37599 21539
rect 37749 21505 37783 21539
rect 38209 21505 38243 21539
rect 38577 21505 38611 21539
rect 38761 21505 38795 21539
rect 39589 21505 39623 21539
rect 39865 21505 39899 21539
rect 40601 21505 40635 21539
rect 40785 21505 40819 21539
rect 40877 21505 40911 21539
rect 41061 21505 41095 21539
rect 43637 21505 43671 21539
rect 43913 21505 43947 21539
rect 44649 21505 44683 21539
rect 45017 21505 45051 21539
rect 45293 21505 45327 21539
rect 45753 21505 45787 21539
rect 46489 21505 46523 21539
rect 22109 21437 22143 21471
rect 22845 21437 22879 21471
rect 24041 21437 24075 21471
rect 25973 21437 26007 21471
rect 29101 21437 29135 21471
rect 29285 21437 29319 21471
rect 30481 21437 30515 21471
rect 36461 21437 36495 21471
rect 39681 21437 39715 21471
rect 43545 21437 43579 21471
rect 32597 21369 32631 21403
rect 38301 21369 38335 21403
rect 39773 21369 39807 21403
rect 40969 21369 41003 21403
rect 41613 21369 41647 21403
rect 41705 21369 41739 21403
rect 25881 21301 25915 21335
rect 28089 21301 28123 21335
rect 28641 21301 28675 21335
rect 29837 21301 29871 21335
rect 34989 21301 35023 21335
rect 36369 21301 36403 21335
rect 37565 21301 37599 21335
rect 39405 21301 39439 21335
rect 42809 21301 42843 21335
rect 45017 21301 45051 21335
rect 46673 21301 46707 21335
rect 23489 21097 23523 21131
rect 25789 21097 25823 21131
rect 32413 21097 32447 21131
rect 38025 21097 38059 21131
rect 41061 21097 41095 21131
rect 41889 21097 41923 21131
rect 46213 21097 46247 21131
rect 28365 21029 28399 21063
rect 38853 21029 38887 21063
rect 27629 20961 27663 20995
rect 30205 20961 30239 20995
rect 32597 20961 32631 20995
rect 33609 20961 33643 20995
rect 36921 20961 36955 20995
rect 39037 20961 39071 20995
rect 40141 20961 40175 20995
rect 42901 20961 42935 20995
rect 23673 20893 23707 20927
rect 23857 20893 23891 20927
rect 25145 20893 25179 20927
rect 25329 20893 25363 20927
rect 25789 20893 25823 20927
rect 25881 20893 25915 20927
rect 30113 20893 30147 20927
rect 32321 20893 32355 20927
rect 33793 20893 33827 20927
rect 33885 20893 33919 20927
rect 35725 20893 35759 20927
rect 36553 20893 36587 20927
rect 36645 20893 36679 20927
rect 37013 20893 37047 20927
rect 38209 20893 38243 20927
rect 39129 20893 39163 20927
rect 40325 20893 40359 20927
rect 41705 20893 41739 20927
rect 42625 20893 42659 20927
rect 42717 20893 42751 20927
rect 42809 20893 42843 20927
rect 43085 20893 43119 20927
rect 43729 20893 43763 20927
rect 43913 20893 43947 20927
rect 45293 20893 45327 20927
rect 45753 20893 45787 20927
rect 26065 20825 26099 20859
rect 27353 20825 27387 20859
rect 35909 20825 35943 20859
rect 37473 20825 37507 20859
rect 38393 20825 38427 20859
rect 39405 20825 39439 20859
rect 39497 20825 39531 20859
rect 45385 20825 45419 20859
rect 24961 20757 24995 20791
rect 26985 20757 27019 20791
rect 27445 20757 27479 20791
rect 29745 20757 29779 20791
rect 31861 20757 31895 20791
rect 32597 20757 32631 20791
rect 33149 20757 33183 20791
rect 33609 20757 33643 20791
rect 35541 20757 35575 20791
rect 36369 20757 36403 20791
rect 36829 20757 36863 20791
rect 40509 20757 40543 20791
rect 42441 20757 42475 20791
rect 43545 20757 43579 20791
rect 44373 20757 44407 20791
rect 28733 20553 28767 20587
rect 35817 20553 35851 20587
rect 37565 20553 37599 20587
rect 38577 20553 38611 20587
rect 39405 20553 39439 20587
rect 44531 20553 44565 20587
rect 23673 20485 23707 20519
rect 32321 20485 32355 20519
rect 35633 20485 35667 20519
rect 38853 20485 38887 20519
rect 40141 20485 40175 20519
rect 40341 20485 40375 20519
rect 42625 20485 42659 20519
rect 44741 20485 44775 20519
rect 45477 20485 45511 20519
rect 25697 20417 25731 20451
rect 27537 20417 27571 20451
rect 27721 20417 27755 20451
rect 29009 20417 29043 20451
rect 30205 20417 30239 20451
rect 30389 20417 30423 20451
rect 31125 20417 31159 20451
rect 31309 20417 31343 20451
rect 31401 20417 31435 20451
rect 31585 20417 31619 20451
rect 31677 20417 31711 20451
rect 32597 20417 32631 20451
rect 32689 20417 32723 20451
rect 32781 20417 32815 20451
rect 32965 20417 32999 20451
rect 33885 20417 33919 20451
rect 34713 20417 34747 20451
rect 35909 20417 35943 20451
rect 36369 20417 36403 20451
rect 36553 20417 36587 20451
rect 37473 20417 37507 20451
rect 37749 20417 37783 20451
rect 39405 20417 39439 20451
rect 39589 20417 39623 20451
rect 40969 20417 41003 20451
rect 41153 20417 41187 20451
rect 41797 20417 41831 20451
rect 41981 20417 42015 20451
rect 42717 20417 42751 20451
rect 42901 20417 42935 20451
rect 43637 20417 43671 20451
rect 43821 20417 43855 20451
rect 45201 20417 45235 20451
rect 45661 20417 45695 20451
rect 22845 20349 22879 20383
rect 24685 20349 24719 20383
rect 28733 20349 28767 20383
rect 28917 20349 28951 20383
rect 34161 20349 34195 20383
rect 36461 20349 36495 20383
rect 27537 20281 27571 20315
rect 35633 20281 35667 20315
rect 37749 20281 37783 20315
rect 43637 20281 43671 20315
rect 29745 20213 29779 20247
rect 30297 20213 30331 20247
rect 33701 20213 33735 20247
rect 34069 20213 34103 20247
rect 34897 20213 34931 20247
rect 40325 20213 40359 20247
rect 40509 20213 40543 20247
rect 41153 20213 41187 20247
rect 41797 20213 41831 20247
rect 44373 20213 44407 20247
rect 44557 20213 44591 20247
rect 23213 20009 23247 20043
rect 23673 20009 23707 20043
rect 24041 20009 24075 20043
rect 25789 20009 25823 20043
rect 27261 20009 27295 20043
rect 27445 20009 27479 20043
rect 30757 20009 30791 20043
rect 32045 20009 32079 20043
rect 33333 20009 33367 20043
rect 34345 20009 34379 20043
rect 46213 20009 46247 20043
rect 25697 19941 25731 19975
rect 26249 19941 26283 19975
rect 27813 19941 27847 19975
rect 35909 19941 35943 19975
rect 41705 19941 41739 19975
rect 42441 19941 42475 19975
rect 44649 19941 44683 19975
rect 22845 19873 22879 19907
rect 26709 19873 26743 19907
rect 28733 19873 28767 19907
rect 31769 19873 31803 19907
rect 32689 19873 32723 19907
rect 41613 19873 41647 19907
rect 44281 19873 44315 19907
rect 44465 19873 44499 19907
rect 45201 19873 45235 19907
rect 23029 19805 23063 19839
rect 23673 19805 23707 19839
rect 23857 19805 23891 19839
rect 26617 19805 26651 19839
rect 28273 19805 28307 19839
rect 28457 19805 28491 19839
rect 28825 19805 28859 19839
rect 30113 19805 30147 19839
rect 30292 19805 30326 19839
rect 30408 19799 30442 19833
rect 30527 19805 30561 19839
rect 31847 19805 31881 19839
rect 33517 19805 33551 19839
rect 33793 19805 33827 19839
rect 35909 19805 35943 19839
rect 36093 19805 36127 19839
rect 36185 19805 36219 19839
rect 37289 19805 37323 19839
rect 37473 19805 37507 19839
rect 37933 19805 37967 19839
rect 38117 19805 38151 19839
rect 38853 19805 38887 19839
rect 38945 19805 38979 19839
rect 39221 19805 39255 19839
rect 40049 19805 40083 19839
rect 40233 19805 40267 19839
rect 40325 19805 40359 19839
rect 40509 19805 40543 19839
rect 40601 19805 40635 19839
rect 41521 19805 41555 19839
rect 41797 19805 41831 19839
rect 41981 19805 42015 19839
rect 42717 19805 42751 19839
rect 43821 19805 43855 19839
rect 44373 19805 44407 19839
rect 45385 19805 45419 19839
rect 45477 19805 45511 19839
rect 45661 19805 45695 19839
rect 45753 19805 45787 19839
rect 25329 19737 25363 19771
rect 27445 19737 27479 19771
rect 33701 19737 33735 19771
rect 39037 19737 39071 19771
rect 42441 19737 42475 19771
rect 44649 19737 44683 19771
rect 35449 19669 35483 19703
rect 36645 19669 36679 19703
rect 37381 19669 37415 19703
rect 38025 19669 38059 19703
rect 38669 19669 38703 19703
rect 41337 19669 41371 19703
rect 42625 19669 42659 19703
rect 43637 19669 43671 19703
rect 23489 19465 23523 19499
rect 27261 19465 27295 19499
rect 37473 19465 37507 19499
rect 40509 19465 40543 19499
rect 44097 19465 44131 19499
rect 44281 19465 44315 19499
rect 45109 19465 45143 19499
rect 46029 19465 46063 19499
rect 36829 19397 36863 19431
rect 41521 19397 41555 19431
rect 42073 19397 42107 19431
rect 23673 19329 23707 19363
rect 23765 19329 23799 19363
rect 24225 19329 24259 19363
rect 24409 19329 24443 19363
rect 25329 19329 25363 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 28641 19329 28675 19363
rect 29285 19329 29319 19363
rect 29469 19329 29503 19363
rect 29561 19329 29595 19363
rect 29745 19329 29779 19363
rect 29837 19329 29871 19363
rect 30297 19329 30331 19363
rect 30481 19329 30515 19363
rect 32597 19329 32631 19363
rect 32689 19329 32723 19363
rect 32965 19329 32999 19363
rect 34345 19329 34379 19363
rect 34437 19329 34471 19363
rect 34621 19329 34655 19363
rect 35357 19329 35391 19363
rect 35449 19329 35483 19363
rect 36369 19329 36403 19363
rect 36553 19329 36587 19363
rect 37749 19329 37783 19363
rect 37841 19329 37875 19363
rect 37933 19329 37967 19363
rect 38117 19329 38151 19363
rect 39129 19329 39163 19363
rect 39221 19329 39255 19363
rect 39313 19329 39347 19363
rect 39497 19329 39531 19363
rect 40417 19329 40451 19363
rect 40601 19329 40635 19363
rect 41245 19329 41279 19363
rect 43085 19329 43119 19363
rect 43269 19329 43303 19363
rect 43913 19329 43947 19363
rect 45569 19329 45603 19363
rect 23489 19261 23523 19295
rect 25421 19261 25455 19295
rect 28825 19261 28859 19295
rect 32413 19261 32447 19295
rect 34529 19261 34563 19295
rect 35541 19261 35575 19295
rect 35633 19261 35667 19295
rect 41521 19261 41555 19295
rect 44005 19261 44039 19295
rect 44373 19261 44407 19295
rect 30297 19193 30331 19227
rect 31493 19193 31527 19227
rect 32873 19193 32907 19227
rect 36185 19193 36219 19227
rect 43729 19193 43763 19227
rect 24317 19125 24351 19159
rect 25697 19125 25731 19159
rect 28457 19125 28491 19159
rect 33425 19125 33459 19159
rect 34161 19125 34195 19159
rect 35173 19125 35207 19159
rect 36737 19125 36771 19159
rect 38853 19125 38887 19159
rect 41337 19125 41371 19159
rect 43085 19125 43119 19159
rect 45293 19125 45327 19159
rect 23581 18921 23615 18955
rect 25973 18921 26007 18955
rect 27629 18921 27663 18955
rect 35449 18921 35483 18955
rect 36185 18921 36219 18955
rect 39497 18921 39531 18955
rect 42717 18921 42751 18955
rect 44373 18921 44407 18955
rect 46213 18921 46247 18955
rect 27813 18853 27847 18887
rect 34897 18853 34931 18887
rect 37473 18853 37507 18887
rect 37565 18853 37599 18887
rect 43453 18853 43487 18887
rect 45293 18853 45327 18887
rect 23397 18785 23431 18819
rect 33977 18785 34011 18819
rect 37197 18785 37231 18819
rect 41245 18785 41279 18819
rect 41889 18785 41923 18819
rect 43177 18785 43211 18819
rect 23305 18717 23339 18751
rect 24777 18717 24811 18751
rect 24961 18717 24995 18751
rect 25789 18717 25823 18751
rect 25973 18717 26007 18751
rect 31033 18717 31067 18751
rect 31125 18717 31159 18751
rect 31217 18717 31251 18751
rect 31401 18717 31435 18751
rect 32229 18717 32263 18751
rect 33057 18717 33091 18751
rect 33149 18717 33183 18751
rect 34161 18717 34195 18751
rect 34345 18717 34379 18751
rect 35022 18717 35056 18751
rect 35541 18717 35575 18751
rect 37390 18711 37424 18745
rect 37657 18717 37691 18751
rect 37841 18717 37875 18751
rect 40754 18717 40788 18751
rect 41153 18717 41187 18751
rect 42349 18717 42383 18751
rect 43361 18717 43395 18751
rect 43545 18717 43579 18751
rect 43637 18717 43671 18751
rect 43821 18717 43855 18751
rect 44465 18717 44499 18751
rect 45201 18717 45235 18751
rect 45661 18717 45695 18751
rect 28089 18649 28123 18683
rect 28549 18649 28583 18683
rect 31861 18649 31895 18683
rect 32045 18649 32079 18683
rect 33425 18649 33459 18683
rect 33517 18649 33551 18683
rect 36369 18649 36403 18683
rect 36553 18649 36587 18683
rect 39129 18649 39163 18683
rect 39313 18649 39347 18683
rect 42533 18649 42567 18683
rect 24593 18581 24627 18615
rect 30757 18581 30791 18615
rect 32873 18581 32907 18615
rect 35081 18581 35115 18615
rect 38669 18581 38703 18615
rect 40049 18581 40083 18615
rect 40601 18581 40635 18615
rect 40785 18581 40819 18615
rect 30373 18377 30407 18411
rect 33241 18377 33275 18411
rect 39681 18377 39715 18411
rect 39773 18377 39807 18411
rect 41061 18377 41095 18411
rect 42809 18377 42843 18411
rect 43821 18377 43855 18411
rect 30573 18309 30607 18343
rect 31125 18309 31159 18343
rect 43361 18309 43395 18343
rect 23581 18241 23615 18275
rect 23857 18241 23891 18275
rect 24593 18241 24627 18275
rect 25697 18241 25731 18275
rect 27537 18241 27571 18275
rect 29009 18241 29043 18275
rect 31401 18241 31435 18275
rect 32781 18241 32815 18275
rect 33241 18241 33275 18275
rect 33425 18241 33459 18275
rect 34713 18241 34747 18275
rect 34897 18241 34931 18275
rect 35909 18241 35943 18275
rect 36001 18241 36035 18275
rect 36185 18241 36219 18275
rect 36277 18241 36311 18275
rect 38301 18241 38335 18275
rect 38485 18241 38519 18275
rect 38761 18241 38795 18275
rect 39497 18241 39531 18275
rect 39865 18241 39899 18275
rect 40877 18241 40911 18275
rect 42809 18241 42843 18275
rect 43821 18241 43855 18275
rect 44005 18241 44039 18275
rect 45109 18241 45143 18275
rect 45385 18241 45419 18275
rect 25605 18173 25639 18207
rect 27629 18173 27663 18207
rect 28733 18173 28767 18207
rect 31125 18173 31159 18207
rect 38578 18173 38612 18207
rect 39405 18173 39439 18207
rect 41245 18173 41279 18207
rect 42717 18173 42751 18207
rect 24317 18105 24351 18139
rect 28825 18105 28859 18139
rect 38669 18105 38703 18139
rect 25329 18037 25363 18071
rect 27261 18037 27295 18071
rect 28917 18037 28951 18071
rect 30205 18037 30239 18071
rect 30389 18037 30423 18071
rect 31309 18037 31343 18071
rect 32321 18037 32355 18071
rect 32597 18037 32631 18071
rect 33885 18037 33919 18071
rect 35081 18037 35115 18071
rect 35725 18037 35759 18071
rect 36829 18037 36863 18071
rect 38945 18037 38979 18071
rect 40141 18037 40175 18071
rect 40693 18037 40727 18071
rect 44465 18037 44499 18071
rect 45477 18037 45511 18071
rect 24685 17833 24719 17867
rect 27169 17833 27203 17867
rect 29745 17833 29779 17867
rect 32965 17833 32999 17867
rect 33425 17833 33459 17867
rect 38209 17833 38243 17867
rect 41521 17833 41555 17867
rect 43545 17833 43579 17867
rect 25513 17765 25547 17799
rect 27353 17765 27387 17799
rect 30113 17765 30147 17799
rect 31861 17765 31895 17799
rect 35541 17765 35575 17799
rect 38853 17765 38887 17799
rect 44189 17765 44223 17799
rect 45201 17765 45235 17799
rect 30021 17697 30055 17731
rect 30941 17697 30975 17731
rect 34069 17697 34103 17731
rect 35449 17697 35483 17731
rect 37933 17697 37967 17731
rect 42257 17697 42291 17731
rect 24593 17629 24627 17663
rect 24777 17629 24811 17663
rect 25697 17629 25731 17663
rect 25881 17629 25915 17663
rect 25973 17629 26007 17663
rect 26433 17629 26467 17663
rect 26617 17629 26651 17663
rect 29929 17629 29963 17663
rect 30205 17629 30239 17663
rect 31401 17629 31435 17663
rect 32045 17629 32079 17663
rect 32137 17629 32171 17663
rect 35968 17629 36002 17663
rect 36829 17629 36863 17663
rect 36922 17629 36956 17663
rect 37105 17629 37139 17663
rect 37335 17629 37369 17663
rect 38393 17629 38427 17663
rect 38853 17629 38887 17663
rect 39129 17629 39163 17663
rect 40141 17629 40175 17663
rect 40417 17629 40451 17663
rect 40969 17639 41003 17673
rect 41061 17629 41095 17663
rect 41245 17629 41279 17663
rect 41334 17629 41368 17663
rect 42717 17629 42751 17663
rect 44465 17629 44499 17663
rect 45201 17629 45235 17663
rect 45385 17629 45419 17663
rect 45845 17629 45879 17663
rect 46029 17629 46063 17663
rect 27629 17561 27663 17595
rect 31861 17561 31895 17595
rect 37197 17561 37231 17595
rect 42395 17561 42429 17595
rect 42533 17561 42567 17595
rect 42625 17561 42659 17595
rect 43529 17561 43563 17595
rect 43729 17561 43763 17595
rect 44189 17561 44223 17595
rect 26525 17493 26559 17527
rect 28181 17493 28215 17527
rect 31217 17493 31251 17527
rect 31309 17493 31343 17527
rect 33793 17493 33827 17527
rect 33885 17493 33919 17527
rect 35909 17493 35943 17527
rect 36093 17493 36127 17527
rect 37473 17493 37507 17527
rect 39037 17493 39071 17527
rect 40325 17493 40359 17527
rect 42901 17493 42935 17527
rect 43361 17493 43395 17527
rect 44373 17493 44407 17527
rect 45845 17493 45879 17527
rect 32321 17289 32355 17323
rect 33425 17289 33459 17323
rect 34069 17289 34103 17323
rect 37657 17289 37691 17323
rect 40785 17289 40819 17323
rect 42073 17289 42107 17323
rect 25237 17221 25271 17255
rect 33241 17221 33275 17255
rect 34437 17221 34471 17255
rect 35249 17221 35283 17255
rect 35449 17221 35483 17255
rect 43269 17221 43303 17255
rect 1869 17153 1903 17187
rect 2421 17153 2455 17187
rect 23673 17153 23707 17187
rect 24225 17153 24259 17187
rect 25605 17153 25639 17187
rect 26065 17153 26099 17187
rect 29193 17153 29227 17187
rect 30113 17153 30147 17187
rect 32597 17153 32631 17187
rect 33517 17153 33551 17187
rect 34253 17153 34287 17187
rect 34345 17153 34379 17187
rect 34621 17153 34655 17187
rect 35909 17153 35943 17187
rect 36093 17153 36127 17187
rect 36553 17153 36587 17187
rect 36737 17153 36771 17187
rect 37473 17153 37507 17187
rect 37749 17153 37783 17187
rect 39221 17153 39255 17187
rect 39405 17153 39439 17187
rect 39865 17153 39899 17187
rect 40693 17153 40727 17187
rect 40969 17153 41003 17187
rect 41429 17153 41463 17187
rect 42625 17153 42659 17187
rect 42809 17153 42843 17187
rect 42901 17153 42935 17187
rect 43039 17153 43073 17187
rect 44311 17153 44345 17187
rect 44465 17153 44499 17187
rect 44925 17153 44959 17187
rect 45385 17153 45419 17187
rect 58081 17153 58115 17187
rect 27629 17085 27663 17119
rect 32321 17085 32355 17119
rect 32505 17085 32539 17119
rect 39957 17085 39991 17119
rect 45017 17085 45051 17119
rect 57437 17085 57471 17119
rect 1685 17017 1719 17051
rect 27261 17017 27295 17051
rect 30665 17017 30699 17051
rect 37473 17017 37507 17051
rect 39405 17017 39439 17051
rect 44097 17017 44131 17051
rect 58265 17017 58299 17051
rect 22845 16949 22879 16983
rect 27169 16949 27203 16983
rect 33241 16949 33275 16983
rect 35081 16949 35115 16983
rect 35265 16949 35299 16983
rect 36001 16949 36035 16983
rect 36553 16949 36587 16983
rect 38485 16949 38519 16983
rect 39957 16949 39991 16983
rect 40233 16949 40267 16983
rect 40969 16949 41003 16983
rect 25053 16745 25087 16779
rect 28641 16745 28675 16779
rect 29009 16745 29043 16779
rect 33977 16745 34011 16779
rect 39221 16745 39255 16779
rect 42349 16745 42383 16779
rect 27629 16677 27663 16711
rect 31677 16677 31711 16711
rect 37933 16677 37967 16711
rect 38209 16677 38243 16711
rect 38301 16677 38335 16711
rect 41061 16677 41095 16711
rect 26893 16609 26927 16643
rect 27997 16609 28031 16643
rect 36277 16609 36311 16643
rect 37013 16609 37047 16643
rect 39037 16609 39071 16643
rect 40049 16609 40083 16643
rect 40325 16609 40359 16643
rect 40417 16609 40451 16643
rect 45201 16609 45235 16643
rect 25237 16541 25271 16575
rect 25329 16541 25363 16575
rect 25513 16541 25547 16575
rect 25605 16541 25639 16575
rect 26801 16541 26835 16575
rect 27813 16541 27847 16575
rect 28549 16541 28583 16575
rect 31585 16541 31619 16575
rect 31953 16541 31987 16575
rect 32229 16541 32263 16575
rect 32413 16541 32447 16575
rect 32597 16541 32631 16575
rect 33057 16541 33091 16575
rect 33333 16541 33367 16575
rect 33977 16541 34011 16575
rect 34253 16541 34287 16575
rect 35633 16541 35667 16575
rect 36369 16541 36403 16575
rect 36921 16541 36955 16575
rect 38117 16541 38151 16575
rect 38393 16541 38427 16575
rect 38577 16541 38611 16575
rect 39313 16541 39347 16575
rect 40233 16541 40267 16575
rect 40509 16541 40543 16575
rect 41245 16541 41279 16575
rect 41337 16541 41371 16575
rect 41521 16541 41555 16575
rect 41613 16541 41647 16575
rect 42165 16541 42199 16575
rect 42257 16541 42291 16575
rect 43361 16541 43395 16575
rect 43453 16541 43487 16575
rect 43637 16541 43671 16575
rect 43729 16541 43763 16575
rect 44373 16541 44407 16575
rect 44557 16541 44591 16575
rect 33241 16473 33275 16507
rect 34161 16473 34195 16507
rect 39037 16473 39071 16507
rect 27169 16405 27203 16439
rect 33155 16405 33189 16439
rect 35541 16405 35575 16439
rect 42533 16405 42567 16439
rect 43913 16405 43947 16439
rect 44373 16405 44407 16439
rect 24869 16201 24903 16235
rect 28365 16201 28399 16235
rect 33333 16201 33367 16235
rect 34621 16201 34655 16235
rect 35449 16201 35483 16235
rect 41521 16201 41555 16235
rect 25053 16133 25087 16167
rect 25789 16133 25823 16167
rect 30573 16133 30607 16167
rect 36461 16133 36495 16167
rect 44189 16133 44223 16167
rect 24777 16065 24811 16099
rect 25513 16065 25547 16099
rect 25605 16065 25639 16099
rect 27445 16065 27479 16099
rect 28549 16065 28583 16099
rect 29469 16065 29503 16099
rect 30389 16065 30423 16099
rect 30665 16065 30699 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 32505 16065 32539 16099
rect 32689 16065 32723 16099
rect 33330 16065 33364 16099
rect 33793 16065 33827 16099
rect 34897 16065 34931 16099
rect 35541 16065 35575 16099
rect 36737 16065 36771 16099
rect 37657 16065 37691 16099
rect 37933 16065 37967 16099
rect 39313 16065 39347 16099
rect 39497 16065 39531 16099
rect 39773 16065 39807 16099
rect 40233 16065 40267 16099
rect 40417 16065 40451 16099
rect 41337 16065 41371 16099
rect 41521 16065 41555 16099
rect 41889 16065 41923 16099
rect 43913 16065 43947 16099
rect 44925 16065 44959 16099
rect 45201 16065 45235 16099
rect 27537 15997 27571 16031
rect 27813 15997 27847 16031
rect 28825 15997 28859 16031
rect 29745 15997 29779 16031
rect 31217 15997 31251 16031
rect 34621 15997 34655 16031
rect 36553 15997 36587 16031
rect 39589 15997 39623 16031
rect 40693 15997 40727 16031
rect 43821 15997 43855 16031
rect 44281 15997 44315 16031
rect 44741 15997 44775 16031
rect 25053 15929 25087 15963
rect 29285 15929 29319 15963
rect 33149 15929 33183 15963
rect 37841 15929 37875 15963
rect 39405 15929 39439 15963
rect 25697 15861 25731 15895
rect 28733 15861 28767 15895
rect 29653 15861 29687 15895
rect 30205 15861 30239 15895
rect 32321 15861 32355 15895
rect 32597 15861 32631 15895
rect 33701 15861 33735 15895
rect 34805 15861 34839 15895
rect 36737 15861 36771 15895
rect 36921 15861 36955 15895
rect 37473 15861 37507 15895
rect 39129 15861 39163 15895
rect 40601 15861 40635 15895
rect 43637 15861 43671 15895
rect 45109 15861 45143 15895
rect 45661 15861 45695 15895
rect 28733 15657 28767 15691
rect 29101 15657 29135 15691
rect 31585 15657 31619 15691
rect 34897 15657 34931 15691
rect 35081 15657 35115 15691
rect 40233 15657 40267 15691
rect 41153 15657 41187 15691
rect 31401 15589 31435 15623
rect 36553 15589 36587 15623
rect 26985 15521 27019 15555
rect 31677 15521 31711 15555
rect 32413 15521 32447 15555
rect 32781 15521 32815 15555
rect 37473 15521 37507 15555
rect 38393 15521 38427 15555
rect 40325 15521 40359 15555
rect 43085 15521 43119 15555
rect 43913 15521 43947 15555
rect 46305 15521 46339 15555
rect 23397 15453 23431 15487
rect 23581 15453 23615 15487
rect 25605 15453 25639 15487
rect 26065 15453 26099 15487
rect 27169 15453 27203 15487
rect 27261 15453 27295 15487
rect 28917 15453 28951 15487
rect 29101 15453 29135 15487
rect 31953 15453 31987 15487
rect 32597 15453 32631 15487
rect 32873 15453 32907 15487
rect 33793 15453 33827 15487
rect 33977 15453 34011 15487
rect 34069 15453 34103 15487
rect 36461 15453 36495 15487
rect 36737 15453 36771 15487
rect 37565 15453 37599 15487
rect 37657 15453 37691 15487
rect 37749 15453 37783 15487
rect 40601 15453 40635 15487
rect 42533 15453 42567 15487
rect 43269 15453 43303 15487
rect 43821 15453 43855 15487
rect 45477 15453 45511 15487
rect 45569 15453 45603 15487
rect 45661 15453 45695 15487
rect 45845 15453 45879 15487
rect 27813 15385 27847 15419
rect 30481 15385 30515 15419
rect 30665 15385 30699 15419
rect 33609 15385 33643 15419
rect 35265 15385 35299 15419
rect 42625 15385 42659 15419
rect 45201 15385 45235 15419
rect 23489 15317 23523 15351
rect 26985 15317 27019 15351
rect 30297 15317 30331 15351
rect 35065 15317 35099 15351
rect 37289 15317 37323 15351
rect 40049 15317 40083 15351
rect 26065 15113 26099 15147
rect 31677 15113 31711 15147
rect 33057 15113 33091 15147
rect 33701 15113 33735 15147
rect 36737 15113 36771 15147
rect 44097 15113 44131 15147
rect 37565 15045 37599 15079
rect 38117 15045 38151 15079
rect 40969 15045 41003 15079
rect 42073 15045 42107 15079
rect 23949 14977 23983 15011
rect 24317 14977 24351 15011
rect 26065 14977 26099 15011
rect 26433 14977 26467 15011
rect 27353 14977 27387 15011
rect 27537 14977 27571 15011
rect 28181 14977 28215 15011
rect 28549 14977 28583 15011
rect 28825 14977 28859 15011
rect 28917 14977 28951 15011
rect 29837 14977 29871 15011
rect 30297 14977 30331 15011
rect 30481 14977 30515 15011
rect 31769 14977 31803 15011
rect 32561 14977 32595 15011
rect 32689 14977 32723 15011
rect 32873 14977 32907 15011
rect 33609 14977 33643 15011
rect 33793 14977 33827 15011
rect 35081 14977 35115 15011
rect 35265 14977 35299 15011
rect 35449 14977 35483 15011
rect 35633 14977 35667 15011
rect 36093 14977 36127 15011
rect 36277 14977 36311 15011
rect 36369 14977 36403 15011
rect 36461 14977 36495 15011
rect 38853 14977 38887 15011
rect 38945 14977 38979 15011
rect 39037 14977 39071 15011
rect 39221 14977 39255 15011
rect 39773 14977 39807 15011
rect 40049 14977 40083 15011
rect 40693 14977 40727 15011
rect 40785 14977 40819 15011
rect 41613 14977 41647 15011
rect 41797 14977 41831 15011
rect 41889 14977 41923 15011
rect 42717 14977 42751 15011
rect 42993 14977 43027 15011
rect 43177 14977 43211 15011
rect 44465 14977 44499 15011
rect 25881 14909 25915 14943
rect 27169 14909 27203 14943
rect 28365 14909 28399 14943
rect 35357 14909 35391 14943
rect 39865 14909 39899 14943
rect 39957 14909 39991 14943
rect 41981 14909 42015 14943
rect 43453 14909 43487 14943
rect 24225 14841 24259 14875
rect 30389 14841 30423 14875
rect 32777 14841 32811 14875
rect 38577 14841 38611 14875
rect 43361 14841 43395 14875
rect 43913 14841 43947 14875
rect 29653 14773 29687 14807
rect 34345 14773 34379 14807
rect 34897 14773 34931 14807
rect 40233 14773 40267 14807
rect 40969 14773 41003 14807
rect 44097 14773 44131 14807
rect 25329 14569 25363 14603
rect 26433 14569 26467 14603
rect 26985 14569 27019 14603
rect 27997 14569 28031 14603
rect 29193 14569 29227 14603
rect 30205 14569 30239 14603
rect 31401 14569 31435 14603
rect 34253 14569 34287 14603
rect 36921 14569 36955 14603
rect 39405 14569 39439 14603
rect 40049 14569 40083 14603
rect 42901 14569 42935 14603
rect 45293 14569 45327 14603
rect 32597 14501 32631 14535
rect 35449 14501 35483 14535
rect 28181 14433 28215 14467
rect 28273 14433 28307 14467
rect 30849 14433 30883 14467
rect 37933 14433 37967 14467
rect 38025 14433 38059 14467
rect 40693 14433 40727 14467
rect 42165 14433 42199 14467
rect 23857 14365 23891 14399
rect 25053 14365 25087 14399
rect 27537 14365 27571 14399
rect 28365 14365 28399 14399
rect 28457 14365 28491 14399
rect 30573 14365 30607 14399
rect 31401 14365 31435 14399
rect 31585 14365 31619 14399
rect 34069 14365 34103 14399
rect 34345 14365 34379 14399
rect 35633 14365 35667 14399
rect 35817 14365 35851 14399
rect 36001 14365 36035 14399
rect 36093 14365 36127 14399
rect 37013 14365 37047 14399
rect 37197 14365 37231 14399
rect 37841 14365 37875 14399
rect 38117 14365 38151 14399
rect 40877 14365 40911 14399
rect 41061 14365 41095 14399
rect 41521 14365 41555 14399
rect 41889 14365 41923 14399
rect 42901 14365 42935 14399
rect 43085 14365 43119 14399
rect 44373 14365 44407 14399
rect 44557 14365 44591 14399
rect 32781 14297 32815 14331
rect 32965 14297 32999 14331
rect 34897 14297 34931 14331
rect 35725 14297 35759 14331
rect 39037 14297 39071 14331
rect 39221 14297 39255 14331
rect 23765 14229 23799 14263
rect 25513 14229 25547 14263
rect 30665 14229 30699 14263
rect 33885 14229 33919 14263
rect 37657 14229 37691 14263
rect 44465 14229 44499 14263
rect 23489 14025 23523 14059
rect 26065 14025 26099 14059
rect 27813 14025 27847 14059
rect 29285 14025 29319 14059
rect 29653 14025 29687 14059
rect 31125 14025 31159 14059
rect 31217 14025 31251 14059
rect 32781 14025 32815 14059
rect 34345 14025 34379 14059
rect 36461 14025 36495 14059
rect 40969 14025 41003 14059
rect 22845 13957 22879 13991
rect 26157 13957 26191 13991
rect 28733 13957 28767 13991
rect 29745 13957 29779 13991
rect 31493 13957 31527 13991
rect 37749 13957 37783 13991
rect 38853 13957 38887 13991
rect 41705 13957 41739 13991
rect 42993 13957 43027 13991
rect 22753 13889 22787 13923
rect 22937 13889 22971 13923
rect 23397 13889 23431 13923
rect 23673 13889 23707 13923
rect 24409 13889 24443 13923
rect 24593 13889 24627 13923
rect 25329 13889 25363 13923
rect 25513 13889 25547 13923
rect 25605 13889 25639 13923
rect 26065 13889 26099 13923
rect 26341 13889 26375 13923
rect 27353 13889 27387 13923
rect 28365 13889 28399 13923
rect 28549 13889 28583 13923
rect 28825 13889 28859 13923
rect 30941 13889 30975 13923
rect 31309 13889 31343 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 34989 13889 35023 13923
rect 35081 13889 35115 13923
rect 35265 13889 35299 13923
rect 35357 13889 35391 13923
rect 36459 13889 36493 13923
rect 37933 13889 37967 13923
rect 38025 13889 38059 13923
rect 38761 13889 38795 13923
rect 39681 13889 39715 13923
rect 40693 13889 40727 13923
rect 40834 13889 40868 13923
rect 41061 13889 41095 13923
rect 41889 13889 41923 13923
rect 42625 13889 42659 13923
rect 42901 13889 42935 13923
rect 44097 13889 44131 13923
rect 44281 13889 44315 13923
rect 44373 13889 44407 13923
rect 44557 13889 44591 13923
rect 45017 13889 45051 13923
rect 45201 13889 45235 13923
rect 24317 13821 24351 13855
rect 25145 13821 25179 13855
rect 27445 13821 27479 13855
rect 29929 13821 29963 13855
rect 32965 13821 32999 13855
rect 33149 13821 33183 13855
rect 36921 13821 36955 13855
rect 44189 13821 44223 13855
rect 36829 13753 36863 13787
rect 45661 13753 45695 13787
rect 23857 13685 23891 13719
rect 27169 13685 27203 13719
rect 34805 13685 34839 13719
rect 36277 13685 36311 13719
rect 37749 13685 37783 13719
rect 39497 13685 39531 13719
rect 40693 13685 40727 13719
rect 41521 13685 41555 13719
rect 43913 13685 43947 13719
rect 45017 13685 45051 13719
rect 28917 13481 28951 13515
rect 29837 13481 29871 13515
rect 31033 13481 31067 13515
rect 32873 13481 32907 13515
rect 33609 13481 33643 13515
rect 33885 13481 33919 13515
rect 36461 13481 36495 13515
rect 38853 13481 38887 13515
rect 40693 13481 40727 13515
rect 41429 13481 41463 13515
rect 26801 13413 26835 13447
rect 30389 13413 30423 13447
rect 36829 13413 36863 13447
rect 37841 13413 37875 13447
rect 41981 13413 42015 13447
rect 43269 13413 43303 13447
rect 43361 13413 43395 13447
rect 44005 13413 44039 13447
rect 23765 13345 23799 13379
rect 25145 13345 25179 13379
rect 27261 13345 27295 13379
rect 27813 13345 27847 13379
rect 31769 13345 31803 13379
rect 34253 13345 34287 13379
rect 35173 13345 35207 13379
rect 36737 13345 36771 13379
rect 37933 13345 37967 13379
rect 41245 13345 41279 13379
rect 23397 13277 23431 13311
rect 23489 13277 23523 13311
rect 24777 13277 24811 13311
rect 25237 13277 25271 13311
rect 26065 13277 26099 13311
rect 26341 13277 26375 13311
rect 27169 13277 27203 13311
rect 27997 13277 28031 13311
rect 28365 13277 28399 13311
rect 29009 13277 29043 13311
rect 30297 13277 30331 13311
rect 30481 13277 30515 13311
rect 31309 13277 31343 13311
rect 32597 13277 32631 13311
rect 33793 13277 33827 13311
rect 34161 13277 34195 13311
rect 35081 13277 35115 13311
rect 35633 13277 35667 13311
rect 36645 13277 36679 13311
rect 36921 13277 36955 13311
rect 37565 13277 37599 13311
rect 37749 13277 37783 13311
rect 38025 13277 38059 13311
rect 38669 13277 38703 13311
rect 40325 13277 40359 13311
rect 40785 13277 40819 13311
rect 41521 13277 41555 13311
rect 42165 13277 42199 13311
rect 42257 13277 42291 13311
rect 42441 13277 42475 13311
rect 42533 13277 42567 13311
rect 42993 13277 43027 13311
rect 43177 13277 43211 13311
rect 43453 13277 43487 13311
rect 44005 13277 44039 13311
rect 44189 13277 44223 13311
rect 31033 13209 31067 13243
rect 32873 13209 32907 13243
rect 38780 13209 38814 13243
rect 38945 13209 38979 13243
rect 40417 13209 40451 13243
rect 41245 13209 41279 13243
rect 23581 13141 23615 13175
rect 23765 13141 23799 13175
rect 24869 13141 24903 13175
rect 24961 13141 24995 13175
rect 25421 13141 25455 13175
rect 25881 13141 25915 13175
rect 26249 13141 26283 13175
rect 28273 13141 28307 13175
rect 31217 13141 31251 13175
rect 32689 13141 32723 13175
rect 38209 13141 38243 13175
rect 40049 13141 40083 13175
rect 40509 13141 40543 13175
rect 25881 12937 25915 12971
rect 26049 12937 26083 12971
rect 28917 12937 28951 12971
rect 33885 12937 33919 12971
rect 34529 12937 34563 12971
rect 35449 12937 35483 12971
rect 36645 12937 36679 12971
rect 38301 12937 38335 12971
rect 41797 12937 41831 12971
rect 26249 12869 26283 12903
rect 27261 12869 27295 12903
rect 27477 12869 27511 12903
rect 30941 12869 30975 12903
rect 31125 12869 31159 12903
rect 40877 12869 40911 12903
rect 42625 12869 42659 12903
rect 23673 12801 23707 12835
rect 24317 12801 24351 12835
rect 28365 12801 28399 12835
rect 28917 12801 28951 12835
rect 29929 12801 29963 12835
rect 30757 12801 30791 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 32689 12801 32723 12835
rect 33701 12801 33735 12835
rect 34437 12801 34471 12835
rect 34713 12801 34747 12835
rect 35633 12801 35667 12835
rect 36553 12801 36587 12835
rect 36737 12801 36771 12835
rect 37657 12801 37691 12835
rect 37841 12801 37875 12835
rect 39405 12801 39439 12835
rect 39681 12801 39715 12835
rect 41061 12801 41095 12835
rect 41245 12801 41279 12835
rect 41337 12801 41371 12835
rect 28457 12733 28491 12767
rect 29852 12733 29886 12767
rect 30297 12733 30331 12767
rect 32597 12733 32631 12767
rect 35909 12733 35943 12767
rect 39221 12733 39255 12767
rect 39497 12733 39531 12767
rect 39589 12733 39623 12767
rect 27629 12665 27663 12699
rect 32321 12665 32355 12699
rect 35817 12665 35851 12699
rect 24961 12597 24995 12631
rect 26065 12597 26099 12631
rect 27445 12597 27479 12631
rect 29653 12597 29687 12631
rect 31585 12597 31619 12631
rect 34713 12597 34747 12631
rect 37657 12597 37691 12631
rect 28549 12393 28583 12427
rect 28917 12393 28951 12427
rect 30205 12393 30239 12427
rect 32597 12393 32631 12427
rect 35633 12393 35667 12427
rect 37013 12393 37047 12427
rect 40877 12393 40911 12427
rect 41705 12393 41739 12427
rect 26893 12325 26927 12359
rect 29837 12325 29871 12359
rect 36369 12325 36403 12359
rect 25053 12257 25087 12291
rect 27813 12257 27847 12291
rect 27905 12257 27939 12291
rect 28641 12257 28675 12291
rect 32045 12257 32079 12291
rect 32873 12257 32907 12291
rect 32965 12257 32999 12291
rect 33977 12257 34011 12291
rect 34069 12257 34103 12291
rect 36553 12257 36587 12291
rect 25237 12189 25271 12223
rect 25881 12189 25915 12223
rect 26157 12189 26191 12223
rect 27721 12189 27755 12223
rect 28549 12189 28583 12223
rect 29745 12189 29779 12223
rect 30021 12189 30055 12223
rect 30941 12189 30975 12223
rect 31125 12189 31159 12223
rect 31217 12189 31251 12223
rect 31309 12189 31343 12223
rect 32781 12189 32815 12223
rect 33057 12189 33091 12223
rect 33885 12189 33919 12223
rect 34161 12189 34195 12223
rect 35449 12189 35483 12223
rect 35541 12189 35575 12223
rect 36277 12189 36311 12223
rect 37749 12189 37783 12223
rect 25421 12053 25455 12087
rect 27353 12053 27387 12087
rect 31585 12053 31619 12087
rect 34345 12053 34379 12087
rect 35817 12053 35851 12087
rect 36553 12053 36587 12087
rect 37657 12053 37691 12087
rect 25697 11849 25731 11883
rect 26157 11849 26191 11883
rect 27629 11849 27663 11883
rect 28825 11849 28859 11883
rect 30481 11849 30515 11883
rect 31125 11849 31159 11883
rect 31493 11849 31527 11883
rect 32781 11849 32815 11883
rect 33517 11849 33551 11883
rect 32597 11781 32631 11815
rect 34437 11781 34471 11815
rect 34621 11781 34655 11815
rect 35541 11781 35575 11815
rect 35757 11781 35791 11815
rect 1869 11713 1903 11747
rect 2421 11713 2455 11747
rect 25513 11713 25547 11747
rect 26341 11713 26375 11747
rect 27537 11713 27571 11747
rect 29009 11713 29043 11747
rect 30481 11713 30515 11747
rect 30665 11713 30699 11747
rect 31309 11713 31343 11747
rect 31585 11713 31619 11747
rect 32873 11713 32907 11747
rect 33333 11713 33367 11747
rect 36737 11713 36771 11747
rect 37841 11713 37875 11747
rect 38209 11713 38243 11747
rect 38485 11713 38519 11747
rect 38853 11713 38887 11747
rect 39313 11713 39347 11747
rect 25053 11645 25087 11679
rect 27813 11645 27847 11679
rect 29193 11645 29227 11679
rect 36645 11645 36679 11679
rect 38025 11645 38059 11679
rect 1685 11577 1719 11611
rect 27169 11577 27203 11611
rect 30021 11577 30055 11611
rect 32597 11577 32631 11611
rect 34805 11509 34839 11543
rect 35725 11509 35759 11543
rect 35909 11509 35943 11543
rect 36369 11509 36403 11543
rect 39405 11509 39439 11543
rect 39773 11509 39807 11543
rect 25697 11305 25731 11339
rect 27445 11305 27479 11339
rect 29929 11305 29963 11339
rect 30481 11305 30515 11339
rect 32965 11305 32999 11339
rect 34989 11305 35023 11339
rect 36185 11305 36219 11339
rect 36829 11305 36863 11339
rect 58173 11305 58207 11339
rect 26249 11237 26283 11271
rect 39129 11237 39163 11271
rect 28549 11169 28583 11203
rect 32413 11169 32447 11203
rect 33885 11169 33919 11203
rect 37013 11169 37047 11203
rect 37105 11169 37139 11203
rect 28641 11101 28675 11135
rect 29745 11101 29779 11135
rect 29929 11101 29963 11135
rect 32137 11101 32171 11135
rect 32229 11101 32263 11135
rect 33609 11101 33643 11135
rect 33701 11101 33735 11135
rect 35081 11101 35115 11135
rect 35541 11101 35575 11135
rect 35725 11101 35759 11135
rect 37197 11101 37231 11135
rect 37289 11101 37323 11135
rect 37841 11101 37875 11135
rect 26893 11033 26927 11067
rect 33885 11033 33919 11067
rect 35633 11033 35667 11067
rect 57621 11033 57655 11067
rect 58265 11033 58299 11067
rect 27997 10965 28031 10999
rect 29009 10965 29043 10999
rect 32413 10965 32447 10999
rect 28917 10761 28951 10795
rect 32321 10761 32355 10795
rect 32489 10761 32523 10795
rect 33149 10761 33183 10795
rect 35449 10761 35483 10795
rect 37473 10761 37507 10795
rect 27445 10693 27479 10727
rect 30021 10693 30055 10727
rect 32689 10693 32723 10727
rect 36277 10693 36311 10727
rect 36461 10693 36495 10727
rect 39497 10693 39531 10727
rect 27169 10625 27203 10659
rect 31769 10625 31803 10659
rect 33333 10625 33367 10659
rect 33517 10625 33551 10659
rect 34621 10625 34655 10659
rect 35357 10625 35391 10659
rect 35541 10625 35575 10659
rect 29745 10557 29779 10591
rect 34437 10557 34471 10591
rect 34713 10557 34747 10591
rect 34805 10557 34839 10591
rect 39129 10489 39163 10523
rect 26433 10421 26467 10455
rect 32505 10421 32539 10455
rect 33333 10421 33367 10455
rect 36093 10421 36127 10455
rect 39037 10421 39071 10455
rect 26893 10217 26927 10251
rect 29101 10217 29135 10251
rect 31309 10217 31343 10251
rect 33241 10217 33275 10251
rect 33885 10217 33919 10251
rect 27445 10149 27479 10183
rect 36829 10149 36863 10183
rect 29837 10081 29871 10115
rect 30297 10081 30331 10115
rect 36093 10081 36127 10115
rect 37289 10081 37323 10115
rect 40141 10081 40175 10115
rect 27905 10013 27939 10047
rect 28089 10013 28123 10047
rect 29929 10013 29963 10047
rect 31217 10013 31251 10047
rect 33885 10013 33919 10047
rect 34069 10013 34103 10047
rect 36001 10013 36035 10047
rect 37197 10013 37231 10047
rect 38301 10013 38335 10047
rect 38577 10013 38611 10047
rect 38761 10013 38795 10047
rect 40233 10013 40267 10047
rect 27905 9877 27939 9911
rect 28641 9877 28675 9911
rect 33701 9877 33735 9911
rect 35633 9877 35667 9911
rect 38117 9877 38151 9911
rect 40601 9877 40635 9911
rect 28917 9673 28951 9707
rect 29653 9605 29687 9639
rect 29837 9605 29871 9639
rect 32505 9605 32539 9639
rect 33057 9605 33091 9639
rect 37657 9605 37691 9639
rect 26617 9537 26651 9571
rect 27169 9537 27203 9571
rect 31033 9537 31067 9571
rect 33701 9537 33735 9571
rect 33885 9537 33919 9571
rect 33977 9537 34011 9571
rect 34437 9537 34471 9571
rect 34897 9537 34931 9571
rect 35081 9537 35115 9571
rect 35541 9537 35575 9571
rect 35725 9537 35759 9571
rect 36921 9537 36955 9571
rect 37473 9537 37507 9571
rect 37749 9537 37783 9571
rect 38577 9537 38611 9571
rect 27445 9469 27479 9503
rect 30573 9469 30607 9503
rect 31125 9469 31159 9503
rect 38485 9469 38519 9503
rect 38945 9469 38979 9503
rect 34345 9401 34379 9435
rect 37473 9401 37507 9435
rect 30021 9333 30055 9367
rect 31125 9333 31159 9367
rect 31401 9333 31435 9367
rect 35081 9333 35115 9367
rect 35633 9333 35667 9367
rect 27169 9129 27203 9163
rect 28273 9129 28307 9163
rect 29101 9129 29135 9163
rect 30849 9129 30883 9163
rect 31401 9129 31435 9163
rect 32965 9129 32999 9163
rect 29837 9061 29871 9095
rect 34253 9061 34287 9095
rect 31585 8993 31619 9027
rect 32873 8993 32907 9027
rect 35633 8993 35667 9027
rect 26617 8925 26651 8959
rect 27077 8925 27111 8959
rect 27261 8925 27295 8959
rect 30021 8925 30055 8959
rect 30665 8925 30699 8959
rect 30941 8925 30975 8959
rect 31677 8925 31711 8959
rect 31769 8925 31803 8959
rect 32597 8925 32631 8959
rect 33885 8925 33919 8959
rect 33977 8925 34011 8959
rect 34069 8925 34103 8959
rect 35541 8925 35575 8959
rect 37657 8925 37691 8959
rect 38025 8925 38059 8959
rect 27997 8857 28031 8891
rect 33701 8857 33735 8891
rect 39497 8857 39531 8891
rect 30481 8789 30515 8823
rect 33149 8789 33183 8823
rect 35909 8789 35943 8823
rect 27905 8585 27939 8619
rect 30205 8585 30239 8619
rect 31125 8585 31159 8619
rect 32689 8585 32723 8619
rect 33793 8585 33827 8619
rect 35081 8585 35115 8619
rect 38025 8517 38059 8551
rect 28457 8449 28491 8483
rect 30941 8449 30975 8483
rect 31217 8449 31251 8483
rect 32505 8449 32539 8483
rect 32781 8449 32815 8483
rect 32965 8449 32999 8483
rect 33609 8449 33643 8483
rect 33885 8449 33919 8483
rect 34897 8449 34931 8483
rect 35173 8449 35207 8483
rect 35909 8449 35943 8483
rect 36093 8449 36127 8483
rect 28733 8381 28767 8415
rect 30757 8381 30791 8415
rect 34713 8381 34747 8415
rect 36921 8381 36955 8415
rect 27353 8313 27387 8347
rect 37749 8313 37783 8347
rect 33425 8245 33459 8279
rect 37565 8245 37599 8279
rect 28181 8041 28215 8075
rect 30389 8041 30423 8075
rect 33977 8041 34011 8075
rect 31401 7973 31435 8007
rect 31033 7905 31067 7939
rect 32873 7837 32907 7871
rect 33057 7837 33091 7871
rect 33241 7837 33275 7871
rect 33333 7837 33367 7871
rect 33961 7769 33995 7803
rect 34161 7769 34195 7803
rect 31493 7701 31527 7735
rect 33793 7701 33827 7735
rect 31401 7361 31435 7395
rect 33701 7361 33735 7395
rect 31309 7293 31343 7327
rect 33793 7293 33827 7327
rect 33333 7225 33367 7259
rect 31769 7157 31803 7191
rect 33701 6953 33735 6987
rect 33517 6885 33551 6919
rect 33241 6749 33275 6783
rect 57529 5865 57563 5899
rect 1869 5661 1903 5695
rect 2421 5661 2455 5695
rect 58081 5661 58115 5695
rect 1685 5525 1719 5559
rect 58265 5525 58299 5559
rect 27997 2601 28031 2635
rect 37565 2601 37599 2635
rect 44097 2601 44131 2635
rect 5733 2465 5767 2499
rect 17693 2465 17727 2499
rect 57437 2465 57471 2499
rect 1869 2397 1903 2431
rect 6009 2397 6043 2431
rect 6561 2397 6595 2431
rect 11989 2397 12023 2431
rect 17141 2397 17175 2431
rect 22293 2397 22327 2431
rect 27445 2397 27479 2431
rect 32965 2397 32999 2431
rect 38117 2397 38151 2431
rect 43453 2397 43487 2431
rect 43913 2397 43947 2431
rect 48513 2397 48547 2431
rect 49065 2397 49099 2431
rect 55505 2397 55539 2431
rect 58081 2397 58115 2431
rect 2421 2329 2455 2363
rect 12541 2329 12575 2363
rect 54861 2329 54895 2363
rect 1685 2261 1719 2295
rect 11805 2261 11839 2295
rect 16957 2261 16991 2295
rect 22109 2261 22143 2295
rect 27261 2261 27295 2295
rect 33149 2261 33183 2295
rect 38301 2261 38335 2295
rect 49249 2261 49283 2295
rect 55689 2261 55723 2295
rect 58265 2261 58299 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1670 57576 1676 57588
rect 1631 57548 1676 57576
rect 1670 57536 1676 57548
rect 1728 57536 1734 57588
rect 8386 57536 8392 57588
rect 8444 57576 8450 57588
rect 9217 57579 9275 57585
rect 9217 57576 9229 57579
rect 8444 57548 9229 57576
rect 8444 57536 8450 57548
rect 9217 57545 9229 57548
rect 9263 57545 9275 57579
rect 9217 57539 9275 57545
rect 13538 57536 13544 57588
rect 13596 57576 13602 57588
rect 14461 57579 14519 57585
rect 14461 57576 14473 57579
rect 13596 57548 14473 57576
rect 13596 57536 13602 57548
rect 14461 57545 14473 57548
rect 14507 57545 14519 57579
rect 14461 57539 14519 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19521 57579 19579 57585
rect 19521 57576 19533 57579
rect 19392 57548 19533 57576
rect 19392 57536 19398 57548
rect 19521 57545 19533 57548
rect 19567 57545 19579 57579
rect 19521 57539 19579 57545
rect 24486 57536 24492 57588
rect 24544 57576 24550 57588
rect 24673 57579 24731 57585
rect 24673 57576 24685 57579
rect 24544 57548 24685 57576
rect 24544 57536 24550 57548
rect 24673 57545 24685 57548
rect 24719 57545 24731 57579
rect 24673 57539 24731 57545
rect 35434 57536 35440 57588
rect 35492 57576 35498 57588
rect 35713 57579 35771 57585
rect 35713 57576 35725 57579
rect 35492 57548 35725 57576
rect 35492 57536 35498 57548
rect 35713 57545 35725 57548
rect 35759 57545 35771 57579
rect 35713 57539 35771 57545
rect 41414 57536 41420 57588
rect 41472 57576 41478 57588
rect 41509 57579 41567 57585
rect 41509 57576 41521 57579
rect 41472 57548 41521 57576
rect 41472 57536 41478 57548
rect 41509 57545 41521 57548
rect 41555 57545 41567 57579
rect 41509 57539 41567 57545
rect 46382 57536 46388 57588
rect 46440 57576 46446 57588
rect 46661 57579 46719 57585
rect 46661 57576 46673 57579
rect 46440 57548 46673 57576
rect 46440 57536 46446 57548
rect 46661 57545 46673 57548
rect 46707 57545 46719 57579
rect 46661 57539 46719 57545
rect 52178 57536 52184 57588
rect 52236 57576 52242 57588
rect 53101 57579 53159 57585
rect 53101 57576 53113 57579
rect 52236 57548 53113 57576
rect 52236 57536 52242 57548
rect 53101 57545 53113 57548
rect 53147 57545 53159 57579
rect 53101 57539 53159 57545
rect 57330 57536 57336 57588
rect 57388 57576 57394 57588
rect 58253 57579 58311 57585
rect 58253 57576 58265 57579
rect 57388 57548 58265 57576
rect 57388 57536 57394 57548
rect 58253 57545 58265 57548
rect 58299 57545 58311 57579
rect 58253 57539 58311 57545
rect 2590 57468 2596 57520
rect 2648 57508 2654 57520
rect 2777 57511 2835 57517
rect 2777 57508 2789 57511
rect 2648 57480 2789 57508
rect 2648 57468 2654 57480
rect 2777 57477 2789 57480
rect 2823 57477 2835 57511
rect 2777 57471 2835 57477
rect 29917 57511 29975 57517
rect 29917 57477 29929 57511
rect 29963 57508 29975 57511
rect 30282 57508 30288 57520
rect 29963 57480 30288 57508
rect 29963 57477 29975 57480
rect 29917 57471 29975 57477
rect 30282 57468 30288 57480
rect 30340 57508 30346 57520
rect 30469 57511 30527 57517
rect 30469 57508 30481 57511
rect 30340 57480 30481 57508
rect 30340 57468 30346 57480
rect 30469 57477 30481 57480
rect 30515 57477 30527 57511
rect 30469 57471 30527 57477
rect 1854 57440 1860 57452
rect 1815 57412 1860 57440
rect 1854 57400 1860 57412
rect 1912 57400 1918 57452
rect 9401 57443 9459 57449
rect 9401 57409 9413 57443
rect 9447 57440 9459 57443
rect 9858 57440 9864 57452
rect 9447 57412 9864 57440
rect 9447 57409 9459 57412
rect 9401 57403 9459 57409
rect 9858 57400 9864 57412
rect 9916 57400 9922 57452
rect 13725 57443 13783 57449
rect 13725 57409 13737 57443
rect 13771 57440 13783 57443
rect 14274 57440 14280 57452
rect 13771 57412 14280 57440
rect 13771 57409 13783 57412
rect 13725 57403 13783 57409
rect 14274 57400 14280 57412
rect 14332 57400 14338 57452
rect 19705 57443 19763 57449
rect 19705 57409 19717 57443
rect 19751 57409 19763 57443
rect 19705 57403 19763 57409
rect 24857 57443 24915 57449
rect 24857 57409 24869 57443
rect 24903 57440 24915 57443
rect 25314 57440 25320 57452
rect 24903 57412 25320 57440
rect 24903 57409 24915 57412
rect 24857 57403 24915 57409
rect 19720 57372 19748 57403
rect 25314 57400 25320 57412
rect 25372 57400 25378 57452
rect 35526 57440 35532 57452
rect 35487 57412 35532 57440
rect 35526 57400 35532 57412
rect 35584 57400 35590 57452
rect 40865 57443 40923 57449
rect 40865 57409 40877 57443
rect 40911 57440 40923 57443
rect 41322 57440 41328 57452
rect 40911 57412 41328 57440
rect 40911 57409 40923 57412
rect 40865 57403 40923 57409
rect 41322 57400 41328 57412
rect 41380 57400 41386 57452
rect 46017 57443 46075 57449
rect 46017 57409 46029 57443
rect 46063 57440 46075 57443
rect 46474 57440 46480 57452
rect 46063 57412 46480 57440
rect 46063 57409 46075 57412
rect 46017 57403 46075 57409
rect 46474 57400 46480 57412
rect 46532 57400 46538 57452
rect 52270 57400 52276 57452
rect 52328 57440 52334 57452
rect 52917 57443 52975 57449
rect 52917 57440 52929 57443
rect 52328 57412 52929 57440
rect 52328 57400 52334 57412
rect 52917 57409 52929 57412
rect 52963 57409 52975 57443
rect 58069 57443 58127 57449
rect 58069 57440 58081 57443
rect 52917 57403 52975 57409
rect 57440 57412 58081 57440
rect 20257 57375 20315 57381
rect 20257 57372 20269 57375
rect 19720 57344 20269 57372
rect 20257 57341 20269 57344
rect 20303 57372 20315 57375
rect 32398 57372 32404 57384
rect 20303 57344 32404 57372
rect 20303 57341 20315 57344
rect 20257 57335 20315 57341
rect 32398 57332 32404 57344
rect 32456 57332 32462 57384
rect 2866 57236 2872 57248
rect 2827 57208 2872 57236
rect 2866 57196 2872 57208
rect 2924 57196 2930 57248
rect 9858 57236 9864 57248
rect 9819 57208 9864 57236
rect 9858 57196 9864 57208
rect 9916 57196 9922 57248
rect 25314 57236 25320 57248
rect 25275 57208 25320 57236
rect 25314 57196 25320 57208
rect 25372 57196 25378 57248
rect 30558 57236 30564 57248
rect 30519 57208 30564 57236
rect 30558 57196 30564 57208
rect 30616 57196 30622 57248
rect 52270 57236 52276 57248
rect 52231 57208 52276 57236
rect 52270 57196 52276 57208
rect 52328 57196 52334 57248
rect 57146 57196 57152 57248
rect 57204 57236 57210 57248
rect 57440 57245 57468 57412
rect 58069 57409 58081 57412
rect 58115 57409 58127 57443
rect 58069 57403 58127 57409
rect 57425 57239 57483 57245
rect 57425 57236 57437 57239
rect 57204 57208 57437 57236
rect 57204 57196 57210 57208
rect 57425 57205 57437 57208
rect 57471 57205 57483 57239
rect 57425 57199 57483 57205
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 2590 57032 2596 57044
rect 2551 57004 2596 57032
rect 2590 56992 2596 57004
rect 2648 56992 2654 57044
rect 35253 57035 35311 57041
rect 35253 57001 35265 57035
rect 35299 57032 35311 57035
rect 35526 57032 35532 57044
rect 35299 57004 35532 57032
rect 35299 57001 35311 57004
rect 35253 56995 35311 57001
rect 35526 56992 35532 57004
rect 35584 56992 35590 57044
rect 58250 57032 58256 57044
rect 58211 57004 58256 57032
rect 58250 56992 58256 57004
rect 58308 56992 58314 57044
rect 35069 56831 35127 56837
rect 35069 56797 35081 56831
rect 35115 56828 35127 56831
rect 58069 56831 58127 56837
rect 58069 56828 58081 56831
rect 35115 56800 35664 56828
rect 35115 56797 35127 56800
rect 35069 56791 35127 56797
rect 35636 56704 35664 56800
rect 57624 56800 58081 56828
rect 57624 56704 57652 56800
rect 58069 56797 58081 56800
rect 58115 56797 58127 56831
rect 58069 56791 58127 56797
rect 1854 56652 1860 56704
rect 1912 56692 1918 56704
rect 1949 56695 2007 56701
rect 1949 56692 1961 56695
rect 1912 56664 1961 56692
rect 1912 56652 1918 56664
rect 1949 56661 1961 56664
rect 1995 56661 2007 56695
rect 1949 56655 2007 56661
rect 35618 56652 35624 56704
rect 35676 56692 35682 56704
rect 35713 56695 35771 56701
rect 35713 56692 35725 56695
rect 35676 56664 35725 56692
rect 35676 56652 35682 56664
rect 35713 56661 35725 56664
rect 35759 56661 35771 56695
rect 57606 56692 57612 56704
rect 57567 56664 57612 56692
rect 35713 56655 35771 56661
rect 57606 56652 57612 56664
rect 57664 56652 57670 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1857 52003 1915 52009
rect 1857 51969 1869 52003
rect 1903 52000 1915 52003
rect 2130 52000 2136 52012
rect 1903 51972 2136 52000
rect 1903 51969 1915 51972
rect 1857 51963 1915 51969
rect 2130 51960 2136 51972
rect 2188 51960 2194 52012
rect 58069 52003 58127 52009
rect 58069 52000 58081 52003
rect 57440 51972 58081 52000
rect 1670 51796 1676 51808
rect 1631 51768 1676 51796
rect 1670 51756 1676 51768
rect 1728 51756 1734 51808
rect 2130 51756 2136 51808
rect 2188 51796 2194 51808
rect 2317 51799 2375 51805
rect 2317 51796 2329 51799
rect 2188 51768 2329 51796
rect 2188 51756 2194 51768
rect 2317 51765 2329 51768
rect 2363 51765 2375 51799
rect 2317 51759 2375 51765
rect 57238 51756 57244 51808
rect 57296 51796 57302 51808
rect 57440 51805 57468 51972
rect 58069 51969 58081 51972
rect 58115 51969 58127 52003
rect 58069 51963 58127 51969
rect 57425 51799 57483 51805
rect 57425 51796 57437 51799
rect 57296 51768 57437 51796
rect 57296 51756 57302 51768
rect 57425 51765 57437 51768
rect 57471 51765 57483 51799
rect 58250 51796 58256 51808
rect 58211 51768 58256 51796
rect 57425 51759 57483 51765
rect 58250 51756 58256 51768
rect 58308 51756 58314 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 29730 47988 29736 48000
rect 29691 47960 29736 47988
rect 29730 47948 29736 47960
rect 29788 47948 29794 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 25958 47744 25964 47796
rect 26016 47784 26022 47796
rect 26016 47756 31754 47784
rect 26016 47744 26022 47756
rect 31726 47728 31754 47756
rect 25041 47719 25099 47725
rect 25041 47685 25053 47719
rect 25087 47716 25099 47719
rect 27246 47716 27252 47728
rect 25087 47688 27252 47716
rect 25087 47685 25099 47688
rect 25041 47679 25099 47685
rect 27246 47676 27252 47688
rect 27304 47716 27310 47728
rect 27304 47688 28764 47716
rect 31726 47688 31760 47728
rect 27304 47676 27310 47688
rect 28258 47648 28264 47660
rect 28219 47620 28264 47648
rect 28258 47608 28264 47620
rect 28316 47608 28322 47660
rect 28442 47648 28448 47660
rect 28403 47620 28448 47648
rect 28442 47608 28448 47620
rect 28500 47608 28506 47660
rect 28736 47657 28764 47688
rect 31754 47676 31760 47688
rect 31812 47676 31818 47728
rect 28721 47651 28779 47657
rect 28721 47617 28733 47651
rect 28767 47617 28779 47651
rect 28721 47611 28779 47617
rect 32582 47608 32588 47660
rect 32640 47648 32646 47660
rect 33413 47651 33471 47657
rect 33413 47648 33425 47651
rect 32640 47620 33425 47648
rect 32640 47608 32646 47620
rect 33413 47617 33425 47620
rect 33459 47648 33471 47651
rect 33459 47620 34008 47648
rect 33459 47617 33471 47620
rect 33413 47611 33471 47617
rect 25593 47583 25651 47589
rect 25593 47580 25605 47583
rect 23676 47552 25605 47580
rect 22370 47444 22376 47456
rect 22331 47416 22376 47444
rect 22370 47404 22376 47416
rect 22428 47404 22434 47456
rect 23017 47447 23075 47453
rect 23017 47413 23029 47447
rect 23063 47444 23075 47447
rect 23198 47444 23204 47456
rect 23063 47416 23204 47444
rect 23063 47413 23075 47416
rect 23017 47407 23075 47413
rect 23198 47404 23204 47416
rect 23256 47444 23262 47456
rect 23676 47453 23704 47552
rect 25593 47549 25605 47552
rect 25639 47549 25651 47583
rect 25593 47543 25651 47549
rect 25774 47540 25780 47592
rect 25832 47580 25838 47592
rect 29273 47583 29331 47589
rect 29273 47580 29285 47583
rect 25832 47552 29285 47580
rect 25832 47540 25838 47552
rect 29273 47549 29285 47552
rect 29319 47580 29331 47583
rect 29362 47580 29368 47592
rect 29319 47552 29368 47580
rect 29319 47549 29331 47552
rect 29273 47543 29331 47549
rect 29362 47540 29368 47552
rect 29420 47540 29426 47592
rect 33226 47580 33232 47592
rect 33187 47552 33232 47580
rect 33226 47540 33232 47552
rect 33284 47540 33290 47592
rect 31018 47512 31024 47524
rect 24964 47484 31024 47512
rect 23661 47447 23719 47453
rect 23661 47444 23673 47447
rect 23256 47416 23673 47444
rect 23256 47404 23262 47416
rect 23661 47413 23673 47416
rect 23707 47413 23719 47447
rect 23661 47407 23719 47413
rect 24670 47404 24676 47456
rect 24728 47444 24734 47456
rect 24964 47453 24992 47484
rect 31018 47472 31024 47484
rect 31076 47472 31082 47524
rect 24949 47447 25007 47453
rect 24949 47444 24961 47447
rect 24728 47416 24961 47444
rect 24728 47404 24734 47416
rect 24949 47413 24961 47416
rect 24995 47413 25007 47447
rect 24949 47407 25007 47413
rect 29730 47404 29736 47456
rect 29788 47444 29794 47456
rect 30285 47447 30343 47453
rect 30285 47444 30297 47447
rect 29788 47416 30297 47444
rect 29788 47404 29794 47416
rect 30285 47413 30297 47416
rect 30331 47413 30343 47447
rect 31294 47444 31300 47456
rect 31255 47416 31300 47444
rect 30285 47407 30343 47413
rect 31294 47404 31300 47416
rect 31352 47404 31358 47456
rect 33980 47453 34008 47620
rect 33965 47447 34023 47453
rect 33965 47413 33977 47447
rect 34011 47444 34023 47447
rect 34422 47444 34428 47456
rect 34011 47416 34428 47444
rect 34011 47413 34023 47416
rect 33965 47407 34023 47413
rect 34422 47404 34428 47416
rect 34480 47404 34486 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 28721 47243 28779 47249
rect 28721 47209 28733 47243
rect 28767 47209 28779 47243
rect 32582 47240 32588 47252
rect 32543 47212 32588 47240
rect 28721 47203 28779 47209
rect 25222 47132 25228 47184
rect 25280 47172 25286 47184
rect 26697 47175 26755 47181
rect 26697 47172 26709 47175
rect 25280 47144 26709 47172
rect 25280 47132 25286 47144
rect 26697 47141 26709 47144
rect 26743 47172 26755 47175
rect 26970 47172 26976 47184
rect 26743 47144 26976 47172
rect 26743 47141 26755 47144
rect 26697 47135 26755 47141
rect 26970 47132 26976 47144
rect 27028 47132 27034 47184
rect 27893 47175 27951 47181
rect 27893 47141 27905 47175
rect 27939 47172 27951 47175
rect 28626 47172 28632 47184
rect 27939 47144 28632 47172
rect 27939 47141 27951 47144
rect 27893 47135 27951 47141
rect 28626 47132 28632 47144
rect 28684 47132 28690 47184
rect 21266 47064 21272 47116
rect 21324 47104 21330 47116
rect 23201 47107 23259 47113
rect 23201 47104 23213 47107
rect 21324 47076 23213 47104
rect 21324 47064 21330 47076
rect 22020 47045 22048 47076
rect 23201 47073 23213 47076
rect 23247 47073 23259 47107
rect 25958 47104 25964 47116
rect 23201 47067 23259 47073
rect 23400 47076 25964 47104
rect 22005 47039 22063 47045
rect 22005 47005 22017 47039
rect 22051 47036 22063 47039
rect 22189 47039 22247 47045
rect 22051 47008 22085 47036
rect 22051 47005 22063 47008
rect 22005 46999 22063 47005
rect 22189 47005 22201 47039
rect 22235 47036 22247 47039
rect 23014 47036 23020 47048
rect 22235 47008 22876 47036
rect 22975 47008 23020 47036
rect 22235 47005 22247 47008
rect 22189 46999 22247 47005
rect 22094 46928 22100 46980
rect 22152 46968 22158 46980
rect 22848 46968 22876 47008
rect 23014 46996 23020 47008
rect 23072 46996 23078 47048
rect 23400 47036 23428 47076
rect 25958 47064 25964 47076
rect 26016 47064 26022 47116
rect 26988 47104 27016 47132
rect 28736 47104 28764 47203
rect 32582 47200 32588 47212
rect 32640 47200 32646 47252
rect 28902 47104 28908 47116
rect 26988 47076 28908 47104
rect 23124 47008 23428 47036
rect 23477 47039 23535 47045
rect 23124 46968 23152 47008
rect 23477 47005 23489 47039
rect 23523 47036 23535 47039
rect 24762 47036 24768 47048
rect 23523 47008 24768 47036
rect 23523 47005 23535 47008
rect 23477 46999 23535 47005
rect 24762 46996 24768 47008
rect 24820 47036 24826 47048
rect 24857 47039 24915 47045
rect 24857 47036 24869 47039
rect 24820 47008 24869 47036
rect 24820 46996 24826 47008
rect 24857 47005 24869 47008
rect 24903 47005 24915 47039
rect 25130 47036 25136 47048
rect 25091 47008 25136 47036
rect 24857 46999 24915 47005
rect 25130 46996 25136 47008
rect 25188 46996 25194 47048
rect 26510 47036 26516 47048
rect 26471 47008 26516 47036
rect 26510 46996 26516 47008
rect 26568 46996 26574 47048
rect 26786 47036 26792 47048
rect 26747 47008 26792 47036
rect 26786 46996 26792 47008
rect 26844 47036 26850 47048
rect 27908 47045 27936 47076
rect 28902 47064 28908 47076
rect 28960 47064 28966 47116
rect 31754 47064 31760 47116
rect 31812 47104 31818 47116
rect 31812 47076 31857 47104
rect 31812 47064 31818 47076
rect 27709 47039 27767 47045
rect 27709 47036 27721 47039
rect 26844 47008 27721 47036
rect 26844 46996 26850 47008
rect 27709 47005 27721 47008
rect 27755 47005 27767 47039
rect 27709 46999 27767 47005
rect 27893 47039 27951 47045
rect 27893 47005 27905 47039
rect 27939 47005 27951 47039
rect 27893 46999 27951 47005
rect 22152 46940 22197 46968
rect 22848 46940 23152 46968
rect 23385 46971 23443 46977
rect 22152 46928 22158 46940
rect 23385 46937 23397 46971
rect 23431 46968 23443 46971
rect 24670 46968 24676 46980
rect 23431 46940 24676 46968
rect 23431 46937 23443 46940
rect 23385 46931 23443 46937
rect 24670 46928 24676 46940
rect 24728 46968 24734 46980
rect 24949 46971 25007 46977
rect 24949 46968 24961 46971
rect 24728 46940 24961 46968
rect 24728 46928 24734 46940
rect 24949 46937 24961 46940
rect 24995 46937 25007 46971
rect 25774 46968 25780 46980
rect 24949 46931 25007 46937
rect 25148 46940 25780 46968
rect 23290 46860 23296 46912
rect 23348 46900 23354 46912
rect 23937 46903 23995 46909
rect 23937 46900 23949 46903
rect 23348 46872 23949 46900
rect 23348 46860 23354 46872
rect 23937 46869 23949 46872
rect 23983 46900 23995 46903
rect 25148 46900 25176 46940
rect 25774 46928 25780 46940
rect 25832 46928 25838 46980
rect 26528 46968 26556 46996
rect 27525 46971 27583 46977
rect 27525 46968 27537 46971
rect 26528 46940 27537 46968
rect 27525 46937 27537 46940
rect 27571 46937 27583 46971
rect 27724 46968 27752 46999
rect 28534 46996 28540 47048
rect 28592 47036 28598 47048
rect 29089 47039 29147 47045
rect 29089 47036 29101 47039
rect 28592 47008 29101 47036
rect 28592 46996 28598 47008
rect 29089 47005 29101 47008
rect 29135 47005 29147 47039
rect 30837 47039 30895 47045
rect 30837 47036 30849 47039
rect 29089 46999 29147 47005
rect 29380 47008 30849 47036
rect 29380 46968 29408 47008
rect 30837 47005 30849 47008
rect 30883 47036 30895 47039
rect 30926 47036 30932 47048
rect 30883 47008 30932 47036
rect 30883 47005 30895 47008
rect 30837 46999 30895 47005
rect 30926 46996 30932 47008
rect 30984 46996 30990 47048
rect 31018 46996 31024 47048
rect 31076 47036 31082 47048
rect 31076 47008 31121 47036
rect 31076 46996 31082 47008
rect 27724 46940 29408 46968
rect 27525 46931 27583 46937
rect 30098 46928 30104 46980
rect 30156 46968 30162 46980
rect 30285 46971 30343 46977
rect 30285 46968 30297 46971
rect 30156 46940 30297 46968
rect 30156 46928 30162 46940
rect 30285 46937 30297 46940
rect 30331 46968 30343 46971
rect 31294 46968 31300 46980
rect 30331 46940 31300 46968
rect 30331 46937 30343 46940
rect 30285 46931 30343 46937
rect 31294 46928 31300 46940
rect 31352 46928 31358 46980
rect 33413 46971 33471 46977
rect 33413 46937 33425 46971
rect 33459 46968 33471 46971
rect 33594 46968 33600 46980
rect 33459 46940 33600 46968
rect 33459 46937 33471 46940
rect 33413 46931 33471 46937
rect 33594 46928 33600 46940
rect 33652 46928 33658 46980
rect 25314 46900 25320 46912
rect 23983 46872 25176 46900
rect 25275 46872 25320 46900
rect 23983 46869 23995 46872
rect 23937 46863 23995 46869
rect 25314 46860 25320 46872
rect 25372 46860 25378 46912
rect 25869 46903 25927 46909
rect 25869 46869 25881 46903
rect 25915 46900 25927 46903
rect 26050 46900 26056 46912
rect 25915 46872 26056 46900
rect 25915 46869 25927 46872
rect 25869 46863 25927 46869
rect 26050 46860 26056 46872
rect 26108 46860 26114 46912
rect 26326 46900 26332 46912
rect 26287 46872 26332 46900
rect 26326 46860 26332 46872
rect 26384 46860 26390 46912
rect 27614 46860 27620 46912
rect 27672 46900 27678 46912
rect 28537 46903 28595 46909
rect 28537 46900 28549 46903
rect 27672 46872 28549 46900
rect 27672 46860 27678 46872
rect 28537 46869 28549 46872
rect 28583 46869 28595 46903
rect 28718 46900 28724 46912
rect 28679 46872 28724 46900
rect 28537 46863 28595 46869
rect 28718 46860 28724 46872
rect 28776 46860 28782 46912
rect 28902 46860 28908 46912
rect 28960 46900 28966 46912
rect 32306 46900 32312 46912
rect 28960 46872 32312 46900
rect 28960 46860 28966 46872
rect 32306 46860 32312 46872
rect 32364 46860 32370 46912
rect 33318 46900 33324 46912
rect 33279 46872 33324 46900
rect 33318 46860 33324 46872
rect 33376 46860 33382 46912
rect 33962 46900 33968 46912
rect 33923 46872 33968 46900
rect 33962 46860 33968 46872
rect 34020 46860 34026 46912
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 27706 46656 27712 46708
rect 27764 46696 27770 46708
rect 28718 46696 28724 46708
rect 27764 46668 28724 46696
rect 27764 46656 27770 46668
rect 28718 46656 28724 46668
rect 28776 46696 28782 46708
rect 30101 46699 30159 46705
rect 30101 46696 30113 46699
rect 28776 46668 30113 46696
rect 28776 46656 28782 46668
rect 30101 46665 30113 46668
rect 30147 46696 30159 46699
rect 33318 46696 33324 46708
rect 30147 46668 33324 46696
rect 30147 46665 30159 46668
rect 30101 46659 30159 46665
rect 33318 46656 33324 46668
rect 33376 46656 33382 46708
rect 24857 46631 24915 46637
rect 24857 46628 24869 46631
rect 23308 46600 24869 46628
rect 1857 46563 1915 46569
rect 1857 46529 1869 46563
rect 1903 46560 1915 46563
rect 2314 46560 2320 46572
rect 1903 46532 2320 46560
rect 1903 46529 1915 46532
rect 1857 46523 1915 46529
rect 2314 46520 2320 46532
rect 2372 46520 2378 46572
rect 21266 46560 21272 46572
rect 21227 46532 21272 46560
rect 21266 46520 21272 46532
rect 21324 46520 21330 46572
rect 21453 46563 21511 46569
rect 21453 46529 21465 46563
rect 21499 46560 21511 46563
rect 21542 46560 21548 46572
rect 21499 46532 21548 46560
rect 21499 46529 21511 46532
rect 21453 46523 21511 46529
rect 21542 46520 21548 46532
rect 21600 46520 21606 46572
rect 22281 46563 22339 46569
rect 22281 46529 22293 46563
rect 22327 46560 22339 46563
rect 22370 46560 22376 46572
rect 22327 46532 22376 46560
rect 22327 46529 22339 46532
rect 22281 46523 22339 46529
rect 22370 46520 22376 46532
rect 22428 46520 22434 46572
rect 23014 46560 23020 46572
rect 22480 46532 23020 46560
rect 22480 46433 22508 46532
rect 23014 46520 23020 46532
rect 23072 46560 23078 46572
rect 23308 46569 23336 46600
rect 24857 46597 24869 46600
rect 24903 46628 24915 46631
rect 25130 46628 25136 46640
rect 24903 46600 25136 46628
rect 24903 46597 24915 46600
rect 24857 46591 24915 46597
rect 25130 46588 25136 46600
rect 25188 46628 25194 46640
rect 26510 46628 26516 46640
rect 25188 46600 26516 46628
rect 25188 46588 25194 46600
rect 23293 46563 23351 46569
rect 23293 46560 23305 46563
rect 23072 46532 23305 46560
rect 23072 46520 23078 46532
rect 23293 46529 23305 46532
rect 23339 46529 23351 46563
rect 24670 46560 24676 46572
rect 23293 46523 23351 46529
rect 24228 46532 24676 46560
rect 22465 46427 22523 46433
rect 22465 46393 22477 46427
rect 22511 46393 22523 46427
rect 24026 46424 24032 46436
rect 23939 46396 24032 46424
rect 22465 46387 22523 46393
rect 24026 46384 24032 46396
rect 24084 46424 24090 46436
rect 24228 46424 24256 46532
rect 24670 46520 24676 46532
rect 24728 46560 24734 46572
rect 25041 46563 25099 46569
rect 25041 46560 25053 46563
rect 24728 46532 25053 46560
rect 24728 46520 24734 46532
rect 25041 46529 25053 46532
rect 25087 46529 25099 46563
rect 25222 46560 25228 46572
rect 25183 46532 25228 46560
rect 25041 46523 25099 46529
rect 25222 46520 25228 46532
rect 25280 46520 25286 46572
rect 26050 46520 26056 46572
rect 26108 46560 26114 46572
rect 26344 46569 26372 46600
rect 26510 46588 26516 46600
rect 26568 46628 26574 46640
rect 27890 46628 27896 46640
rect 26568 46600 27896 46628
rect 26568 46588 26574 46600
rect 27890 46588 27896 46600
rect 27948 46628 27954 46640
rect 30650 46628 30656 46640
rect 27948 46600 28304 46628
rect 27948 46588 27954 46600
rect 26145 46563 26203 46569
rect 26145 46560 26157 46563
rect 26108 46532 26157 46560
rect 26108 46520 26114 46532
rect 26145 46529 26157 46532
rect 26191 46529 26203 46563
rect 26145 46523 26203 46529
rect 26329 46563 26387 46569
rect 26329 46529 26341 46563
rect 26375 46529 26387 46563
rect 26329 46523 26387 46529
rect 26605 46563 26663 46569
rect 26605 46529 26617 46563
rect 26651 46560 26663 46563
rect 26694 46560 26700 46572
rect 26651 46532 26700 46560
rect 26651 46529 26663 46532
rect 26605 46523 26663 46529
rect 26694 46520 26700 46532
rect 26752 46560 26758 46572
rect 27706 46560 27712 46572
rect 26752 46532 27712 46560
rect 26752 46520 26758 46532
rect 27706 46520 27712 46532
rect 27764 46520 27770 46572
rect 28077 46563 28135 46569
rect 28077 46529 28089 46563
rect 28123 46529 28135 46563
rect 28276 46558 28304 46600
rect 29012 46600 30656 46628
rect 28445 46563 28503 46569
rect 28445 46560 28457 46563
rect 28368 46558 28457 46560
rect 28276 46532 28457 46558
rect 28276 46530 28396 46532
rect 28077 46523 28135 46529
rect 28445 46529 28457 46532
rect 28491 46560 28503 46563
rect 28534 46560 28540 46572
rect 28491 46532 28540 46560
rect 28491 46529 28503 46532
rect 28445 46523 28503 46529
rect 24302 46452 24308 46504
rect 24360 46492 24366 46504
rect 24762 46492 24768 46504
rect 24360 46464 24768 46492
rect 24360 46452 24366 46464
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 28092 46492 28120 46523
rect 28534 46520 28540 46532
rect 28592 46520 28598 46572
rect 29012 46492 29040 46600
rect 30650 46588 30656 46600
rect 30708 46588 30714 46640
rect 32306 46588 32312 46640
rect 32364 46628 32370 46640
rect 33134 46628 33140 46640
rect 32364 46600 33140 46628
rect 32364 46588 32370 46600
rect 33134 46588 33140 46600
rect 33192 46628 33198 46640
rect 33505 46631 33563 46637
rect 33505 46628 33517 46631
rect 33192 46600 33517 46628
rect 33192 46588 33198 46600
rect 33505 46597 33517 46600
rect 33551 46597 33563 46631
rect 33505 46591 33563 46597
rect 29178 46520 29184 46572
rect 29236 46560 29242 46572
rect 29730 46560 29736 46572
rect 29236 46532 29736 46560
rect 29236 46520 29242 46532
rect 29730 46520 29736 46532
rect 29788 46560 29794 46572
rect 29917 46563 29975 46569
rect 29917 46560 29929 46563
rect 29788 46532 29929 46560
rect 29788 46520 29794 46532
rect 29917 46529 29929 46532
rect 29963 46529 29975 46563
rect 29917 46523 29975 46529
rect 30193 46563 30251 46569
rect 30193 46529 30205 46563
rect 30239 46529 30251 46563
rect 30193 46523 30251 46529
rect 31113 46563 31171 46569
rect 31113 46529 31125 46563
rect 31159 46560 31171 46563
rect 31294 46560 31300 46572
rect 31159 46532 31300 46560
rect 31159 46529 31171 46532
rect 31113 46523 31171 46529
rect 28092 46464 29040 46492
rect 30208 46492 30236 46523
rect 31294 46520 31300 46532
rect 31352 46560 31358 46572
rect 32401 46563 32459 46569
rect 31352 46532 32260 46560
rect 31352 46520 31358 46532
rect 32232 46492 32260 46532
rect 32401 46529 32413 46563
rect 32447 46529 32459 46563
rect 32401 46523 32459 46529
rect 32306 46492 32312 46504
rect 30208 46464 31754 46492
rect 32232 46464 32312 46492
rect 25130 46424 25136 46436
rect 24084 46396 24256 46424
rect 25091 46396 25136 46424
rect 24084 46384 24090 46396
rect 25130 46384 25136 46396
rect 25188 46384 25194 46436
rect 26421 46427 26479 46433
rect 25240 46396 26280 46424
rect 1670 46356 1676 46368
rect 1631 46328 1676 46356
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 2314 46356 2320 46368
rect 2275 46328 2320 46356
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 20806 46316 20812 46368
rect 20864 46356 20870 46368
rect 21453 46359 21511 46365
rect 21453 46356 21465 46359
rect 20864 46328 21465 46356
rect 20864 46316 20870 46328
rect 21453 46325 21465 46328
rect 21499 46325 21511 46359
rect 21453 46319 21511 46325
rect 22094 46316 22100 46368
rect 22152 46356 22158 46368
rect 23109 46359 23167 46365
rect 23109 46356 23121 46359
rect 22152 46328 23121 46356
rect 22152 46316 22158 46328
rect 23109 46325 23121 46328
rect 23155 46356 23167 46359
rect 23658 46356 23664 46368
rect 23155 46328 23664 46356
rect 23155 46325 23167 46328
rect 23109 46319 23167 46325
rect 23658 46316 23664 46328
rect 23716 46316 23722 46368
rect 23842 46356 23848 46368
rect 23803 46328 23848 46356
rect 23842 46316 23848 46328
rect 23900 46316 23906 46368
rect 24762 46316 24768 46368
rect 24820 46356 24826 46368
rect 25240 46356 25268 46396
rect 25866 46356 25872 46368
rect 24820 46328 25268 46356
rect 25827 46328 25872 46356
rect 24820 46316 24826 46328
rect 25866 46316 25872 46328
rect 25924 46316 25930 46368
rect 26252 46365 26280 46396
rect 26421 46393 26433 46427
rect 26467 46424 26479 46427
rect 26786 46424 26792 46436
rect 26467 46396 26792 46424
rect 26467 46393 26479 46396
rect 26421 46387 26479 46393
rect 26786 46384 26792 46396
rect 26844 46384 26850 46436
rect 28092 46424 28120 46464
rect 27080 46396 28120 46424
rect 26237 46359 26295 46365
rect 26237 46325 26249 46359
rect 26283 46356 26295 46359
rect 27080 46356 27108 46396
rect 28258 46384 28264 46436
rect 28316 46424 28322 46436
rect 28902 46424 28908 46436
rect 28316 46396 28908 46424
rect 28316 46384 28322 46396
rect 28902 46384 28908 46396
rect 28960 46424 28966 46436
rect 30208 46424 30236 46464
rect 28960 46396 30236 46424
rect 28960 46384 28966 46396
rect 30282 46384 30288 46436
rect 30340 46424 30346 46436
rect 31573 46427 31631 46433
rect 31573 46424 31585 46427
rect 30340 46396 31585 46424
rect 30340 46384 30346 46396
rect 31573 46393 31585 46396
rect 31619 46393 31631 46427
rect 31726 46424 31754 46464
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32416 46492 32444 46523
rect 32490 46520 32496 46572
rect 32548 46560 32554 46572
rect 33229 46563 33287 46569
rect 33229 46560 33241 46563
rect 32548 46532 33241 46560
rect 32548 46520 32554 46532
rect 33229 46529 33241 46532
rect 33275 46529 33287 46563
rect 33229 46523 33287 46529
rect 32582 46492 32588 46504
rect 32416 46464 32588 46492
rect 32582 46452 32588 46464
rect 32640 46452 32646 46504
rect 31726 46396 32720 46424
rect 31573 46387 31631 46393
rect 26283 46328 27108 46356
rect 26283 46325 26295 46328
rect 26237 46319 26295 46325
rect 27430 46316 27436 46368
rect 27488 46356 27494 46368
rect 27525 46359 27583 46365
rect 27525 46356 27537 46359
rect 27488 46328 27537 46356
rect 27488 46316 27494 46328
rect 27525 46325 27537 46328
rect 27571 46325 27583 46359
rect 28442 46356 28448 46368
rect 28403 46328 28448 46356
rect 27525 46319 27583 46325
rect 28442 46316 28448 46328
rect 28500 46316 28506 46368
rect 28534 46316 28540 46368
rect 28592 46356 28598 46368
rect 28629 46359 28687 46365
rect 28629 46356 28641 46359
rect 28592 46328 28641 46356
rect 28592 46316 28598 46328
rect 28629 46325 28641 46328
rect 28675 46325 28687 46359
rect 29270 46356 29276 46368
rect 29231 46328 29276 46356
rect 28629 46319 28687 46325
rect 29270 46316 29276 46328
rect 29328 46316 29334 46368
rect 29730 46356 29736 46368
rect 29691 46328 29736 46356
rect 29730 46316 29736 46328
rect 29788 46316 29794 46368
rect 30650 46316 30656 46368
rect 30708 46356 30714 46368
rect 30929 46359 30987 46365
rect 30929 46356 30941 46359
rect 30708 46328 30941 46356
rect 30708 46316 30714 46328
rect 30929 46325 30941 46328
rect 30975 46325 30987 46359
rect 31588 46356 31616 46387
rect 31846 46356 31852 46368
rect 31588 46328 31852 46356
rect 30929 46319 30987 46325
rect 31846 46316 31852 46328
rect 31904 46316 31910 46368
rect 32692 46365 32720 46396
rect 32677 46359 32735 46365
rect 32677 46325 32689 46359
rect 32723 46356 32735 46359
rect 33778 46356 33784 46368
rect 32723 46328 33784 46356
rect 32723 46325 32735 46328
rect 32677 46319 32735 46325
rect 33778 46316 33784 46328
rect 33836 46316 33842 46368
rect 34146 46356 34152 46368
rect 34107 46328 34152 46356
rect 34146 46316 34152 46328
rect 34204 46316 34210 46368
rect 34698 46356 34704 46368
rect 34659 46328 34704 46356
rect 34698 46316 34704 46328
rect 34756 46316 34762 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 29270 46112 29276 46164
rect 29328 46152 29334 46164
rect 31202 46152 31208 46164
rect 29328 46124 31208 46152
rect 29328 46112 29334 46124
rect 31202 46112 31208 46124
rect 31260 46112 31266 46164
rect 22370 46044 22376 46096
rect 22428 46084 22434 46096
rect 27338 46084 27344 46096
rect 22428 46056 27344 46084
rect 22428 46044 22434 46056
rect 27338 46044 27344 46056
rect 27396 46044 27402 46096
rect 27982 46044 27988 46096
rect 28040 46084 28046 46096
rect 30742 46084 30748 46096
rect 28040 46056 28856 46084
rect 30703 46056 30748 46084
rect 28040 46044 28046 46056
rect 24026 46016 24032 46028
rect 23768 45988 24032 46016
rect 22554 45948 22560 45960
rect 22515 45920 22560 45948
rect 22554 45908 22560 45920
rect 22612 45908 22618 45960
rect 22833 45951 22891 45957
rect 22833 45917 22845 45951
rect 22879 45948 22891 45951
rect 23198 45948 23204 45960
rect 22879 45920 23204 45948
rect 22879 45917 22891 45920
rect 22833 45911 22891 45917
rect 23198 45908 23204 45920
rect 23256 45908 23262 45960
rect 23768 45957 23796 45988
rect 24026 45976 24032 45988
rect 24084 45976 24090 46028
rect 24578 45976 24584 46028
rect 24636 46016 24642 46028
rect 25869 46019 25927 46025
rect 25869 46016 25881 46019
rect 24636 45988 25881 46016
rect 24636 45976 24642 45988
rect 25869 45985 25881 45988
rect 25915 46016 25927 46019
rect 27430 46016 27436 46028
rect 25915 45988 27436 46016
rect 25915 45985 25927 45988
rect 25869 45979 25927 45985
rect 27430 45976 27436 45988
rect 27488 45976 27494 46028
rect 27798 46016 27804 46028
rect 27646 45988 27804 46016
rect 23753 45951 23811 45957
rect 23753 45917 23765 45951
rect 23799 45917 23811 45951
rect 23753 45911 23811 45917
rect 23937 45951 23995 45957
rect 23937 45917 23949 45951
rect 23983 45948 23995 45951
rect 24302 45948 24308 45960
rect 23983 45920 24308 45948
rect 23983 45917 23995 45920
rect 23937 45911 23995 45917
rect 24302 45908 24308 45920
rect 24360 45908 24366 45960
rect 24765 45951 24823 45957
rect 24765 45917 24777 45951
rect 24811 45917 24823 45951
rect 24946 45948 24952 45960
rect 24907 45920 24952 45948
rect 24765 45911 24823 45917
rect 21545 45883 21603 45889
rect 21545 45880 21557 45883
rect 20456 45852 21557 45880
rect 20456 45824 20484 45852
rect 21545 45849 21557 45852
rect 21591 45849 21603 45883
rect 21545 45843 21603 45849
rect 21913 45883 21971 45889
rect 21913 45849 21925 45883
rect 21959 45880 21971 45883
rect 22278 45880 22284 45892
rect 21959 45852 22284 45880
rect 21959 45849 21971 45852
rect 21913 45843 21971 45849
rect 22278 45840 22284 45852
rect 22336 45840 22342 45892
rect 23566 45840 23572 45892
rect 23624 45880 23630 45892
rect 24581 45883 24639 45889
rect 24581 45880 24593 45883
rect 23624 45852 24593 45880
rect 23624 45840 23630 45852
rect 24581 45849 24593 45852
rect 24627 45849 24639 45883
rect 24780 45880 24808 45911
rect 24946 45908 24952 45920
rect 25004 45908 25010 45960
rect 25041 45951 25099 45957
rect 25041 45917 25053 45951
rect 25087 45948 25099 45951
rect 26142 45948 26148 45960
rect 25087 45920 26148 45948
rect 25087 45917 25099 45920
rect 25041 45911 25099 45917
rect 26142 45908 26148 45920
rect 26200 45908 26206 45960
rect 26513 45951 26571 45957
rect 26513 45917 26525 45951
rect 26559 45948 26571 45951
rect 26694 45948 26700 45960
rect 26559 45920 26700 45948
rect 26559 45917 26571 45920
rect 26513 45911 26571 45917
rect 26694 45908 26700 45920
rect 26752 45908 26758 45960
rect 26970 45948 26976 45960
rect 26931 45920 26976 45948
rect 26970 45908 26976 45920
rect 27028 45948 27034 45960
rect 27646 45957 27674 45988
rect 27798 45976 27804 45988
rect 27856 46016 27862 46028
rect 28258 46016 28264 46028
rect 27856 45988 28264 46016
rect 27856 45976 27862 45988
rect 28258 45976 28264 45988
rect 28316 45976 28322 46028
rect 28828 46025 28856 46056
rect 30742 46044 30748 46056
rect 30800 46044 30806 46096
rect 28813 46019 28871 46025
rect 28813 45985 28825 46019
rect 28859 46016 28871 46019
rect 28859 45988 30604 46016
rect 28859 45985 28871 45988
rect 28813 45979 28871 45985
rect 27617 45951 27675 45957
rect 27028 45920 27568 45948
rect 27028 45908 27034 45920
rect 26602 45880 26608 45892
rect 24780 45852 26608 45880
rect 24581 45843 24639 45849
rect 26602 45840 26608 45852
rect 26660 45880 26666 45892
rect 27433 45883 27491 45889
rect 27433 45880 27445 45883
rect 26660 45852 27445 45880
rect 26660 45840 26666 45852
rect 27433 45849 27445 45852
rect 27479 45849 27491 45883
rect 27540 45880 27568 45920
rect 27617 45917 27629 45951
rect 27663 45917 27675 45951
rect 27617 45911 27675 45917
rect 27706 45908 27712 45960
rect 27764 45948 27770 45960
rect 27890 45948 27896 45960
rect 27764 45920 27809 45948
rect 27851 45920 27896 45948
rect 27764 45908 27770 45920
rect 27890 45908 27896 45920
rect 27948 45908 27954 45960
rect 27985 45951 28043 45957
rect 27985 45917 27997 45951
rect 28031 45917 28043 45951
rect 27985 45911 28043 45917
rect 28000 45880 28028 45911
rect 28902 45908 28908 45960
rect 28960 45948 28966 45960
rect 28997 45951 29055 45957
rect 28997 45948 29009 45951
rect 28960 45920 29009 45948
rect 28960 45908 28966 45920
rect 28997 45917 29009 45920
rect 29043 45917 29055 45951
rect 28997 45911 29055 45917
rect 29730 45908 29736 45960
rect 29788 45948 29794 45960
rect 29917 45951 29975 45957
rect 29917 45948 29929 45951
rect 29788 45920 29929 45948
rect 29788 45908 29794 45920
rect 29917 45917 29929 45920
rect 29963 45917 29975 45951
rect 29917 45911 29975 45917
rect 30193 45951 30251 45957
rect 30193 45917 30205 45951
rect 30239 45948 30251 45951
rect 30282 45948 30288 45960
rect 30239 45920 30288 45948
rect 30239 45917 30251 45920
rect 30193 45911 30251 45917
rect 29178 45880 29184 45892
rect 27540 45852 28028 45880
rect 29091 45852 29184 45880
rect 27433 45843 27491 45849
rect 29178 45840 29184 45852
rect 29236 45840 29242 45892
rect 29362 45840 29368 45892
rect 29420 45880 29426 45892
rect 30208 45880 30236 45911
rect 30282 45908 30288 45920
rect 30340 45908 30346 45960
rect 30576 45957 30604 45988
rect 30650 45976 30656 46028
rect 30708 46016 30714 46028
rect 31846 46016 31852 46028
rect 30708 45988 30753 46016
rect 31807 45988 31852 46016
rect 30708 45976 30714 45988
rect 31846 45976 31852 45988
rect 31904 45976 31910 46028
rect 33318 45976 33324 46028
rect 33376 46016 33382 46028
rect 33376 45988 33916 46016
rect 33376 45976 33382 45988
rect 30561 45951 30619 45957
rect 30561 45917 30573 45951
rect 30607 45917 30619 45951
rect 30561 45911 30619 45917
rect 32125 45951 32183 45957
rect 32125 45917 32137 45951
rect 32171 45948 32183 45951
rect 32490 45948 32496 45960
rect 32171 45920 32496 45948
rect 32171 45917 32183 45920
rect 32125 45911 32183 45917
rect 32490 45908 32496 45920
rect 32548 45908 32554 45960
rect 32585 45951 32643 45957
rect 32585 45917 32597 45951
rect 32631 45917 32643 45951
rect 32585 45911 32643 45917
rect 32953 45951 33011 45957
rect 32953 45917 32965 45951
rect 32999 45948 33011 45951
rect 33594 45948 33600 45960
rect 32999 45920 33600 45948
rect 32999 45917 33011 45920
rect 32953 45911 33011 45917
rect 29420 45852 30236 45880
rect 32600 45880 32628 45911
rect 33594 45908 33600 45920
rect 33652 45908 33658 45960
rect 33689 45951 33747 45957
rect 33689 45917 33701 45951
rect 33735 45948 33747 45951
rect 33778 45948 33784 45960
rect 33735 45920 33784 45948
rect 33735 45917 33747 45920
rect 33689 45911 33747 45917
rect 33704 45880 33732 45911
rect 33778 45908 33784 45920
rect 33836 45908 33842 45960
rect 33888 45957 33916 45988
rect 33873 45951 33931 45957
rect 33873 45917 33885 45951
rect 33919 45917 33931 45951
rect 58069 45951 58127 45957
rect 58069 45948 58081 45951
rect 33873 45911 33931 45917
rect 57532 45920 58081 45948
rect 32600 45852 33732 45880
rect 29420 45840 29426 45852
rect 1854 45772 1860 45824
rect 1912 45812 1918 45824
rect 20438 45812 20444 45824
rect 1912 45784 20444 45812
rect 1912 45772 1918 45784
rect 20438 45772 20444 45784
rect 20496 45772 20502 45824
rect 20993 45815 21051 45821
rect 20993 45781 21005 45815
rect 21039 45812 21051 45815
rect 21082 45812 21088 45824
rect 21039 45784 21088 45812
rect 21039 45781 21051 45784
rect 20993 45775 21051 45781
rect 21082 45772 21088 45784
rect 21140 45772 21146 45824
rect 22370 45812 22376 45824
rect 22331 45784 22376 45812
rect 22370 45772 22376 45784
rect 22428 45772 22434 45824
rect 22738 45812 22744 45824
rect 22699 45784 22744 45812
rect 22738 45772 22744 45784
rect 22796 45772 22802 45824
rect 23474 45772 23480 45824
rect 23532 45812 23538 45824
rect 23845 45815 23903 45821
rect 23845 45812 23857 45815
rect 23532 45784 23857 45812
rect 23532 45772 23538 45784
rect 23845 45781 23857 45784
rect 23891 45781 23903 45815
rect 23845 45775 23903 45781
rect 24026 45772 24032 45824
rect 24084 45812 24090 45824
rect 26513 45815 26571 45821
rect 26513 45812 26525 45815
rect 24084 45784 26525 45812
rect 24084 45772 24090 45784
rect 26513 45781 26525 45784
rect 26559 45781 26571 45815
rect 26513 45775 26571 45781
rect 27338 45772 27344 45824
rect 27396 45812 27402 45824
rect 29196 45812 29224 45840
rect 31294 45812 31300 45824
rect 27396 45784 31300 45812
rect 27396 45772 27402 45784
rect 31294 45772 31300 45784
rect 31352 45772 31358 45824
rect 33870 45812 33876 45824
rect 33831 45784 33876 45812
rect 33870 45772 33876 45784
rect 33928 45772 33934 45824
rect 33962 45772 33968 45824
rect 34020 45812 34026 45824
rect 34698 45812 34704 45824
rect 34020 45784 34704 45812
rect 34020 45772 34026 45784
rect 34698 45772 34704 45784
rect 34756 45812 34762 45824
rect 34885 45815 34943 45821
rect 34885 45812 34897 45815
rect 34756 45784 34897 45812
rect 34756 45772 34762 45784
rect 34885 45781 34897 45784
rect 34931 45781 34943 45815
rect 34885 45775 34943 45781
rect 57330 45772 57336 45824
rect 57388 45812 57394 45824
rect 57532 45821 57560 45920
rect 58069 45917 58081 45920
rect 58115 45917 58127 45951
rect 58069 45911 58127 45917
rect 57517 45815 57575 45821
rect 57517 45812 57529 45815
rect 57388 45784 57529 45812
rect 57388 45772 57394 45784
rect 57517 45781 57529 45784
rect 57563 45781 57575 45815
rect 58250 45812 58256 45824
rect 58211 45784 58256 45812
rect 57517 45775 57575 45781
rect 58250 45772 58256 45784
rect 58308 45772 58314 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 22281 45611 22339 45617
rect 22281 45577 22293 45611
rect 22327 45608 22339 45611
rect 22370 45608 22376 45620
rect 22327 45580 22376 45608
rect 22327 45577 22339 45580
rect 22281 45571 22339 45577
rect 22370 45568 22376 45580
rect 22428 45568 22434 45620
rect 22554 45568 22560 45620
rect 22612 45608 22618 45620
rect 25130 45608 25136 45620
rect 22612 45580 25136 45608
rect 22612 45568 22618 45580
rect 25130 45568 25136 45580
rect 25188 45568 25194 45620
rect 30926 45608 30932 45620
rect 27264 45580 29868 45608
rect 30887 45580 30932 45608
rect 27264 45552 27292 45580
rect 21450 45540 21456 45552
rect 21008 45512 21456 45540
rect 20714 45432 20720 45484
rect 20772 45472 20778 45484
rect 20809 45475 20867 45481
rect 20809 45472 20821 45475
rect 20772 45444 20821 45472
rect 20772 45432 20778 45444
rect 20809 45441 20821 45444
rect 20855 45472 20867 45475
rect 20898 45472 20904 45484
rect 20855 45444 20904 45472
rect 20855 45441 20867 45444
rect 20809 45435 20867 45441
rect 20898 45432 20904 45444
rect 20956 45432 20962 45484
rect 21008 45481 21036 45512
rect 21450 45500 21456 45512
rect 21508 45500 21514 45552
rect 24854 45500 24860 45552
rect 24912 45540 24918 45552
rect 25685 45543 25743 45549
rect 25685 45540 25697 45543
rect 24912 45512 25697 45540
rect 24912 45500 24918 45512
rect 25685 45509 25697 45512
rect 25731 45509 25743 45543
rect 27246 45540 27252 45552
rect 27207 45512 27252 45540
rect 25685 45503 25743 45509
rect 27246 45500 27252 45512
rect 27304 45500 27310 45552
rect 29086 45540 29092 45552
rect 28552 45512 29092 45540
rect 20993 45475 21051 45481
rect 20993 45441 21005 45475
rect 21039 45441 21051 45475
rect 20993 45435 21051 45441
rect 21269 45475 21327 45481
rect 21269 45441 21281 45475
rect 21315 45472 21327 45475
rect 21358 45472 21364 45484
rect 21315 45444 21364 45472
rect 21315 45441 21327 45444
rect 21269 45435 21327 45441
rect 21358 45432 21364 45444
rect 21416 45432 21422 45484
rect 22186 45472 22192 45484
rect 22147 45444 22192 45472
rect 22186 45432 22192 45444
rect 22244 45432 22250 45484
rect 22370 45432 22376 45484
rect 22428 45472 22434 45484
rect 22465 45475 22523 45481
rect 22465 45472 22477 45475
rect 22428 45444 22477 45472
rect 22428 45432 22434 45444
rect 22465 45441 22477 45444
rect 22511 45441 22523 45475
rect 23290 45472 23296 45484
rect 23251 45444 23296 45472
rect 22465 45435 22523 45441
rect 23290 45432 23296 45444
rect 23348 45432 23354 45484
rect 24581 45475 24639 45481
rect 24581 45472 24593 45475
rect 23492 45444 24593 45472
rect 23492 45416 23520 45444
rect 24581 45441 24593 45444
rect 24627 45441 24639 45475
rect 25041 45475 25099 45481
rect 25041 45472 25053 45475
rect 24581 45435 24639 45441
rect 24688 45444 25053 45472
rect 21082 45404 21088 45416
rect 20995 45376 21088 45404
rect 21082 45364 21088 45376
rect 21140 45364 21146 45416
rect 21177 45407 21235 45413
rect 21177 45373 21189 45407
rect 21223 45404 21235 45407
rect 23474 45404 23480 45416
rect 21223 45376 23480 45404
rect 21223 45373 21235 45376
rect 21177 45367 21235 45373
rect 23474 45364 23480 45376
rect 23532 45364 23538 45416
rect 23569 45407 23627 45413
rect 23569 45373 23581 45407
rect 23615 45404 23627 45407
rect 24302 45404 24308 45416
rect 23615 45376 24308 45404
rect 23615 45373 23627 45376
rect 23569 45367 23627 45373
rect 24302 45364 24308 45376
rect 24360 45364 24366 45416
rect 24688 45404 24716 45444
rect 25041 45441 25053 45444
rect 25087 45441 25099 45475
rect 25498 45472 25504 45484
rect 25411 45444 25504 45472
rect 25041 45435 25099 45441
rect 25498 45432 25504 45444
rect 25556 45432 25562 45484
rect 25777 45475 25835 45481
rect 25777 45441 25789 45475
rect 25823 45472 25835 45475
rect 26142 45472 26148 45484
rect 25823 45444 26148 45472
rect 25823 45441 25835 45444
rect 25777 45435 25835 45441
rect 26142 45432 26148 45444
rect 26200 45432 26206 45484
rect 26418 45472 26424 45484
rect 26379 45444 26424 45472
rect 26418 45432 26424 45444
rect 26476 45432 26482 45484
rect 26602 45472 26608 45484
rect 26563 45444 26608 45472
rect 26602 45432 26608 45444
rect 26660 45432 26666 45484
rect 28552 45481 28580 45512
rect 29086 45500 29092 45512
rect 29144 45540 29150 45552
rect 29730 45540 29736 45552
rect 29144 45512 29736 45540
rect 29144 45500 29150 45512
rect 29730 45500 29736 45512
rect 29788 45500 29794 45552
rect 28537 45475 28595 45481
rect 28537 45441 28549 45475
rect 28583 45441 28595 45475
rect 28537 45435 28595 45441
rect 28813 45475 28871 45481
rect 28813 45441 28825 45475
rect 28859 45441 28871 45475
rect 28813 45435 28871 45441
rect 24504 45376 24716 45404
rect 24765 45407 24823 45413
rect 21100 45336 21128 45364
rect 24504 45336 24532 45376
rect 24765 45373 24777 45407
rect 24811 45373 24823 45407
rect 24765 45367 24823 45373
rect 24857 45407 24915 45413
rect 24857 45373 24869 45407
rect 24903 45404 24915 45407
rect 24946 45404 24952 45416
rect 24903 45376 24952 45404
rect 24903 45373 24915 45376
rect 24857 45367 24915 45373
rect 24670 45336 24676 45348
rect 21100 45308 23244 45336
rect 23216 45280 23244 45308
rect 23492 45308 24532 45336
rect 24631 45308 24676 45336
rect 21174 45228 21180 45280
rect 21232 45268 21238 45280
rect 21453 45271 21511 45277
rect 21453 45268 21465 45271
rect 21232 45240 21465 45268
rect 21232 45228 21238 45240
rect 21453 45237 21465 45240
rect 21499 45237 21511 45271
rect 22646 45268 22652 45280
rect 22607 45240 22652 45268
rect 21453 45231 21511 45237
rect 22646 45228 22652 45240
rect 22704 45228 22710 45280
rect 23106 45268 23112 45280
rect 23067 45240 23112 45268
rect 23106 45228 23112 45240
rect 23164 45228 23170 45280
rect 23198 45228 23204 45280
rect 23256 45268 23262 45280
rect 23492 45277 23520 45308
rect 24670 45296 24676 45308
rect 24728 45296 24734 45348
rect 24780 45336 24808 45367
rect 24946 45364 24952 45376
rect 25004 45404 25010 45416
rect 25516 45404 25544 45432
rect 25004 45376 25452 45404
rect 25516 45376 25820 45404
rect 25004 45364 25010 45376
rect 25222 45336 25228 45348
rect 24780 45308 25228 45336
rect 25222 45296 25228 45308
rect 25280 45296 25286 45348
rect 25424 45336 25452 45376
rect 25682 45336 25688 45348
rect 25424 45308 25688 45336
rect 25682 45296 25688 45308
rect 25740 45296 25746 45348
rect 25792 45336 25820 45376
rect 27430 45364 27436 45416
rect 27488 45404 27494 45416
rect 28828 45404 28856 45435
rect 28902 45432 28908 45484
rect 28960 45472 28966 45484
rect 28997 45475 29055 45481
rect 28997 45472 29009 45475
rect 28960 45444 29009 45472
rect 28960 45432 28966 45444
rect 28997 45441 29009 45444
rect 29043 45441 29055 45475
rect 29840 45472 29868 45580
rect 30926 45568 30932 45580
rect 30984 45568 30990 45620
rect 31018 45568 31024 45620
rect 31076 45608 31082 45620
rect 31076 45580 31121 45608
rect 31076 45568 31082 45580
rect 31202 45568 31208 45620
rect 31260 45608 31266 45620
rect 33410 45608 33416 45620
rect 31260 45580 33416 45608
rect 31260 45568 31266 45580
rect 33410 45568 33416 45580
rect 33468 45568 33474 45620
rect 34520 45552 34572 45558
rect 30208 45512 33640 45540
rect 30208 45481 30236 45512
rect 33612 45484 33640 45512
rect 34520 45494 34572 45500
rect 30193 45475 30251 45481
rect 30193 45472 30205 45475
rect 29840 45444 30205 45472
rect 28997 45435 29055 45441
rect 30193 45441 30205 45444
rect 30239 45441 30251 45475
rect 30193 45435 30251 45441
rect 30650 45432 30656 45484
rect 30708 45472 30714 45484
rect 30837 45475 30895 45481
rect 30837 45472 30849 45475
rect 30708 45444 30849 45472
rect 30708 45432 30714 45444
rect 30837 45441 30849 45444
rect 30883 45441 30895 45475
rect 30837 45435 30895 45441
rect 31018 45432 31024 45484
rect 31076 45472 31082 45484
rect 31205 45475 31263 45481
rect 31205 45472 31217 45475
rect 31076 45444 31217 45472
rect 31076 45432 31082 45444
rect 31205 45441 31217 45444
rect 31251 45441 31263 45475
rect 31205 45435 31263 45441
rect 31294 45432 31300 45484
rect 31352 45472 31358 45484
rect 32586 45475 32644 45481
rect 32586 45472 32598 45475
rect 31352 45444 32598 45472
rect 31352 45432 31358 45444
rect 32586 45441 32598 45444
rect 32632 45441 32644 45475
rect 32586 45435 32644 45441
rect 32953 45475 33011 45481
rect 32953 45441 32965 45475
rect 32999 45472 33011 45475
rect 33318 45472 33324 45484
rect 32999 45444 33324 45472
rect 32999 45441 33011 45444
rect 32953 45435 33011 45441
rect 33318 45432 33324 45444
rect 33376 45432 33382 45484
rect 33594 45472 33600 45484
rect 33555 45444 33600 45472
rect 33594 45432 33600 45444
rect 33652 45432 33658 45484
rect 33962 45472 33968 45484
rect 33796 45444 33968 45472
rect 33045 45407 33103 45413
rect 33045 45404 33057 45407
rect 27488 45376 31340 45404
rect 27488 45364 27494 45376
rect 26878 45336 26884 45348
rect 25792 45308 26884 45336
rect 26878 45296 26884 45308
rect 26936 45296 26942 45348
rect 27617 45339 27675 45345
rect 27617 45305 27629 45339
rect 27663 45336 27675 45339
rect 27798 45336 27804 45348
rect 27663 45308 27804 45336
rect 27663 45305 27675 45308
rect 27617 45299 27675 45305
rect 27798 45296 27804 45308
rect 27856 45336 27862 45348
rect 28074 45336 28080 45348
rect 27856 45308 28080 45336
rect 27856 45296 27862 45308
rect 28074 45296 28080 45308
rect 28132 45296 28138 45348
rect 30653 45339 30711 45345
rect 30653 45305 30665 45339
rect 30699 45336 30711 45339
rect 30834 45336 30840 45348
rect 30699 45308 30840 45336
rect 30699 45305 30711 45308
rect 30653 45299 30711 45305
rect 30834 45296 30840 45308
rect 30892 45296 30898 45348
rect 31312 45280 31340 45376
rect 32600 45376 33057 45404
rect 32600 45348 32628 45376
rect 33045 45373 33057 45376
rect 33091 45404 33103 45407
rect 33796 45404 33824 45444
rect 33962 45432 33968 45444
rect 34020 45432 34026 45484
rect 34422 45472 34428 45484
rect 34383 45444 34428 45472
rect 34422 45432 34428 45444
rect 34480 45432 34486 45484
rect 33091 45376 33824 45404
rect 33091 45373 33103 45376
rect 33045 45367 33103 45373
rect 32306 45296 32312 45348
rect 32364 45336 32370 45348
rect 32401 45339 32459 45345
rect 32401 45336 32413 45339
rect 32364 45308 32413 45336
rect 32364 45296 32370 45308
rect 32401 45305 32413 45308
rect 32447 45305 32459 45339
rect 32401 45299 32459 45305
rect 32582 45296 32588 45348
rect 32640 45296 32646 45348
rect 23477 45271 23535 45277
rect 23477 45268 23489 45271
rect 23256 45240 23489 45268
rect 23256 45228 23262 45240
rect 23477 45237 23489 45240
rect 23523 45237 23535 45271
rect 24394 45268 24400 45280
rect 24355 45240 24400 45268
rect 23477 45231 23535 45237
rect 24394 45228 24400 45240
rect 24452 45228 24458 45280
rect 25774 45268 25780 45280
rect 25735 45240 25780 45268
rect 25774 45228 25780 45240
rect 25832 45228 25838 45280
rect 26510 45268 26516 45280
rect 26471 45240 26516 45268
rect 26510 45228 26516 45240
rect 26568 45228 26574 45280
rect 27522 45228 27528 45280
rect 27580 45268 27586 45280
rect 27709 45271 27767 45277
rect 27709 45268 27721 45271
rect 27580 45240 27721 45268
rect 27580 45228 27586 45240
rect 27709 45237 27721 45240
rect 27755 45237 27767 45271
rect 28350 45268 28356 45280
rect 28311 45240 28356 45268
rect 27709 45231 27767 45237
rect 28350 45228 28356 45240
rect 28408 45228 28414 45280
rect 29730 45268 29736 45280
rect 29691 45240 29736 45268
rect 29730 45228 29736 45240
rect 29788 45228 29794 45280
rect 30098 45268 30104 45280
rect 30059 45240 30104 45268
rect 30098 45228 30104 45240
rect 30156 45228 30162 45280
rect 31294 45228 31300 45280
rect 31352 45268 31358 45280
rect 31665 45271 31723 45277
rect 31665 45268 31677 45271
rect 31352 45240 31677 45268
rect 31352 45228 31358 45240
rect 31665 45237 31677 45240
rect 31711 45237 31723 45271
rect 31665 45231 31723 45237
rect 34422 45228 34428 45280
rect 34480 45268 34486 45280
rect 35894 45268 35900 45280
rect 34480 45240 35900 45268
rect 34480 45228 34486 45240
rect 35894 45228 35900 45240
rect 35952 45228 35958 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 21453 45067 21511 45073
rect 21453 45033 21465 45067
rect 21499 45033 21511 45067
rect 21453 45027 21511 45033
rect 20073 44931 20131 44937
rect 20073 44897 20085 44931
rect 20119 44928 20131 44931
rect 21082 44928 21088 44940
rect 20119 44900 21088 44928
rect 20119 44897 20131 44900
rect 20073 44891 20131 44897
rect 21082 44888 21088 44900
rect 21140 44888 21146 44940
rect 21468 44928 21496 45027
rect 22186 45024 22192 45076
rect 22244 45064 22250 45076
rect 23293 45067 23351 45073
rect 23293 45064 23305 45067
rect 22244 45036 23305 45064
rect 22244 45024 22250 45036
rect 23293 45033 23305 45036
rect 23339 45033 23351 45067
rect 23293 45027 23351 45033
rect 26878 45024 26884 45076
rect 26936 45064 26942 45076
rect 34146 45064 34152 45076
rect 26936 45036 29960 45064
rect 34107 45036 34152 45064
rect 26936 45024 26942 45036
rect 22370 44956 22376 45008
rect 22428 44996 22434 45008
rect 22428 44968 26004 44996
rect 22428 44956 22434 44968
rect 21468 44900 22140 44928
rect 20625 44863 20683 44869
rect 20625 44829 20637 44863
rect 20671 44860 20683 44863
rect 20990 44860 20996 44872
rect 20671 44832 20996 44860
rect 20671 44829 20683 44832
rect 20625 44823 20683 44829
rect 20990 44820 20996 44832
rect 21048 44820 21054 44872
rect 21361 44863 21419 44869
rect 21361 44829 21373 44863
rect 21407 44829 21419 44863
rect 21361 44823 21419 44829
rect 21376 44792 21404 44823
rect 21450 44820 21456 44872
rect 21508 44860 21514 44872
rect 22112 44860 22140 44900
rect 22186 44888 22192 44940
rect 22244 44928 22250 44940
rect 22244 44900 22784 44928
rect 22244 44888 22250 44900
rect 22462 44860 22468 44872
rect 21508 44832 21553 44860
rect 22112 44832 22468 44860
rect 21508 44820 21514 44832
rect 22462 44820 22468 44832
rect 22520 44820 22526 44872
rect 22756 44869 22784 44900
rect 23382 44888 23388 44940
rect 23440 44928 23446 44940
rect 23652 44931 23710 44937
rect 23652 44928 23664 44931
rect 23440 44900 23664 44928
rect 23440 44888 23446 44900
rect 23652 44897 23664 44900
rect 23698 44897 23710 44931
rect 23652 44891 23710 44897
rect 23753 44931 23811 44937
rect 23753 44897 23765 44931
rect 23799 44928 23811 44931
rect 24854 44928 24860 44940
rect 23799 44900 24860 44928
rect 23799 44897 23811 44900
rect 23753 44891 23811 44897
rect 22557 44863 22615 44869
rect 22557 44829 22569 44863
rect 22603 44860 22615 44863
rect 22741 44863 22799 44869
rect 22603 44832 22692 44860
rect 22603 44829 22615 44832
rect 22557 44823 22615 44829
rect 22002 44792 22008 44804
rect 21376 44764 22008 44792
rect 22002 44752 22008 44764
rect 22060 44792 22066 44804
rect 22094 44792 22100 44804
rect 22060 44764 22100 44792
rect 22060 44752 22066 44764
rect 22094 44752 22100 44764
rect 22152 44752 22158 44804
rect 19521 44727 19579 44733
rect 19521 44693 19533 44727
rect 19567 44724 19579 44727
rect 20530 44724 20536 44736
rect 19567 44696 20536 44724
rect 19567 44693 19579 44696
rect 19521 44687 19579 44693
rect 20530 44684 20536 44696
rect 20588 44684 20594 44736
rect 20622 44684 20628 44736
rect 20680 44724 20686 44736
rect 21085 44727 21143 44733
rect 21085 44724 21097 44727
rect 20680 44696 21097 44724
rect 20680 44684 20686 44696
rect 21085 44693 21097 44696
rect 21131 44693 21143 44727
rect 21085 44687 21143 44693
rect 22281 44727 22339 44733
rect 22281 44693 22293 44727
rect 22327 44724 22339 44727
rect 22462 44724 22468 44736
rect 22327 44696 22468 44724
rect 22327 44693 22339 44696
rect 22281 44687 22339 44693
rect 22462 44684 22468 44696
rect 22520 44684 22526 44736
rect 22664 44724 22692 44832
rect 22741 44829 22753 44863
rect 22787 44829 22799 44863
rect 22741 44823 22799 44829
rect 22830 44820 22836 44872
rect 22888 44860 22894 44872
rect 23474 44860 23480 44872
rect 22888 44832 22933 44860
rect 23435 44832 23480 44860
rect 22888 44820 22894 44832
rect 23474 44820 23480 44832
rect 23532 44820 23538 44872
rect 23569 44863 23627 44869
rect 23569 44829 23581 44863
rect 23615 44860 23627 44863
rect 23934 44860 23940 44872
rect 23615 44832 23940 44860
rect 23615 44829 23627 44832
rect 23569 44823 23627 44829
rect 23934 44820 23940 44832
rect 23992 44820 23998 44872
rect 22848 44792 22876 44820
rect 24044 44792 24072 44900
rect 24854 44888 24860 44900
rect 24912 44888 24918 44940
rect 25222 44888 25228 44940
rect 25280 44928 25286 44940
rect 25976 44928 26004 44968
rect 26142 44956 26148 45008
rect 26200 44996 26206 45008
rect 28261 44999 28319 45005
rect 28261 44996 28273 44999
rect 26200 44968 28273 44996
rect 26200 44956 26206 44968
rect 28261 44965 28273 44968
rect 28307 44996 28319 44999
rect 28718 44996 28724 45008
rect 28307 44968 28724 44996
rect 28307 44965 28319 44968
rect 28261 44959 28319 44965
rect 28718 44956 28724 44968
rect 28776 44956 28782 45008
rect 26418 44928 26424 44940
rect 25280 44900 25728 44928
rect 25280 44888 25286 44900
rect 25590 44860 25596 44872
rect 25551 44832 25596 44860
rect 25590 44820 25596 44832
rect 25648 44820 25654 44872
rect 25700 44869 25728 44900
rect 25976 44900 26424 44928
rect 25685 44863 25743 44869
rect 25685 44829 25697 44863
rect 25731 44829 25743 44863
rect 25685 44823 25743 44829
rect 25774 44820 25780 44872
rect 25832 44860 25838 44872
rect 25976 44869 26004 44900
rect 26418 44888 26424 44900
rect 26476 44888 26482 44940
rect 27249 44931 27307 44937
rect 27249 44897 27261 44931
rect 27295 44928 27307 44931
rect 27798 44928 27804 44940
rect 27295 44900 27804 44928
rect 27295 44897 27307 44900
rect 27249 44891 27307 44897
rect 27798 44888 27804 44900
rect 27856 44888 27862 44940
rect 29932 44928 29960 45036
rect 34146 45024 34152 45036
rect 34204 45064 34210 45076
rect 34885 45067 34943 45073
rect 34885 45064 34897 45067
rect 34204 45036 34897 45064
rect 34204 45024 34210 45036
rect 34885 45033 34897 45036
rect 34931 45033 34943 45067
rect 34885 45027 34943 45033
rect 32122 44996 32128 45008
rect 32083 44968 32128 44996
rect 32122 44956 32128 44968
rect 32180 44956 32186 45008
rect 30558 44928 30564 44940
rect 29932 44900 30564 44928
rect 25961 44863 26019 44869
rect 25832 44832 25877 44860
rect 25832 44820 25838 44832
rect 25961 44829 25973 44863
rect 26007 44829 26019 44863
rect 26697 44863 26755 44869
rect 26697 44860 26709 44863
rect 25961 44823 26019 44829
rect 26068 44832 26709 44860
rect 22848 44764 24072 44792
rect 24857 44795 24915 44801
rect 24857 44761 24869 44795
rect 24903 44792 24915 44795
rect 25498 44792 25504 44804
rect 24903 44764 25504 44792
rect 24903 44761 24915 44764
rect 24857 44755 24915 44761
rect 25498 44752 25504 44764
rect 25556 44792 25562 44804
rect 26068 44792 26096 44832
rect 26697 44829 26709 44832
rect 26743 44829 26755 44863
rect 26697 44823 26755 44829
rect 27522 44820 27528 44872
rect 27580 44860 27586 44872
rect 27617 44863 27675 44869
rect 27617 44860 27629 44863
rect 27580 44832 27629 44860
rect 27580 44820 27586 44832
rect 27617 44829 27629 44832
rect 27663 44860 27675 44863
rect 27890 44860 27896 44872
rect 27663 44832 27896 44860
rect 27663 44829 27675 44832
rect 27617 44823 27675 44829
rect 27890 44820 27896 44832
rect 27948 44820 27954 44872
rect 28074 44860 28080 44872
rect 28035 44832 28080 44860
rect 28074 44820 28080 44832
rect 28132 44820 28138 44872
rect 28997 44863 29055 44869
rect 28997 44829 29009 44863
rect 29043 44860 29055 44863
rect 29086 44860 29092 44872
rect 29043 44832 29092 44860
rect 29043 44829 29055 44832
rect 28997 44823 29055 44829
rect 29086 44820 29092 44832
rect 29144 44820 29150 44872
rect 29181 44863 29239 44869
rect 29181 44829 29193 44863
rect 29227 44860 29239 44863
rect 29362 44860 29368 44872
rect 29227 44832 29368 44860
rect 29227 44829 29239 44832
rect 29181 44823 29239 44829
rect 29362 44820 29368 44832
rect 29420 44820 29426 44872
rect 29822 44860 29828 44872
rect 29564 44832 29828 44860
rect 27430 44792 27436 44804
rect 25556 44764 26096 44792
rect 27391 44764 27436 44792
rect 25556 44752 25562 44764
rect 27430 44752 27436 44764
rect 27488 44752 27494 44804
rect 29564 44792 29592 44832
rect 29822 44820 29828 44832
rect 29880 44820 29886 44872
rect 29932 44869 29960 44900
rect 30558 44888 30564 44900
rect 30616 44888 30622 44940
rect 32490 44888 32496 44940
rect 32548 44928 32554 44940
rect 32861 44931 32919 44937
rect 32861 44928 32873 44931
rect 32548 44900 32873 44928
rect 32548 44888 32554 44900
rect 32861 44897 32873 44900
rect 32907 44897 32919 44931
rect 32861 44891 32919 44897
rect 29917 44863 29975 44869
rect 29917 44829 29929 44863
rect 29963 44829 29975 44863
rect 29917 44823 29975 44829
rect 30101 44863 30159 44869
rect 30101 44829 30113 44863
rect 30147 44860 30159 44863
rect 30282 44860 30288 44872
rect 30147 44832 30288 44860
rect 30147 44829 30159 44832
rect 30101 44823 30159 44829
rect 30282 44820 30288 44832
rect 30340 44860 30346 44872
rect 30926 44860 30932 44872
rect 30340 44832 30932 44860
rect 30340 44820 30346 44832
rect 30926 44820 30932 44832
rect 30984 44860 30990 44872
rect 32033 44863 32091 44869
rect 32033 44860 32045 44863
rect 30984 44832 32045 44860
rect 30984 44820 30990 44832
rect 32033 44829 32045 44832
rect 32079 44829 32091 44863
rect 32033 44823 32091 44829
rect 32217 44863 32275 44869
rect 32217 44829 32229 44863
rect 32263 44860 32275 44863
rect 32953 44863 33011 44869
rect 32953 44860 32965 44863
rect 32263 44832 32965 44860
rect 32263 44829 32275 44832
rect 32217 44823 32275 44829
rect 32953 44829 32965 44832
rect 32999 44860 33011 44863
rect 33134 44860 33140 44872
rect 32999 44832 33140 44860
rect 32999 44829 33011 44832
rect 32953 44823 33011 44829
rect 28920 44764 29592 44792
rect 28920 44736 28948 44764
rect 29638 44752 29644 44804
rect 29696 44792 29702 44804
rect 29733 44795 29791 44801
rect 29733 44792 29745 44795
rect 29696 44764 29745 44792
rect 29696 44752 29702 44764
rect 29733 44761 29745 44764
rect 29779 44761 29791 44795
rect 29733 44755 29791 44761
rect 30650 44752 30656 44804
rect 30708 44792 30714 44804
rect 31021 44795 31079 44801
rect 31021 44792 31033 44795
rect 30708 44764 31033 44792
rect 30708 44752 30714 44764
rect 31021 44761 31033 44764
rect 31067 44761 31079 44795
rect 32048 44792 32076 44823
rect 33134 44820 33140 44832
rect 33192 44860 33198 44872
rect 33502 44860 33508 44872
rect 33192 44832 33508 44860
rect 33192 44820 33198 44832
rect 33502 44820 33508 44832
rect 33560 44820 33566 44872
rect 33594 44820 33600 44872
rect 33652 44860 33658 44872
rect 33652 44832 33697 44860
rect 33652 44820 33658 44832
rect 33226 44792 33232 44804
rect 32048 44764 33232 44792
rect 31021 44755 31079 44761
rect 33226 44752 33232 44764
rect 33284 44752 33290 44804
rect 22738 44724 22744 44736
rect 22664 44696 22744 44724
rect 22738 44684 22744 44696
rect 22796 44724 22802 44736
rect 23014 44724 23020 44736
rect 22796 44696 23020 44724
rect 22796 44684 22802 44696
rect 23014 44684 23020 44696
rect 23072 44684 23078 44736
rect 25314 44724 25320 44736
rect 25275 44696 25320 44724
rect 25314 44684 25320 44696
rect 25372 44684 25378 44736
rect 25682 44684 25688 44736
rect 25740 44724 25746 44736
rect 28902 44724 28908 44736
rect 25740 44696 28908 44724
rect 25740 44684 25746 44696
rect 28902 44684 28908 44696
rect 28960 44684 28966 44736
rect 29089 44727 29147 44733
rect 29089 44693 29101 44727
rect 29135 44724 29147 44727
rect 30006 44724 30012 44736
rect 29135 44696 30012 44724
rect 29135 44693 29147 44696
rect 29089 44687 29147 44693
rect 30006 44684 30012 44696
rect 30064 44684 30070 44736
rect 31294 44724 31300 44736
rect 31255 44696 31300 44724
rect 31294 44684 31300 44696
rect 31352 44684 31358 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 21450 44480 21456 44532
rect 21508 44520 21514 44532
rect 22830 44520 22836 44532
rect 21508 44492 22836 44520
rect 21508 44480 21514 44492
rect 22830 44480 22836 44492
rect 22888 44480 22894 44532
rect 23474 44480 23480 44532
rect 23532 44520 23538 44532
rect 24302 44520 24308 44532
rect 23532 44492 24308 44520
rect 23532 44480 23538 44492
rect 24302 44480 24308 44492
rect 24360 44480 24366 44532
rect 25317 44523 25375 44529
rect 25317 44489 25329 44523
rect 25363 44520 25375 44523
rect 25682 44520 25688 44532
rect 25363 44492 25688 44520
rect 25363 44489 25375 44492
rect 25317 44483 25375 44489
rect 25682 44480 25688 44492
rect 25740 44520 25746 44532
rect 25740 44492 29776 44520
rect 25740 44480 25746 44492
rect 20438 44452 20444 44464
rect 20399 44424 20444 44452
rect 20438 44412 20444 44424
rect 20496 44412 20502 44464
rect 21082 44452 21088 44464
rect 20916 44424 21088 44452
rect 18690 44344 18696 44396
rect 18748 44384 18754 44396
rect 20916 44393 20944 44424
rect 21082 44412 21088 44424
rect 21140 44412 21146 44464
rect 21177 44455 21235 44461
rect 21177 44421 21189 44455
rect 21223 44452 21235 44455
rect 29638 44452 29644 44464
rect 21223 44424 29644 44452
rect 21223 44421 21235 44424
rect 21177 44415 21235 44421
rect 19245 44387 19303 44393
rect 19245 44384 19257 44387
rect 18748 44356 19257 44384
rect 18748 44344 18754 44356
rect 19245 44353 19257 44356
rect 19291 44384 19303 44387
rect 20901 44387 20959 44393
rect 19291 44356 20484 44384
rect 19291 44353 19303 44356
rect 19245 44347 19303 44353
rect 19426 44316 19432 44328
rect 19387 44288 19432 44316
rect 19426 44276 19432 44288
rect 19484 44276 19490 44328
rect 19061 44183 19119 44189
rect 19061 44149 19073 44183
rect 19107 44180 19119 44183
rect 19150 44180 19156 44192
rect 19107 44152 19156 44180
rect 19107 44149 19119 44152
rect 19061 44143 19119 44149
rect 19150 44140 19156 44152
rect 19208 44140 19214 44192
rect 20456 44180 20484 44356
rect 20901 44353 20913 44387
rect 20947 44353 20959 44387
rect 20901 44347 20959 44353
rect 20993 44387 21051 44393
rect 20993 44353 21005 44387
rect 21039 44353 21051 44387
rect 22002 44384 22008 44396
rect 21963 44356 22008 44384
rect 20993 44347 21051 44353
rect 20530 44276 20536 44328
rect 20588 44316 20594 44328
rect 21008 44316 21036 44347
rect 22002 44344 22008 44356
rect 22060 44344 22066 44396
rect 22186 44344 22192 44396
rect 22244 44384 22250 44396
rect 22741 44387 22799 44393
rect 22244 44356 22337 44384
rect 22244 44344 22250 44356
rect 22741 44353 22753 44387
rect 22787 44384 22799 44387
rect 22830 44384 22836 44396
rect 22787 44356 22836 44384
rect 22787 44353 22799 44356
rect 22741 44347 22799 44353
rect 22830 44344 22836 44356
rect 22888 44344 22894 44396
rect 22925 44387 22983 44393
rect 22925 44353 22937 44387
rect 22971 44353 22983 44387
rect 22925 44347 22983 44353
rect 20588 44288 21036 44316
rect 20588 44276 20594 44288
rect 21008 44248 21036 44288
rect 21726 44276 21732 44328
rect 21784 44316 21790 44328
rect 22204 44316 22232 44344
rect 21784 44288 22232 44316
rect 21784 44276 21790 44288
rect 22278 44276 22284 44328
rect 22336 44316 22342 44328
rect 22940 44316 22968 44347
rect 23750 44344 23756 44396
rect 23808 44384 23814 44396
rect 24121 44387 24179 44393
rect 24121 44384 24133 44387
rect 23808 44356 24133 44384
rect 23808 44344 23814 44356
rect 24121 44353 24133 44356
rect 24167 44384 24179 44387
rect 24210 44384 24216 44396
rect 24167 44356 24216 44384
rect 24167 44353 24179 44356
rect 24121 44347 24179 44353
rect 24210 44344 24216 44356
rect 24268 44344 24274 44396
rect 24305 44387 24363 44393
rect 24305 44353 24317 44387
rect 24351 44384 24363 44387
rect 24578 44384 24584 44396
rect 24351 44356 24584 44384
rect 24351 44353 24363 44356
rect 24305 44347 24363 44353
rect 22336 44288 22968 44316
rect 22336 44276 22342 44288
rect 23658 44276 23664 44328
rect 23716 44316 23722 44328
rect 24320 44316 24348 44347
rect 24578 44344 24584 44356
rect 24636 44344 24642 44396
rect 25130 44384 25136 44396
rect 25091 44356 25136 44384
rect 25130 44344 25136 44356
rect 25188 44344 25194 44396
rect 25409 44387 25467 44393
rect 25409 44353 25421 44387
rect 25455 44384 25467 44387
rect 25958 44384 25964 44396
rect 25455 44356 25964 44384
rect 25455 44353 25467 44356
rect 25409 44347 25467 44353
rect 25958 44344 25964 44356
rect 26016 44344 26022 44396
rect 26252 44393 26280 44424
rect 26237 44387 26295 44393
rect 26237 44353 26249 44387
rect 26283 44353 26295 44387
rect 26694 44384 26700 44396
rect 26237 44347 26295 44353
rect 26344 44356 26700 44384
rect 23716 44288 24348 44316
rect 24489 44319 24547 44325
rect 23716 44276 23722 44288
rect 24489 44285 24501 44319
rect 24535 44316 24547 44319
rect 26344 44316 26372 44356
rect 26694 44344 26700 44356
rect 26752 44384 26758 44396
rect 27249 44387 27307 44393
rect 27249 44384 27261 44387
rect 26752 44356 27261 44384
rect 26752 44344 26758 44356
rect 27249 44353 27261 44356
rect 27295 44353 27307 44387
rect 27249 44347 27307 44353
rect 27433 44387 27491 44393
rect 27433 44353 27445 44387
rect 27479 44353 27491 44387
rect 27890 44384 27896 44396
rect 27851 44356 27896 44384
rect 27433 44347 27491 44353
rect 24535 44288 26372 44316
rect 26513 44319 26571 44325
rect 24535 44285 24547 44288
rect 24489 44279 24547 44285
rect 26513 44285 26525 44319
rect 26559 44316 26571 44319
rect 27154 44316 27160 44328
rect 26559 44288 27160 44316
rect 26559 44285 26571 44288
rect 26513 44279 26571 44285
rect 27154 44276 27160 44288
rect 27212 44276 27218 44328
rect 27448 44316 27476 44347
rect 27890 44344 27896 44356
rect 27948 44344 27954 44396
rect 28092 44393 28120 44424
rect 28077 44387 28135 44393
rect 28077 44353 28089 44387
rect 28123 44353 28135 44387
rect 28902 44384 28908 44396
rect 28863 44356 28908 44384
rect 28077 44347 28135 44353
rect 28902 44344 28908 44356
rect 28960 44344 28966 44396
rect 29104 44393 29132 44424
rect 29638 44412 29644 44424
rect 29696 44412 29702 44464
rect 29748 44452 29776 44492
rect 29822 44480 29828 44532
rect 29880 44520 29886 44532
rect 32306 44520 32312 44532
rect 29880 44492 32312 44520
rect 29880 44480 29886 44492
rect 32306 44480 32312 44492
rect 32364 44480 32370 44532
rect 34146 44480 34152 44532
rect 34204 44480 34210 44532
rect 31846 44452 31852 44464
rect 29748 44424 31852 44452
rect 29089 44387 29147 44393
rect 29089 44353 29101 44387
rect 29135 44353 29147 44387
rect 29546 44384 29552 44396
rect 29507 44356 29552 44384
rect 29089 44347 29147 44353
rect 29546 44344 29552 44356
rect 29604 44344 29610 44396
rect 29748 44393 29776 44424
rect 31846 44412 31852 44424
rect 31904 44412 31910 44464
rect 34164 44452 34192 44480
rect 32508 44424 34192 44452
rect 29733 44387 29791 44393
rect 29733 44353 29745 44387
rect 29779 44353 29791 44387
rect 30282 44384 30288 44396
rect 30243 44356 30288 44384
rect 29733 44347 29791 44353
rect 30282 44344 30288 44356
rect 30340 44344 30346 44396
rect 30469 44387 30527 44393
rect 30469 44353 30481 44387
rect 30515 44384 30527 44387
rect 31110 44384 31116 44396
rect 30515 44356 31116 44384
rect 30515 44353 30527 44356
rect 30469 44347 30527 44353
rect 31110 44344 31116 44356
rect 31168 44344 31174 44396
rect 31297 44387 31355 44393
rect 31297 44353 31309 44387
rect 31343 44384 31355 44387
rect 31386 44384 31392 44396
rect 31343 44356 31392 44384
rect 31343 44353 31355 44356
rect 31297 44347 31355 44353
rect 31386 44344 31392 44356
rect 31444 44384 31450 44396
rect 32508 44393 32536 44424
rect 34422 44412 34428 44464
rect 34480 44452 34486 44464
rect 34609 44455 34667 44461
rect 34609 44452 34621 44455
rect 34480 44424 34621 44452
rect 34480 44412 34486 44424
rect 34609 44421 34621 44424
rect 34655 44421 34667 44455
rect 34809 44455 34867 44461
rect 34809 44452 34821 44455
rect 34609 44415 34667 44421
rect 34716 44424 34821 44452
rect 32493 44387 32551 44393
rect 32493 44384 32505 44387
rect 31444 44356 32505 44384
rect 31444 44344 31450 44356
rect 32493 44353 32505 44356
rect 32539 44353 32551 44387
rect 32493 44347 32551 44353
rect 33318 44344 33324 44396
rect 33376 44384 33382 44396
rect 33413 44387 33471 44393
rect 33413 44384 33425 44387
rect 33376 44356 33425 44384
rect 33376 44344 33382 44356
rect 33413 44353 33425 44356
rect 33459 44353 33471 44387
rect 33413 44347 33471 44353
rect 27522 44316 27528 44328
rect 27435 44288 27528 44316
rect 27522 44276 27528 44288
rect 27580 44316 27586 44328
rect 30374 44316 30380 44328
rect 27580 44288 30380 44316
rect 27580 44276 27586 44288
rect 30374 44276 30380 44288
rect 30432 44276 30438 44328
rect 33226 44316 33232 44328
rect 33139 44288 33232 44316
rect 33226 44276 33232 44288
rect 33284 44276 33290 44328
rect 33428 44316 33456 44347
rect 33502 44344 33508 44396
rect 33560 44384 33566 44396
rect 33965 44387 34023 44393
rect 33965 44384 33977 44387
rect 33560 44356 33977 44384
rect 33560 44344 33566 44356
rect 33965 44353 33977 44356
rect 34011 44384 34023 44387
rect 34716 44384 34744 44424
rect 34809 44421 34821 44424
rect 34855 44421 34867 44455
rect 34809 44415 34867 44421
rect 34011 44356 34744 44384
rect 34011 44353 34023 44356
rect 33965 44347 34023 44353
rect 34422 44316 34428 44328
rect 33428 44288 34428 44316
rect 34422 44276 34428 44288
rect 34480 44276 34486 44328
rect 22002 44248 22008 44260
rect 21008 44220 22008 44248
rect 22002 44208 22008 44220
rect 22060 44248 22066 44260
rect 22833 44251 22891 44257
rect 22060 44220 22784 44248
rect 22060 44208 22066 44220
rect 21177 44183 21235 44189
rect 21177 44180 21189 44183
rect 20456 44152 21189 44180
rect 21177 44149 21189 44152
rect 21223 44149 21235 44183
rect 22186 44180 22192 44192
rect 22147 44152 22192 44180
rect 21177 44143 21235 44149
rect 22186 44140 22192 44152
rect 22244 44140 22250 44192
rect 22756 44180 22784 44220
rect 22833 44217 22845 44251
rect 22879 44248 22891 44251
rect 22879 44220 23888 44248
rect 22879 44217 22891 44220
rect 22833 44211 22891 44217
rect 23569 44183 23627 44189
rect 23569 44180 23581 44183
rect 22756 44152 23581 44180
rect 23569 44149 23581 44152
rect 23615 44180 23627 44183
rect 23658 44180 23664 44192
rect 23615 44152 23664 44180
rect 23615 44149 23627 44152
rect 23569 44143 23627 44149
rect 23658 44140 23664 44152
rect 23716 44140 23722 44192
rect 23860 44180 23888 44220
rect 23934 44208 23940 44260
rect 23992 44248 23998 44260
rect 29730 44248 29736 44260
rect 23992 44220 29736 44248
rect 23992 44208 23998 44220
rect 29730 44208 29736 44220
rect 29788 44208 29794 44260
rect 24118 44180 24124 44192
rect 23860 44152 24124 44180
rect 24118 44140 24124 44152
rect 24176 44140 24182 44192
rect 24946 44180 24952 44192
rect 24907 44152 24952 44180
rect 24946 44140 24952 44152
rect 25004 44140 25010 44192
rect 25222 44140 25228 44192
rect 25280 44180 25286 44192
rect 26329 44183 26387 44189
rect 26329 44180 26341 44183
rect 25280 44152 26341 44180
rect 25280 44140 25286 44152
rect 26329 44149 26341 44152
rect 26375 44149 26387 44183
rect 26329 44143 26387 44149
rect 26418 44140 26424 44192
rect 26476 44180 26482 44192
rect 26476 44152 26521 44180
rect 26476 44140 26482 44152
rect 27154 44140 27160 44192
rect 27212 44180 27218 44192
rect 27249 44183 27307 44189
rect 27249 44180 27261 44183
rect 27212 44152 27261 44180
rect 27212 44140 27218 44152
rect 27249 44149 27261 44152
rect 27295 44149 27307 44183
rect 28074 44180 28080 44192
rect 28035 44152 28080 44180
rect 27249 44143 27307 44149
rect 28074 44140 28080 44152
rect 28132 44140 28138 44192
rect 29086 44180 29092 44192
rect 29047 44152 29092 44180
rect 29086 44140 29092 44152
rect 29144 44140 29150 44192
rect 29362 44140 29368 44192
rect 29420 44180 29426 44192
rect 29641 44183 29699 44189
rect 29641 44180 29653 44183
rect 29420 44152 29653 44180
rect 29420 44140 29426 44152
rect 29641 44149 29653 44152
rect 29687 44149 29699 44183
rect 31018 44180 31024 44192
rect 30979 44152 31024 44180
rect 29641 44143 29699 44149
rect 31018 44140 31024 44152
rect 31076 44140 31082 44192
rect 32398 44180 32404 44192
rect 32359 44152 32404 44180
rect 32398 44140 32404 44152
rect 32456 44140 32462 44192
rect 33244 44180 33272 44276
rect 33870 44248 33876 44260
rect 33831 44220 33876 44248
rect 33870 44208 33876 44220
rect 33928 44208 33934 44260
rect 34793 44183 34851 44189
rect 34793 44180 34805 44183
rect 33244 44152 34805 44180
rect 34793 44149 34805 44152
rect 34839 44149 34851 44183
rect 34793 44143 34851 44149
rect 34977 44183 35035 44189
rect 34977 44149 34989 44183
rect 35023 44180 35035 44183
rect 35342 44180 35348 44192
rect 35023 44152 35348 44180
rect 35023 44149 35035 44152
rect 34977 44143 35035 44149
rect 35342 44140 35348 44152
rect 35400 44140 35406 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 20530 43936 20536 43988
rect 20588 43976 20594 43988
rect 21361 43979 21419 43985
rect 20588 43948 21036 43976
rect 20588 43936 20594 43948
rect 18417 43911 18475 43917
rect 18417 43877 18429 43911
rect 18463 43908 18475 43911
rect 21008 43908 21036 43948
rect 21361 43945 21373 43979
rect 21407 43976 21419 43979
rect 22186 43976 22192 43988
rect 21407 43948 22192 43976
rect 21407 43945 21419 43948
rect 21361 43939 21419 43945
rect 22186 43936 22192 43948
rect 22244 43936 22250 43988
rect 23842 43976 23848 43988
rect 23803 43948 23848 43976
rect 23842 43936 23848 43948
rect 23900 43936 23906 43988
rect 24302 43936 24308 43988
rect 24360 43976 24366 43988
rect 24360 43948 26188 43976
rect 24360 43936 24366 43948
rect 25961 43911 26019 43917
rect 25961 43908 25973 43911
rect 18463 43880 20944 43908
rect 21008 43880 25973 43908
rect 18463 43877 18475 43880
rect 18417 43871 18475 43877
rect 19426 43840 19432 43852
rect 18892 43812 19432 43840
rect 18690 43772 18696 43784
rect 18651 43744 18696 43772
rect 18690 43732 18696 43744
rect 18748 43732 18754 43784
rect 18892 43781 18920 43812
rect 19426 43800 19432 43812
rect 19484 43840 19490 43852
rect 20622 43840 20628 43852
rect 19484 43812 20628 43840
rect 19484 43800 19490 43812
rect 20088 43781 20116 43812
rect 20622 43800 20628 43812
rect 20680 43800 20686 43852
rect 20916 43840 20944 43880
rect 25961 43877 25973 43880
rect 26007 43877 26019 43911
rect 26160 43908 26188 43948
rect 26234 43936 26240 43988
rect 26292 43976 26298 43988
rect 29914 43976 29920 43988
rect 26292 43948 29920 43976
rect 26292 43936 26298 43948
rect 29914 43936 29920 43948
rect 29972 43936 29978 43988
rect 30558 43936 30564 43988
rect 30616 43976 30622 43988
rect 30837 43979 30895 43985
rect 30837 43976 30849 43979
rect 30616 43948 30849 43976
rect 30616 43936 30622 43948
rect 30837 43945 30849 43948
rect 30883 43976 30895 43979
rect 31202 43976 31208 43988
rect 30883 43948 31208 43976
rect 30883 43945 30895 43948
rect 30837 43939 30895 43945
rect 31202 43936 31208 43948
rect 31260 43976 31266 43988
rect 32677 43979 32735 43985
rect 32677 43976 32689 43979
rect 31260 43948 32689 43976
rect 31260 43936 31266 43948
rect 32677 43945 32689 43948
rect 32723 43945 32735 43979
rect 32677 43939 32735 43945
rect 33410 43936 33416 43988
rect 33468 43976 33474 43988
rect 33505 43979 33563 43985
rect 33505 43976 33517 43979
rect 33468 43948 33517 43976
rect 33468 43936 33474 43948
rect 33505 43945 33517 43948
rect 33551 43976 33563 43979
rect 33870 43976 33876 43988
rect 33551 43948 33876 43976
rect 33551 43945 33563 43948
rect 33505 43939 33563 43945
rect 33870 43936 33876 43948
rect 33928 43936 33934 43988
rect 26160 43880 28212 43908
rect 25961 43871 26019 43877
rect 21910 43840 21916 43852
rect 20916 43812 21916 43840
rect 21910 43800 21916 43812
rect 21968 43840 21974 43852
rect 25869 43843 25927 43849
rect 25869 43840 25881 43843
rect 21968 43812 25881 43840
rect 21968 43800 21974 43812
rect 25869 43809 25881 43812
rect 25915 43840 25927 43843
rect 26145 43843 26203 43849
rect 25915 43812 26096 43840
rect 25915 43809 25927 43812
rect 25869 43803 25927 43809
rect 18877 43775 18935 43781
rect 18877 43741 18889 43775
rect 18923 43741 18935 43775
rect 18877 43735 18935 43741
rect 20073 43775 20131 43781
rect 20073 43741 20085 43775
rect 20119 43741 20131 43775
rect 20346 43772 20352 43784
rect 20307 43744 20352 43772
rect 20073 43735 20131 43741
rect 20346 43732 20352 43744
rect 20404 43732 20410 43784
rect 20533 43775 20591 43781
rect 20533 43741 20545 43775
rect 20579 43772 20591 43775
rect 20993 43775 21051 43781
rect 20993 43772 21005 43775
rect 20579 43744 21005 43772
rect 20579 43741 20591 43744
rect 20533 43735 20591 43741
rect 20993 43741 21005 43744
rect 21039 43741 21051 43775
rect 20993 43735 21051 43741
rect 21177 43775 21235 43781
rect 21177 43741 21189 43775
rect 21223 43741 21235 43775
rect 21177 43735 21235 43741
rect 20165 43707 20223 43713
rect 20165 43673 20177 43707
rect 20211 43673 20223 43707
rect 20165 43667 20223 43673
rect 20257 43707 20315 43713
rect 20257 43673 20269 43707
rect 20303 43704 20315 43707
rect 20438 43704 20444 43716
rect 20303 43676 20444 43704
rect 20303 43673 20315 43676
rect 20257 43667 20315 43673
rect 18598 43636 18604 43648
rect 18559 43608 18604 43636
rect 18598 43596 18604 43608
rect 18656 43596 18662 43648
rect 19334 43596 19340 43648
rect 19392 43636 19398 43648
rect 19889 43639 19947 43645
rect 19889 43636 19901 43639
rect 19392 43608 19901 43636
rect 19392 43596 19398 43608
rect 19889 43605 19901 43608
rect 19935 43605 19947 43639
rect 20180 43636 20208 43667
rect 20438 43664 20444 43676
rect 20496 43704 20502 43716
rect 20622 43704 20628 43716
rect 20496 43676 20628 43704
rect 20496 43664 20502 43676
rect 20622 43664 20628 43676
rect 20680 43664 20686 43716
rect 21192 43704 21220 43735
rect 21358 43732 21364 43784
rect 21416 43772 21422 43784
rect 21453 43775 21511 43781
rect 21453 43772 21465 43775
rect 21416 43744 21465 43772
rect 21416 43732 21422 43744
rect 21453 43741 21465 43744
rect 21499 43741 21511 43775
rect 23290 43772 23296 43784
rect 21453 43735 21511 43741
rect 21560 43744 23296 43772
rect 21560 43704 21588 43744
rect 23290 43732 23296 43744
rect 23348 43732 23354 43784
rect 23661 43775 23719 43781
rect 23661 43741 23673 43775
rect 23707 43766 23719 43775
rect 24029 43775 24087 43781
rect 23707 43741 23736 43766
rect 23661 43735 23736 43741
rect 24029 43741 24041 43775
rect 24075 43772 24087 43775
rect 24302 43772 24308 43784
rect 24075 43744 24308 43772
rect 24075 43741 24087 43744
rect 24029 43735 24087 43741
rect 21192 43676 21588 43704
rect 21818 43664 21824 43716
rect 21876 43704 21882 43716
rect 22097 43707 22155 43713
rect 22097 43704 22109 43707
rect 21876 43676 22109 43704
rect 21876 43664 21882 43676
rect 22097 43673 22109 43676
rect 22143 43673 22155 43707
rect 22097 43667 22155 43673
rect 22370 43664 22376 43716
rect 22428 43704 22434 43716
rect 22465 43707 22523 43713
rect 22465 43704 22477 43707
rect 22428 43676 22477 43704
rect 22428 43664 22434 43676
rect 22465 43673 22477 43676
rect 22511 43673 22523 43707
rect 23708 43704 23736 43735
rect 24302 43732 24308 43744
rect 24360 43732 24366 43784
rect 25590 43772 25596 43784
rect 25551 43744 25596 43772
rect 25590 43732 25596 43744
rect 25648 43732 25654 43784
rect 25774 43732 25780 43784
rect 25832 43772 25838 43784
rect 25958 43772 25964 43784
rect 25832 43744 25964 43772
rect 25832 43732 25838 43744
rect 25958 43732 25964 43744
rect 26016 43732 26022 43784
rect 26068 43772 26096 43812
rect 26145 43809 26157 43843
rect 26191 43840 26203 43843
rect 27709 43843 27767 43849
rect 27709 43840 27721 43843
rect 26191 43812 27721 43840
rect 26191 43809 26203 43812
rect 26145 43803 26203 43809
rect 27709 43809 27721 43812
rect 27755 43809 27767 43843
rect 27709 43803 27767 43809
rect 28184 43840 28212 43880
rect 29086 43868 29092 43920
rect 29144 43908 29150 43920
rect 30101 43911 30159 43917
rect 30101 43908 30113 43911
rect 29144 43880 30113 43908
rect 29144 43868 29150 43880
rect 30101 43877 30113 43880
rect 30147 43877 30159 43911
rect 31110 43908 31116 43920
rect 30101 43871 30159 43877
rect 30760 43880 31116 43908
rect 29178 43840 29184 43852
rect 28184 43812 29184 43840
rect 26234 43772 26240 43784
rect 26068 43744 26240 43772
rect 26234 43732 26240 43744
rect 26292 43732 26298 43784
rect 26421 43775 26479 43781
rect 26421 43741 26433 43775
rect 26467 43772 26479 43775
rect 26510 43772 26516 43784
rect 26467 43744 26516 43772
rect 26467 43741 26479 43744
rect 26421 43735 26479 43741
rect 26510 43732 26516 43744
rect 26568 43732 26574 43784
rect 27154 43772 27160 43784
rect 27115 43744 27160 43772
rect 27154 43732 27160 43744
rect 27212 43732 27218 43784
rect 27249 43775 27307 43781
rect 27249 43741 27261 43775
rect 27295 43741 27307 43775
rect 27249 43735 27307 43741
rect 27433 43775 27491 43781
rect 27433 43741 27445 43775
rect 27479 43741 27491 43775
rect 27433 43735 27491 43741
rect 27525 43775 27583 43781
rect 27525 43741 27537 43775
rect 27571 43772 27583 43775
rect 27982 43772 27988 43784
rect 27571 43744 27988 43772
rect 27571 43741 27583 43744
rect 27525 43735 27583 43741
rect 23708 43676 24072 43704
rect 22465 43667 22523 43673
rect 24044 43648 24072 43676
rect 24118 43664 24124 43716
rect 24176 43704 24182 43716
rect 27264 43704 27292 43735
rect 24176 43676 27292 43704
rect 27448 43704 27476 43735
rect 27982 43732 27988 43744
rect 28040 43732 28046 43784
rect 28184 43781 28212 43812
rect 29178 43800 29184 43812
rect 29236 43800 29242 43852
rect 30760 43849 30788 43880
rect 31110 43868 31116 43880
rect 31168 43868 31174 43920
rect 31846 43908 31852 43920
rect 31807 43880 31852 43908
rect 31846 43868 31852 43880
rect 31904 43868 31910 43920
rect 30745 43843 30803 43849
rect 30745 43840 30757 43843
rect 29564 43812 30757 43840
rect 28169 43775 28227 43781
rect 28169 43741 28181 43775
rect 28215 43741 28227 43775
rect 28169 43735 28227 43741
rect 28258 43732 28264 43784
rect 28316 43772 28322 43784
rect 28353 43775 28411 43781
rect 28353 43772 28365 43775
rect 28316 43744 28365 43772
rect 28316 43732 28322 43744
rect 28353 43741 28365 43744
rect 28399 43741 28411 43775
rect 28353 43735 28411 43741
rect 28626 43732 28632 43784
rect 28684 43772 28690 43784
rect 28813 43775 28871 43781
rect 28813 43772 28825 43775
rect 28684 43744 28825 43772
rect 28684 43732 28690 43744
rect 28813 43741 28825 43744
rect 28859 43741 28871 43775
rect 28813 43735 28871 43741
rect 28997 43775 29055 43781
rect 28997 43741 29009 43775
rect 29043 43772 29055 43775
rect 29564 43772 29592 43812
rect 30745 43809 30757 43812
rect 30791 43809 30803 43843
rect 34974 43840 34980 43852
rect 34935 43812 34980 43840
rect 30745 43803 30803 43809
rect 34974 43800 34980 43812
rect 35032 43800 35038 43852
rect 29043 43744 29592 43772
rect 29043 43741 29055 43744
rect 28997 43735 29055 43741
rect 29822 43732 29828 43784
rect 29880 43772 29886 43784
rect 29917 43775 29975 43781
rect 29917 43772 29929 43775
rect 29880 43744 29929 43772
rect 29880 43732 29886 43744
rect 29917 43741 29929 43744
rect 29963 43741 29975 43775
rect 29917 43735 29975 43741
rect 30006 43732 30012 43784
rect 30064 43772 30070 43784
rect 30193 43775 30251 43781
rect 30064 43744 30157 43772
rect 30064 43732 30070 43744
rect 30193 43741 30205 43775
rect 30239 43772 30251 43775
rect 30650 43772 30656 43784
rect 30239 43744 30656 43772
rect 30239 43741 30251 43744
rect 30193 43735 30251 43741
rect 30650 43732 30656 43744
rect 30708 43732 30714 43784
rect 31018 43772 31024 43784
rect 30979 43744 31024 43772
rect 31018 43732 31024 43744
rect 31076 43732 31082 43784
rect 31110 43732 31116 43784
rect 31168 43772 31174 43784
rect 31294 43772 31300 43784
rect 31168 43744 31300 43772
rect 31168 43732 31174 43744
rect 31294 43732 31300 43744
rect 31352 43772 31358 43784
rect 31665 43775 31723 43781
rect 31665 43772 31677 43775
rect 31352 43744 31677 43772
rect 31352 43732 31358 43744
rect 31665 43741 31677 43744
rect 31711 43741 31723 43775
rect 31665 43735 31723 43741
rect 32398 43732 32404 43784
rect 32456 43772 32462 43784
rect 34885 43775 34943 43781
rect 34885 43772 34897 43775
rect 32456 43744 34897 43772
rect 32456 43732 32462 43744
rect 34885 43741 34897 43744
rect 34931 43741 34943 43775
rect 34885 43735 34943 43741
rect 35069 43775 35127 43781
rect 35069 43741 35081 43775
rect 35115 43772 35127 43775
rect 35342 43772 35348 43784
rect 35115 43744 35348 43772
rect 35115 43741 35127 43744
rect 35069 43735 35127 43741
rect 35342 43732 35348 43744
rect 35400 43732 35406 43784
rect 29454 43704 29460 43716
rect 27448 43676 29460 43704
rect 24176 43664 24182 43676
rect 29454 43664 29460 43676
rect 29512 43664 29518 43716
rect 30024 43704 30052 43732
rect 30466 43704 30472 43716
rect 30024 43676 30472 43704
rect 30466 43664 30472 43676
rect 30524 43664 30530 43716
rect 32582 43704 32588 43716
rect 32543 43676 32588 43704
rect 32582 43664 32588 43676
rect 32640 43664 32646 43716
rect 33318 43664 33324 43716
rect 33376 43704 33382 43716
rect 33781 43707 33839 43713
rect 33781 43704 33793 43707
rect 33376 43676 33793 43704
rect 33376 43664 33382 43676
rect 33781 43673 33793 43676
rect 33827 43673 33839 43707
rect 33781 43667 33839 43673
rect 22554 43636 22560 43648
rect 20180 43608 22560 43636
rect 19889 43599 19947 43605
rect 22554 43596 22560 43608
rect 22612 43596 22618 43648
rect 23474 43636 23480 43648
rect 23435 43608 23480 43636
rect 23474 43596 23480 43608
rect 23532 43596 23538 43648
rect 24026 43596 24032 43648
rect 24084 43596 24090 43648
rect 24765 43639 24823 43645
rect 24765 43605 24777 43639
rect 24811 43636 24823 43639
rect 25038 43636 25044 43648
rect 24811 43608 25044 43636
rect 24811 43605 24823 43608
rect 24765 43599 24823 43605
rect 25038 43596 25044 43608
rect 25096 43596 25102 43648
rect 28258 43636 28264 43648
rect 28219 43608 28264 43636
rect 28258 43596 28264 43608
rect 28316 43596 28322 43648
rect 28902 43636 28908 43648
rect 28863 43608 28908 43636
rect 28902 43596 28908 43608
rect 28960 43596 28966 43648
rect 29730 43636 29736 43648
rect 29691 43608 29736 43636
rect 29730 43596 29736 43608
rect 29788 43596 29794 43648
rect 31205 43639 31263 43645
rect 31205 43605 31217 43639
rect 31251 43636 31263 43639
rect 31478 43636 31484 43648
rect 31251 43608 31484 43636
rect 31251 43605 31263 43608
rect 31205 43599 31263 43605
rect 31478 43596 31484 43608
rect 31536 43596 31542 43648
rect 35621 43639 35679 43645
rect 35621 43605 35633 43639
rect 35667 43636 35679 43639
rect 35802 43636 35808 43648
rect 35667 43608 35808 43636
rect 35667 43605 35679 43608
rect 35621 43599 35679 43605
rect 35802 43596 35808 43608
rect 35860 43596 35866 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 23385 43435 23443 43441
rect 23385 43432 23397 43435
rect 20456 43404 23397 43432
rect 18598 43324 18604 43376
rect 18656 43364 18662 43376
rect 18656 43336 20208 43364
rect 18656 43324 18662 43336
rect 18892 43305 18920 43336
rect 18509 43299 18567 43305
rect 18509 43265 18521 43299
rect 18555 43265 18567 43299
rect 18509 43259 18567 43265
rect 18877 43299 18935 43305
rect 18877 43265 18889 43299
rect 18923 43265 18935 43299
rect 18877 43259 18935 43265
rect 19061 43299 19119 43305
rect 19061 43265 19073 43299
rect 19107 43296 19119 43299
rect 19978 43296 19984 43308
rect 19107 43268 19984 43296
rect 19107 43265 19119 43268
rect 19061 43259 19119 43265
rect 18524 43228 18552 43259
rect 19978 43256 19984 43268
rect 20036 43256 20042 43308
rect 20180 43305 20208 43336
rect 20073 43299 20131 43305
rect 20073 43265 20085 43299
rect 20119 43265 20131 43299
rect 20073 43259 20131 43265
rect 20165 43299 20223 43305
rect 20165 43265 20177 43299
rect 20211 43265 20223 43299
rect 20165 43259 20223 43265
rect 19150 43228 19156 43240
rect 18524 43200 19156 43228
rect 19150 43188 19156 43200
rect 19208 43228 19214 43240
rect 20088 43228 20116 43259
rect 20254 43256 20260 43308
rect 20312 43296 20318 43308
rect 20456 43305 20484 43404
rect 23385 43401 23397 43404
rect 23431 43401 23443 43435
rect 24118 43432 24124 43444
rect 23385 43395 23443 43401
rect 23492 43404 24124 43432
rect 20901 43367 20959 43373
rect 20901 43333 20913 43367
rect 20947 43364 20959 43367
rect 22094 43364 22100 43376
rect 20947 43336 22100 43364
rect 20947 43333 20959 43336
rect 20901 43327 20959 43333
rect 22094 43324 22100 43336
rect 22152 43364 22158 43376
rect 22278 43364 22284 43376
rect 22152 43336 22284 43364
rect 22152 43324 22158 43336
rect 22278 43324 22284 43336
rect 22336 43324 22342 43376
rect 23492 43364 23520 43404
rect 24118 43392 24124 43404
rect 24176 43392 24182 43444
rect 25409 43435 25467 43441
rect 25409 43401 25421 43435
rect 25455 43432 25467 43435
rect 25590 43432 25596 43444
rect 25455 43404 25596 43432
rect 25455 43401 25467 43404
rect 25409 43395 25467 43401
rect 25590 43392 25596 43404
rect 25648 43392 25654 43444
rect 26510 43392 26516 43444
rect 26568 43432 26574 43444
rect 26568 43404 28212 43432
rect 26568 43392 26574 43404
rect 22756 43336 23520 43364
rect 23661 43367 23719 43373
rect 20441 43299 20499 43305
rect 20312 43268 20357 43296
rect 20312 43256 20318 43268
rect 20441 43265 20453 43299
rect 20487 43265 20499 43299
rect 20441 43259 20499 43265
rect 20456 43228 20484 43259
rect 20990 43256 20996 43308
rect 21048 43296 21054 43308
rect 21085 43299 21143 43305
rect 21085 43296 21097 43299
rect 21048 43268 21097 43296
rect 21048 43256 21054 43268
rect 21085 43265 21097 43268
rect 21131 43265 21143 43299
rect 21085 43259 21143 43265
rect 21174 43256 21180 43308
rect 21232 43296 21238 43308
rect 22462 43296 22468 43308
rect 21232 43268 21277 43296
rect 22423 43268 22468 43296
rect 21232 43256 21238 43268
rect 22462 43256 22468 43268
rect 22520 43256 22526 43308
rect 22756 43305 22784 43336
rect 23661 43333 23673 43367
rect 23707 43364 23719 43367
rect 24762 43364 24768 43376
rect 23707 43336 24768 43364
rect 23707 43333 23719 43336
rect 23661 43327 23719 43333
rect 24762 43324 24768 43336
rect 24820 43324 24826 43376
rect 26326 43324 26332 43376
rect 26384 43364 26390 43376
rect 27309 43367 27367 43373
rect 27309 43364 27321 43367
rect 26384 43336 27321 43364
rect 26384 43324 26390 43336
rect 27309 43333 27321 43336
rect 27355 43333 27367 43367
rect 27522 43364 27528 43376
rect 27483 43336 27528 43364
rect 27309 43327 27367 43333
rect 27522 43324 27528 43336
rect 27580 43324 27586 43376
rect 28184 43373 28212 43404
rect 29178 43392 29184 43444
rect 29236 43432 29242 43444
rect 32122 43432 32128 43444
rect 29236 43404 32128 43432
rect 29236 43392 29242 43404
rect 32122 43392 32128 43404
rect 32180 43392 32186 43444
rect 28169 43367 28227 43373
rect 28169 43333 28181 43367
rect 28215 43333 28227 43367
rect 31205 43367 31263 43373
rect 31205 43364 31217 43367
rect 28169 43327 28227 43333
rect 30392 43336 31217 43364
rect 22557 43299 22615 43305
rect 22557 43265 22569 43299
rect 22603 43265 22615 43299
rect 22557 43259 22615 43265
rect 22741 43299 22799 43305
rect 22741 43265 22753 43299
rect 22787 43265 22799 43299
rect 22741 43259 22799 43265
rect 22833 43299 22891 43305
rect 22833 43265 22845 43299
rect 22879 43296 22891 43299
rect 22879 43268 23428 43296
rect 22879 43265 22891 43268
rect 22833 43259 22891 43265
rect 19208 43200 20116 43228
rect 20272 43200 20484 43228
rect 19208 43188 19214 43200
rect 19337 43163 19395 43169
rect 19337 43129 19349 43163
rect 19383 43160 19395 43163
rect 20272 43160 20300 43200
rect 19383 43132 20300 43160
rect 19383 43129 19395 43132
rect 19337 43123 19395 43129
rect 20346 43120 20352 43172
rect 20404 43160 20410 43172
rect 20901 43163 20959 43169
rect 20901 43160 20913 43163
rect 20404 43132 20913 43160
rect 20404 43120 20410 43132
rect 20901 43129 20913 43132
rect 20947 43129 20959 43163
rect 20901 43123 20959 43129
rect 22186 43120 22192 43172
rect 22244 43160 22250 43172
rect 22572 43160 22600 43259
rect 23400 43228 23428 43268
rect 23474 43256 23480 43308
rect 23532 43305 23538 43308
rect 23532 43299 23581 43305
rect 23532 43265 23535 43299
rect 23569 43265 23581 43299
rect 23750 43296 23756 43308
rect 23711 43268 23756 43296
rect 23532 43259 23581 43265
rect 23532 43256 23538 43259
rect 23750 43256 23756 43268
rect 23808 43256 23814 43308
rect 23934 43296 23940 43308
rect 23895 43268 23940 43296
rect 23934 43256 23940 43268
rect 23992 43256 23998 43308
rect 24029 43299 24087 43305
rect 24029 43265 24041 43299
rect 24075 43296 24087 43299
rect 24118 43296 24124 43308
rect 24075 43268 24124 43296
rect 24075 43265 24087 43268
rect 24029 43259 24087 43265
rect 24118 43256 24124 43268
rect 24176 43256 24182 43308
rect 24210 43256 24216 43308
rect 24268 43296 24274 43308
rect 24489 43299 24547 43305
rect 24489 43296 24501 43299
rect 24268 43268 24501 43296
rect 24268 43256 24274 43268
rect 24489 43265 24501 43268
rect 24535 43265 24547 43299
rect 24670 43296 24676 43308
rect 24631 43268 24676 43296
rect 24489 43259 24547 43265
rect 24670 43256 24676 43268
rect 24728 43256 24734 43308
rect 25498 43256 25504 43308
rect 25556 43296 25562 43308
rect 25593 43299 25651 43305
rect 25593 43296 25605 43299
rect 25556 43268 25605 43296
rect 25556 43256 25562 43268
rect 25593 43265 25605 43268
rect 25639 43265 25651 43299
rect 25593 43259 25651 43265
rect 25685 43299 25743 43305
rect 25685 43265 25697 43299
rect 25731 43296 25743 43299
rect 25774 43296 25780 43308
rect 25731 43268 25780 43296
rect 25731 43265 25743 43268
rect 25685 43259 25743 43265
rect 25774 43256 25780 43268
rect 25832 43256 25838 43308
rect 25869 43299 25927 43305
rect 25869 43265 25881 43299
rect 25915 43296 25927 43299
rect 25958 43296 25964 43308
rect 25915 43268 25964 43296
rect 25915 43265 25927 43268
rect 25869 43259 25927 43265
rect 25958 43256 25964 43268
rect 26016 43256 26022 43308
rect 28258 43296 28264 43308
rect 28219 43268 28264 43296
rect 28258 43256 28264 43268
rect 28316 43256 28322 43308
rect 28537 43299 28595 43305
rect 28997 43302 29055 43305
rect 28537 43265 28549 43299
rect 28583 43265 28595 43299
rect 28828 43299 29055 43302
rect 28828 43296 29009 43299
rect 28537 43259 28595 43265
rect 28644 43274 29009 43296
rect 28644 43268 28856 43274
rect 27062 43228 27068 43240
rect 23400 43200 23612 43228
rect 23584 43172 23612 43200
rect 25792 43200 27068 43228
rect 22244 43132 22600 43160
rect 22244 43120 22250 43132
rect 23566 43120 23572 43172
rect 23624 43120 23630 43172
rect 25590 43120 25596 43172
rect 25648 43160 25654 43172
rect 25792 43169 25820 43200
rect 27062 43188 27068 43200
rect 27120 43228 27126 43240
rect 28442 43228 28448 43240
rect 27120 43200 28448 43228
rect 27120 43188 27126 43200
rect 28442 43188 28448 43200
rect 28500 43188 28506 43240
rect 25777 43163 25835 43169
rect 25777 43160 25789 43163
rect 25648 43132 25789 43160
rect 25648 43120 25654 43132
rect 25777 43129 25789 43132
rect 25823 43129 25835 43163
rect 25777 43123 25835 43129
rect 26513 43163 26571 43169
rect 26513 43129 26525 43163
rect 26559 43160 26571 43163
rect 26602 43160 26608 43172
rect 26559 43132 26608 43160
rect 26559 43129 26571 43132
rect 26513 43123 26571 43129
rect 26602 43120 26608 43132
rect 26660 43120 26666 43172
rect 27154 43160 27160 43172
rect 27115 43132 27160 43160
rect 27154 43120 27160 43132
rect 27212 43120 27218 43172
rect 27246 43120 27252 43172
rect 27304 43160 27310 43172
rect 28258 43160 28264 43172
rect 27304 43132 28264 43160
rect 27304 43120 27310 43132
rect 28258 43120 28264 43132
rect 28316 43160 28322 43172
rect 28552 43160 28580 43259
rect 28316 43132 28580 43160
rect 28316 43120 28322 43132
rect 19242 43092 19248 43104
rect 19203 43064 19248 43092
rect 19242 43052 19248 43064
rect 19300 43052 19306 43104
rect 19426 43052 19432 43104
rect 19484 43092 19490 43104
rect 19797 43095 19855 43101
rect 19797 43092 19809 43095
rect 19484 43064 19809 43092
rect 19484 43052 19490 43064
rect 19797 43061 19809 43064
rect 19843 43061 19855 43095
rect 19797 43055 19855 43061
rect 22281 43095 22339 43101
rect 22281 43061 22293 43095
rect 22327 43092 22339 43095
rect 22554 43092 22560 43104
rect 22327 43064 22560 43092
rect 22327 43061 22339 43064
rect 22281 43055 22339 43061
rect 22554 43052 22560 43064
rect 22612 43052 22618 43104
rect 24673 43095 24731 43101
rect 24673 43061 24685 43095
rect 24719 43092 24731 43095
rect 24762 43092 24768 43104
rect 24719 43064 24768 43092
rect 24719 43061 24731 43064
rect 24673 43055 24731 43061
rect 24762 43052 24768 43064
rect 24820 43052 24826 43104
rect 26050 43052 26056 43104
rect 26108 43092 26114 43104
rect 27341 43095 27399 43101
rect 27341 43092 27353 43095
rect 26108 43064 27353 43092
rect 26108 43052 26114 43064
rect 27341 43061 27353 43064
rect 27387 43061 27399 43095
rect 27341 43055 27399 43061
rect 27890 43052 27896 43104
rect 27948 43092 27954 43104
rect 28644 43092 28672 43268
rect 28997 43265 29009 43274
rect 29043 43265 29055 43299
rect 29362 43296 29368 43308
rect 29323 43268 29368 43296
rect 28997 43259 29055 43265
rect 29362 43256 29368 43268
rect 29420 43256 29426 43308
rect 29454 43256 29460 43308
rect 29512 43296 29518 43308
rect 29733 43299 29791 43305
rect 29733 43296 29745 43299
rect 29512 43268 29745 43296
rect 29512 43256 29518 43268
rect 29733 43265 29745 43268
rect 29779 43265 29791 43299
rect 29733 43259 29791 43265
rect 29822 43120 29828 43172
rect 29880 43160 29886 43172
rect 30190 43160 30196 43172
rect 29880 43132 30196 43160
rect 29880 43120 29886 43132
rect 30190 43120 30196 43132
rect 30248 43120 30254 43172
rect 27948 43064 28672 43092
rect 27948 43052 27954 43064
rect 30006 43052 30012 43104
rect 30064 43092 30070 43104
rect 30392 43092 30420 43336
rect 31205 43333 31217 43336
rect 31251 43333 31263 43367
rect 32398 43364 32404 43376
rect 32359 43336 32404 43364
rect 31205 43327 31263 43333
rect 32398 43324 32404 43336
rect 32456 43324 32462 43376
rect 30469 43299 30527 43305
rect 30469 43265 30481 43299
rect 30515 43265 30527 43299
rect 33686 43296 33692 43308
rect 33647 43268 33692 43296
rect 30469 43259 30527 43265
rect 30484 43228 30512 43259
rect 33686 43256 33692 43268
rect 33744 43296 33750 43308
rect 35161 43299 35219 43305
rect 35161 43296 35173 43299
rect 33744 43268 35173 43296
rect 33744 43256 33750 43268
rect 35161 43265 35173 43268
rect 35207 43296 35219 43299
rect 35434 43296 35440 43308
rect 35207 43268 35440 43296
rect 35207 43265 35219 43268
rect 35161 43259 35219 43265
rect 35434 43256 35440 43268
rect 35492 43256 35498 43308
rect 31662 43228 31668 43240
rect 30484 43200 31668 43228
rect 31662 43188 31668 43200
rect 31720 43188 31726 43240
rect 33502 43188 33508 43240
rect 33560 43228 33566 43240
rect 33873 43231 33931 43237
rect 33873 43228 33885 43231
rect 33560 43200 33885 43228
rect 33560 43188 33566 43200
rect 33873 43197 33885 43200
rect 33919 43197 33931 43231
rect 33873 43191 33931 43197
rect 34701 43163 34759 43169
rect 34701 43129 34713 43163
rect 34747 43160 34759 43163
rect 35986 43160 35992 43172
rect 34747 43132 35992 43160
rect 34747 43129 34759 43132
rect 34701 43123 34759 43129
rect 35986 43120 35992 43132
rect 36044 43120 36050 43172
rect 30561 43095 30619 43101
rect 30561 43092 30573 43095
rect 30064 43064 30573 43092
rect 30064 43052 30070 43064
rect 30561 43061 30573 43064
rect 30607 43061 30619 43095
rect 31294 43092 31300 43104
rect 31255 43064 31300 43092
rect 30561 43055 30619 43061
rect 31294 43052 31300 43064
rect 31352 43052 31358 43104
rect 32674 43092 32680 43104
rect 32635 43064 32680 43092
rect 32674 43052 32680 43064
rect 32732 43052 32738 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 20254 42848 20260 42900
rect 20312 42888 20318 42900
rect 24670 42888 24676 42900
rect 20312 42860 24676 42888
rect 20312 42848 20318 42860
rect 24670 42848 24676 42860
rect 24728 42848 24734 42900
rect 25041 42891 25099 42897
rect 25041 42857 25053 42891
rect 25087 42888 25099 42891
rect 25498 42888 25504 42900
rect 25087 42860 25504 42888
rect 25087 42857 25099 42860
rect 25041 42851 25099 42857
rect 25498 42848 25504 42860
rect 25556 42848 25562 42900
rect 29914 42848 29920 42900
rect 29972 42888 29978 42900
rect 30009 42891 30067 42897
rect 30009 42888 30021 42891
rect 29972 42860 30021 42888
rect 29972 42848 29978 42860
rect 30009 42857 30021 42860
rect 30055 42888 30067 42891
rect 30282 42888 30288 42900
rect 30055 42860 30288 42888
rect 30055 42857 30067 42860
rect 30009 42851 30067 42857
rect 30282 42848 30288 42860
rect 30340 42848 30346 42900
rect 30650 42848 30656 42900
rect 30708 42888 30714 42900
rect 31205 42891 31263 42897
rect 31205 42888 31217 42891
rect 30708 42860 31217 42888
rect 30708 42848 30714 42860
rect 31205 42857 31217 42860
rect 31251 42857 31263 42891
rect 31205 42851 31263 42857
rect 31389 42891 31447 42897
rect 31389 42857 31401 42891
rect 31435 42857 31447 42891
rect 31389 42851 31447 42857
rect 21818 42780 21824 42832
rect 21876 42820 21882 42832
rect 25590 42820 25596 42832
rect 21876 42792 25596 42820
rect 21876 42780 21882 42792
rect 25590 42780 25596 42792
rect 25648 42780 25654 42832
rect 26326 42820 26332 42832
rect 25700 42792 26332 42820
rect 20622 42752 20628 42764
rect 20456 42724 20628 42752
rect 20456 42693 20484 42724
rect 20622 42712 20628 42724
rect 20680 42712 20686 42764
rect 20898 42712 20904 42764
rect 20956 42752 20962 42764
rect 21910 42752 21916 42764
rect 20956 42724 21916 42752
rect 20956 42712 20962 42724
rect 21910 42712 21916 42724
rect 21968 42752 21974 42764
rect 21968 42724 22508 42752
rect 21968 42712 21974 42724
rect 20441 42687 20499 42693
rect 20441 42653 20453 42687
rect 20487 42653 20499 42687
rect 20441 42647 20499 42653
rect 20533 42687 20591 42693
rect 20533 42653 20545 42687
rect 20579 42653 20591 42687
rect 20714 42684 20720 42696
rect 20675 42656 20720 42684
rect 20533 42647 20591 42653
rect 19797 42619 19855 42625
rect 19797 42585 19809 42619
rect 19843 42616 19855 42619
rect 20346 42616 20352 42628
rect 19843 42588 20352 42616
rect 19843 42585 19855 42588
rect 19797 42579 19855 42585
rect 20346 42576 20352 42588
rect 20404 42616 20410 42628
rect 20548 42616 20576 42647
rect 20714 42644 20720 42656
rect 20772 42644 20778 42696
rect 20809 42687 20867 42693
rect 20809 42653 20821 42687
rect 20855 42684 20867 42687
rect 21082 42684 21088 42696
rect 20855 42656 21088 42684
rect 20855 42653 20867 42656
rect 20809 42647 20867 42653
rect 21082 42644 21088 42656
rect 21140 42644 21146 42696
rect 21450 42684 21456 42696
rect 21411 42656 21456 42684
rect 21450 42644 21456 42656
rect 21508 42644 21514 42696
rect 21726 42684 21732 42696
rect 21687 42656 21732 42684
rect 21726 42644 21732 42656
rect 21784 42644 21790 42696
rect 22480 42693 22508 42724
rect 22646 42712 22652 42764
rect 22704 42752 22710 42764
rect 23198 42752 23204 42764
rect 22704 42724 23204 42752
rect 22704 42712 22710 42724
rect 23198 42712 23204 42724
rect 23256 42752 23262 42764
rect 23293 42755 23351 42761
rect 23293 42752 23305 42755
rect 23256 42724 23305 42752
rect 23256 42712 23262 42724
rect 23293 42721 23305 42724
rect 23339 42752 23351 42755
rect 23339 42724 24532 42752
rect 23339 42721 23351 42724
rect 23293 42715 23351 42721
rect 22189 42687 22247 42693
rect 22189 42653 22201 42687
rect 22235 42653 22247 42687
rect 22189 42647 22247 42653
rect 22465 42687 22523 42693
rect 22465 42653 22477 42687
rect 22511 42653 22523 42687
rect 22738 42684 22744 42696
rect 22465 42647 22523 42653
rect 22572 42656 22744 42684
rect 20990 42616 20996 42628
rect 20404 42588 20996 42616
rect 20404 42576 20410 42588
rect 20990 42576 20996 42588
rect 21048 42576 21054 42628
rect 21361 42619 21419 42625
rect 21361 42585 21373 42619
rect 21407 42616 21419 42619
rect 22204 42616 22232 42647
rect 22572 42616 22600 42656
rect 22738 42644 22744 42656
rect 22796 42644 22802 42696
rect 23382 42644 23388 42696
rect 23440 42684 23446 42696
rect 23658 42684 23664 42696
rect 23440 42656 23664 42684
rect 23440 42644 23446 42656
rect 23658 42644 23664 42656
rect 23716 42644 23722 42696
rect 23750 42644 23756 42696
rect 23808 42684 23814 42696
rect 24504 42684 24532 42724
rect 24670 42712 24676 42764
rect 24728 42752 24734 42764
rect 25700 42761 25728 42792
rect 26326 42780 26332 42792
rect 26384 42780 26390 42832
rect 26970 42780 26976 42832
rect 27028 42820 27034 42832
rect 28077 42823 28135 42829
rect 28077 42820 28089 42823
rect 27028 42792 28089 42820
rect 27028 42780 27034 42792
rect 28077 42789 28089 42792
rect 28123 42789 28135 42823
rect 29086 42820 29092 42832
rect 28077 42783 28135 42789
rect 28276 42792 29092 42820
rect 25501 42755 25559 42761
rect 25501 42752 25513 42755
rect 24728 42724 25513 42752
rect 24728 42712 24734 42724
rect 25501 42721 25513 42724
rect 25547 42721 25559 42755
rect 25501 42715 25559 42721
rect 25685 42755 25743 42761
rect 25685 42721 25697 42755
rect 25731 42721 25743 42755
rect 25685 42715 25743 42721
rect 25961 42755 26019 42761
rect 25961 42721 25973 42755
rect 26007 42752 26019 42755
rect 26418 42752 26424 42764
rect 26007 42724 26424 42752
rect 26007 42721 26019 42724
rect 25961 42715 26019 42721
rect 26418 42712 26424 42724
rect 26476 42712 26482 42764
rect 26786 42712 26792 42764
rect 26844 42752 26850 42764
rect 27157 42755 27215 42761
rect 27157 42752 27169 42755
rect 26844 42724 27169 42752
rect 26844 42712 26850 42724
rect 27157 42721 27169 42724
rect 27203 42721 27215 42755
rect 27157 42715 27215 42721
rect 27430 42712 27436 42764
rect 27488 42752 27494 42764
rect 28166 42752 28172 42764
rect 27488 42724 28172 42752
rect 27488 42712 27494 42724
rect 28166 42712 28172 42724
rect 28224 42712 28230 42764
rect 28276 42761 28304 42792
rect 29086 42780 29092 42792
rect 29144 42780 29150 42832
rect 31404 42820 31432 42851
rect 30116 42792 31432 42820
rect 28261 42755 28319 42761
rect 28261 42721 28273 42755
rect 28307 42721 28319 42755
rect 28261 42715 28319 42721
rect 28721 42755 28779 42761
rect 28721 42721 28733 42755
rect 28767 42752 28779 42755
rect 29454 42752 29460 42764
rect 28767 42724 29460 42752
rect 28767 42721 28779 42724
rect 28721 42715 28779 42721
rect 29454 42712 29460 42724
rect 29512 42712 29518 42764
rect 25038 42684 25044 42696
rect 23808 42656 24440 42684
rect 24504 42656 25044 42684
rect 23808 42644 23814 42656
rect 21407 42588 21680 42616
rect 22204 42588 22600 42616
rect 22649 42619 22707 42625
rect 21407 42585 21419 42588
rect 21361 42579 21419 42585
rect 21652 42560 21680 42588
rect 22649 42585 22661 42619
rect 22695 42616 22707 42619
rect 24118 42616 24124 42628
rect 22695 42588 24124 42616
rect 22695 42585 22707 42588
rect 22649 42579 22707 42585
rect 24118 42576 24124 42588
rect 24176 42576 24182 42628
rect 24412 42616 24440 42656
rect 25038 42644 25044 42656
rect 25096 42644 25102 42696
rect 25774 42684 25780 42696
rect 25735 42656 25780 42684
rect 25774 42644 25780 42656
rect 25832 42644 25838 42696
rect 25869 42687 25927 42693
rect 25869 42653 25881 42687
rect 25915 42684 25927 42687
rect 26050 42684 26056 42696
rect 25915 42656 26056 42684
rect 25915 42653 25927 42656
rect 25869 42647 25927 42653
rect 26050 42644 26056 42656
rect 26108 42644 26114 42696
rect 26436 42684 26464 42712
rect 27065 42687 27123 42693
rect 27065 42684 27077 42687
rect 26436 42656 27077 42684
rect 27065 42653 27077 42656
rect 27111 42653 27123 42687
rect 27246 42684 27252 42696
rect 27207 42656 27252 42684
rect 27065 42647 27123 42653
rect 27246 42644 27252 42656
rect 27304 42644 27310 42696
rect 27338 42644 27344 42696
rect 27396 42684 27402 42696
rect 27985 42687 28043 42693
rect 27396 42656 27441 42684
rect 27396 42644 27402 42656
rect 27985 42653 27997 42687
rect 28031 42653 28043 42687
rect 27985 42647 28043 42653
rect 28905 42687 28963 42693
rect 28905 42653 28917 42687
rect 28951 42684 28963 42687
rect 29270 42684 29276 42696
rect 28951 42656 29276 42684
rect 28951 42653 28963 42656
rect 28905 42647 28963 42653
rect 28000 42616 28028 42647
rect 29270 42644 29276 42656
rect 29328 42644 29334 42696
rect 29730 42644 29736 42696
rect 29788 42684 29794 42696
rect 29917 42687 29975 42693
rect 29917 42684 29929 42687
rect 29788 42656 29929 42684
rect 29788 42644 29794 42656
rect 29917 42653 29929 42656
rect 29963 42653 29975 42687
rect 29917 42647 29975 42653
rect 30006 42644 30012 42696
rect 30064 42684 30070 42696
rect 30116 42693 30144 42792
rect 31938 42780 31944 42832
rect 31996 42820 32002 42832
rect 31996 42792 32628 42820
rect 31996 42780 32002 42792
rect 32600 42764 32628 42792
rect 32950 42780 32956 42832
rect 33008 42820 33014 42832
rect 33689 42823 33747 42829
rect 33689 42820 33701 42823
rect 33008 42792 33701 42820
rect 33008 42780 33014 42792
rect 33689 42789 33701 42792
rect 33735 42789 33747 42823
rect 33689 42783 33747 42789
rect 31481 42755 31539 42761
rect 31481 42721 31493 42755
rect 31527 42752 31539 42755
rect 32398 42752 32404 42764
rect 31527 42724 32404 42752
rect 31527 42721 31539 42724
rect 31481 42715 31539 42721
rect 32398 42712 32404 42724
rect 32456 42712 32462 42764
rect 32582 42712 32588 42764
rect 32640 42752 32646 42764
rect 35802 42752 35808 42764
rect 32640 42724 35808 42752
rect 32640 42712 32646 42724
rect 30101 42687 30159 42693
rect 30101 42684 30113 42687
rect 30064 42656 30113 42684
rect 30064 42644 30070 42656
rect 30101 42653 30113 42656
rect 30147 42653 30159 42687
rect 30101 42647 30159 42653
rect 31573 42687 31631 42693
rect 31573 42653 31585 42687
rect 31619 42684 31631 42687
rect 31754 42684 31760 42696
rect 31619 42656 31760 42684
rect 31619 42653 31631 42656
rect 31573 42647 31631 42653
rect 31754 42644 31760 42656
rect 31812 42684 31818 42696
rect 33428 42693 33456 42724
rect 35802 42712 35808 42724
rect 35860 42712 35866 42764
rect 32493 42687 32551 42693
rect 32493 42684 32505 42687
rect 31812 42656 32505 42684
rect 31812 42644 31818 42656
rect 32493 42653 32505 42656
rect 32539 42653 32551 42687
rect 32493 42647 32551 42653
rect 32677 42687 32735 42693
rect 32677 42653 32689 42687
rect 32723 42653 32735 42687
rect 32677 42647 32735 42653
rect 33413 42687 33471 42693
rect 33413 42653 33425 42687
rect 33459 42653 33471 42687
rect 33413 42647 33471 42653
rect 24412 42588 28028 42616
rect 29089 42619 29147 42625
rect 29089 42585 29101 42619
rect 29135 42585 29147 42619
rect 29089 42579 29147 42585
rect 20254 42548 20260 42560
rect 20215 42520 20260 42548
rect 20254 42508 20260 42520
rect 20312 42508 20318 42560
rect 21634 42508 21640 42560
rect 21692 42548 21698 42560
rect 22186 42548 22192 42560
rect 21692 42520 22192 42548
rect 21692 42508 21698 42520
rect 22186 42508 22192 42520
rect 22244 42548 22250 42560
rect 22281 42551 22339 42557
rect 22281 42548 22293 42551
rect 22244 42520 22293 42548
rect 22244 42508 22250 42520
rect 22281 42517 22293 42520
rect 22327 42517 22339 42551
rect 22281 42511 22339 42517
rect 22830 42508 22836 42560
rect 22888 42548 22894 42560
rect 24029 42551 24087 42557
rect 24029 42548 24041 42551
rect 22888 42520 24041 42548
rect 22888 42508 22894 42520
rect 24029 42517 24041 42520
rect 24075 42548 24087 42551
rect 26142 42548 26148 42560
rect 24075 42520 26148 42548
rect 24075 42517 24087 42520
rect 24029 42511 24087 42517
rect 26142 42508 26148 42520
rect 26200 42548 26206 42560
rect 27154 42548 27160 42560
rect 26200 42520 27160 42548
rect 26200 42508 26206 42520
rect 27154 42508 27160 42520
rect 27212 42508 27218 42560
rect 27522 42548 27528 42560
rect 27483 42520 27528 42548
rect 27522 42508 27528 42520
rect 27580 42508 27586 42560
rect 28258 42548 28264 42560
rect 28219 42520 28264 42548
rect 28258 42508 28264 42520
rect 28316 42508 28322 42560
rect 28442 42508 28448 42560
rect 28500 42548 28506 42560
rect 29104 42548 29132 42579
rect 31846 42576 31852 42628
rect 31904 42616 31910 42628
rect 32692 42616 32720 42647
rect 33778 42644 33784 42696
rect 33836 42684 33842 42696
rect 34149 42687 34207 42693
rect 34149 42684 34161 42687
rect 33836 42656 34161 42684
rect 33836 42644 33842 42656
rect 34149 42653 34161 42656
rect 34195 42684 34207 42687
rect 34885 42687 34943 42693
rect 34885 42684 34897 42687
rect 34195 42656 34897 42684
rect 34195 42653 34207 42656
rect 34149 42647 34207 42653
rect 34885 42653 34897 42656
rect 34931 42653 34943 42687
rect 34885 42647 34943 42653
rect 33042 42616 33048 42628
rect 31904 42588 33048 42616
rect 31904 42576 31910 42588
rect 33042 42576 33048 42588
rect 33100 42576 33106 42628
rect 33502 42576 33508 42628
rect 33560 42616 33566 42628
rect 35069 42619 35127 42625
rect 35069 42616 35081 42619
rect 33560 42588 35081 42616
rect 33560 42576 33566 42588
rect 35069 42585 35081 42588
rect 35115 42585 35127 42619
rect 35069 42579 35127 42585
rect 29822 42548 29828 42560
rect 28500 42520 29828 42548
rect 28500 42508 28506 42520
rect 29822 42508 29828 42520
rect 29880 42508 29886 42560
rect 32585 42551 32643 42557
rect 32585 42517 32597 42551
rect 32631 42548 32643 42551
rect 33410 42548 33416 42560
rect 32631 42520 33416 42548
rect 32631 42517 32643 42520
rect 32585 42511 32643 42517
rect 33410 42508 33416 42520
rect 33468 42508 33474 42560
rect 33686 42508 33692 42560
rect 33744 42548 33750 42560
rect 35253 42551 35311 42557
rect 35253 42548 35265 42551
rect 33744 42520 35265 42548
rect 33744 42508 33750 42520
rect 35253 42517 35265 42520
rect 35299 42517 35311 42551
rect 35802 42548 35808 42560
rect 35715 42520 35808 42548
rect 35253 42511 35311 42517
rect 35802 42508 35808 42520
rect 35860 42548 35866 42560
rect 37090 42548 37096 42560
rect 35860 42520 37096 42548
rect 35860 42508 35866 42520
rect 37090 42508 37096 42520
rect 37148 42508 37154 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 20441 42347 20499 42353
rect 20441 42313 20453 42347
rect 20487 42344 20499 42347
rect 20622 42344 20628 42356
rect 20487 42316 20628 42344
rect 20487 42313 20499 42316
rect 20441 42307 20499 42313
rect 20622 42304 20628 42316
rect 20680 42304 20686 42356
rect 21726 42304 21732 42356
rect 21784 42344 21790 42356
rect 21784 42316 22508 42344
rect 21784 42304 21790 42316
rect 20162 42276 20168 42288
rect 19720 42248 20168 42276
rect 19720 42217 19748 42248
rect 20162 42236 20168 42248
rect 20220 42276 20226 42288
rect 20898 42276 20904 42288
rect 20220 42248 20484 42276
rect 20220 42236 20226 42248
rect 20456 42220 20484 42248
rect 20640 42248 20904 42276
rect 19705 42211 19763 42217
rect 19705 42177 19717 42211
rect 19751 42177 19763 42211
rect 19705 42171 19763 42177
rect 20349 42211 20407 42217
rect 20349 42177 20361 42211
rect 20395 42177 20407 42211
rect 20349 42171 20407 42177
rect 19613 42143 19671 42149
rect 19613 42109 19625 42143
rect 19659 42109 19671 42143
rect 19613 42103 19671 42109
rect 19797 42143 19855 42149
rect 19797 42109 19809 42143
rect 19843 42140 19855 42143
rect 20364 42140 20392 42171
rect 20438 42168 20444 42220
rect 20496 42168 20502 42220
rect 20640 42217 20668 42248
rect 20898 42236 20904 42248
rect 20956 42236 20962 42288
rect 21818 42236 21824 42288
rect 21876 42276 21882 42288
rect 22480 42276 22508 42316
rect 23658 42304 23664 42356
rect 23716 42344 23722 42356
rect 26050 42344 26056 42356
rect 23716 42316 26056 42344
rect 23716 42304 23722 42316
rect 26050 42304 26056 42316
rect 26108 42304 26114 42356
rect 27709 42347 27767 42353
rect 27709 42313 27721 42347
rect 27755 42344 27767 42347
rect 27982 42344 27988 42356
rect 27755 42316 27988 42344
rect 27755 42313 27767 42316
rect 27709 42307 27767 42313
rect 27982 42304 27988 42316
rect 28040 42344 28046 42356
rect 28810 42344 28816 42356
rect 28040 42316 28816 42344
rect 28040 42304 28046 42316
rect 28810 42304 28816 42316
rect 28868 42304 28874 42356
rect 29638 42344 29644 42356
rect 29048 42316 29644 42344
rect 23474 42276 23480 42288
rect 21876 42248 22413 42276
rect 21876 42236 21882 42248
rect 20625 42211 20683 42217
rect 20625 42177 20637 42211
rect 20671 42177 20683 42211
rect 20625 42171 20683 42177
rect 20714 42168 20720 42220
rect 20772 42208 20778 42220
rect 21361 42211 21419 42217
rect 21361 42208 21373 42211
rect 20772 42180 21373 42208
rect 20772 42168 20778 42180
rect 21361 42177 21373 42180
rect 21407 42177 21419 42211
rect 21361 42171 21419 42177
rect 22002 42168 22008 42220
rect 22060 42208 22066 42220
rect 22385 42217 22413 42248
rect 22480 42248 23480 42276
rect 22480 42217 22508 42248
rect 23474 42236 23480 42248
rect 23532 42236 23538 42288
rect 23842 42236 23848 42288
rect 23900 42276 23906 42288
rect 27798 42276 27804 42288
rect 23900 42248 24624 42276
rect 23900 42236 23906 42248
rect 22281 42211 22339 42217
rect 22281 42208 22293 42211
rect 22060 42180 22293 42208
rect 22060 42168 22066 42180
rect 22281 42177 22293 42180
rect 22327 42177 22339 42211
rect 22281 42171 22339 42177
rect 22373 42211 22431 42217
rect 22373 42177 22385 42211
rect 22419 42177 22431 42211
rect 22373 42171 22431 42177
rect 22465 42211 22523 42217
rect 22465 42177 22477 42211
rect 22511 42177 22523 42211
rect 22465 42171 22523 42177
rect 22649 42211 22707 42217
rect 22649 42177 22661 42211
rect 22695 42208 22707 42211
rect 22738 42208 22744 42220
rect 22695 42180 22744 42208
rect 22695 42177 22707 42180
rect 22649 42171 22707 42177
rect 22738 42168 22744 42180
rect 22796 42168 22802 42220
rect 23658 42208 23664 42220
rect 23619 42180 23664 42208
rect 23658 42168 23664 42180
rect 23716 42168 23722 42220
rect 24596 42217 24624 42248
rect 25148 42248 27804 42276
rect 24397 42211 24455 42217
rect 23768 42180 24348 42208
rect 23768 42149 23796 42180
rect 23385 42143 23443 42149
rect 23385 42140 23397 42143
rect 19843 42112 23397 42140
rect 19843 42109 19855 42112
rect 19797 42103 19855 42109
rect 23385 42109 23397 42112
rect 23431 42109 23443 42143
rect 23385 42103 23443 42109
rect 23569 42143 23627 42149
rect 23569 42109 23581 42143
rect 23615 42109 23627 42143
rect 23569 42103 23627 42109
rect 23753 42143 23811 42149
rect 23753 42109 23765 42143
rect 23799 42109 23811 42143
rect 23753 42103 23811 42109
rect 23845 42143 23903 42149
rect 23845 42109 23857 42143
rect 23891 42140 23903 42143
rect 24210 42140 24216 42152
rect 23891 42112 24216 42140
rect 23891 42109 23903 42112
rect 23845 42103 23903 42109
rect 19628 42072 19656 42103
rect 21910 42072 21916 42084
rect 19628 42044 21916 42072
rect 21910 42032 21916 42044
rect 21968 42072 21974 42084
rect 22005 42075 22063 42081
rect 22005 42072 22017 42075
rect 21968 42044 22017 42072
rect 21968 42032 21974 42044
rect 22005 42041 22017 42044
rect 22051 42041 22063 42075
rect 22005 42035 22063 42041
rect 22370 42032 22376 42084
rect 22428 42072 22434 42084
rect 23014 42072 23020 42084
rect 22428 42044 23020 42072
rect 22428 42032 22434 42044
rect 23014 42032 23020 42044
rect 23072 42032 23078 42084
rect 23585 42072 23613 42103
rect 24210 42100 24216 42112
rect 24268 42100 24274 42152
rect 23934 42072 23940 42084
rect 23585 42044 23940 42072
rect 23934 42032 23940 42044
rect 23992 42032 23998 42084
rect 24320 42072 24348 42180
rect 24397 42177 24409 42211
rect 24443 42177 24455 42211
rect 24397 42171 24455 42177
rect 24581 42211 24639 42217
rect 24581 42177 24593 42211
rect 24627 42208 24639 42211
rect 24670 42208 24676 42220
rect 24627 42180 24676 42208
rect 24627 42177 24639 42180
rect 24581 42171 24639 42177
rect 24412 42140 24440 42171
rect 24670 42168 24676 42180
rect 24728 42168 24734 42220
rect 25038 42208 25044 42220
rect 24951 42180 25044 42208
rect 25038 42168 25044 42180
rect 25096 42208 25102 42220
rect 25148 42208 25176 42248
rect 27798 42236 27804 42248
rect 27856 42236 27862 42288
rect 28626 42276 28632 42288
rect 28587 42248 28632 42276
rect 28626 42236 28632 42248
rect 28684 42236 28690 42288
rect 29048 42276 29076 42316
rect 29638 42304 29644 42316
rect 29696 42304 29702 42356
rect 31846 42344 31852 42356
rect 31680 42316 31852 42344
rect 30006 42276 30012 42288
rect 29012 42248 29076 42276
rect 29104 42248 30012 42276
rect 25096 42180 25176 42208
rect 25225 42211 25283 42217
rect 25096 42168 25102 42180
rect 25225 42177 25237 42211
rect 25271 42208 25283 42211
rect 25682 42208 25688 42220
rect 25271 42180 25688 42208
rect 25271 42177 25283 42180
rect 25225 42171 25283 42177
rect 25682 42168 25688 42180
rect 25740 42168 25746 42220
rect 25866 42208 25872 42220
rect 25827 42180 25872 42208
rect 25866 42168 25872 42180
rect 25924 42168 25930 42220
rect 26053 42211 26111 42217
rect 26053 42177 26065 42211
rect 26099 42208 26111 42211
rect 26234 42208 26240 42220
rect 26099 42180 26240 42208
rect 26099 42177 26111 42180
rect 26053 42171 26111 42177
rect 26234 42168 26240 42180
rect 26292 42168 26298 42220
rect 27706 42211 27764 42217
rect 27706 42177 27718 42211
rect 27752 42208 27764 42211
rect 28074 42208 28080 42220
rect 27752 42180 28080 42208
rect 27752 42177 27764 42180
rect 27706 42171 27764 42177
rect 28074 42168 28080 42180
rect 28132 42208 28138 42220
rect 28132 42198 28718 42208
rect 28132 42180 28764 42198
rect 28132 42168 28138 42180
rect 28690 42170 28764 42180
rect 26326 42140 26332 42152
rect 24412 42112 26332 42140
rect 25056 42084 25084 42112
rect 26326 42100 26332 42112
rect 26384 42140 26390 42152
rect 28169 42143 28227 42149
rect 28169 42140 28181 42143
rect 26384 42112 28181 42140
rect 26384 42100 26390 42112
rect 28169 42109 28181 42112
rect 28215 42109 28227 42143
rect 28736 42140 28764 42170
rect 28810 42168 28816 42220
rect 28868 42214 28874 42220
rect 29012 42217 29040 42248
rect 29104 42220 29132 42248
rect 30006 42236 30012 42248
rect 30064 42236 30070 42288
rect 30742 42236 30748 42288
rect 30800 42276 30806 42288
rect 31680 42276 31708 42316
rect 31846 42304 31852 42316
rect 31904 42304 31910 42356
rect 33134 42304 33140 42356
rect 33192 42344 33198 42356
rect 33192 42316 34376 42344
rect 33192 42304 33198 42316
rect 30800 42248 31708 42276
rect 30800 42236 30806 42248
rect 28905 42214 28963 42217
rect 28868 42211 28963 42214
rect 28868 42186 28917 42211
rect 28868 42168 28874 42186
rect 28905 42177 28917 42186
rect 28951 42177 28963 42211
rect 28905 42171 28963 42177
rect 28997 42211 29055 42217
rect 28997 42177 29009 42211
rect 29043 42177 29055 42211
rect 28997 42171 29055 42177
rect 29086 42168 29092 42220
rect 29144 42208 29150 42220
rect 29273 42211 29331 42217
rect 29144 42180 29237 42208
rect 29144 42168 29150 42180
rect 29273 42177 29285 42211
rect 29319 42208 29331 42211
rect 29454 42208 29460 42220
rect 29319 42180 29460 42208
rect 29319 42177 29331 42180
rect 29273 42171 29331 42177
rect 29454 42168 29460 42180
rect 29512 42168 29518 42220
rect 30282 42168 30288 42220
rect 30340 42208 30346 42220
rect 30377 42211 30435 42217
rect 30377 42208 30389 42211
rect 30340 42180 30389 42208
rect 30340 42168 30346 42180
rect 30377 42177 30389 42180
rect 30423 42177 30435 42211
rect 30377 42171 30435 42177
rect 30466 42168 30472 42220
rect 30524 42208 30530 42220
rect 30650 42208 30656 42220
rect 30524 42180 30569 42208
rect 30611 42180 30656 42208
rect 30524 42168 30530 42180
rect 30650 42168 30656 42180
rect 30708 42168 30714 42220
rect 31570 42217 31576 42220
rect 31389 42211 31447 42217
rect 31389 42177 31401 42211
rect 31435 42177 31447 42211
rect 31389 42171 31447 42177
rect 31554 42211 31576 42217
rect 31554 42177 31566 42211
rect 31554 42171 31576 42177
rect 31404 42140 31432 42171
rect 31570 42168 31576 42171
rect 31628 42168 31634 42220
rect 31680 42217 31708 42248
rect 32306 42236 32312 42288
rect 32364 42276 32370 42288
rect 32364 42248 32904 42276
rect 32364 42236 32370 42248
rect 31665 42211 31723 42217
rect 31665 42177 31677 42211
rect 31711 42177 31723 42211
rect 31665 42171 31723 42177
rect 31757 42211 31815 42217
rect 31938 42211 31944 42220
rect 31757 42177 31769 42211
rect 31803 42183 31944 42211
rect 31803 42177 31815 42183
rect 31757 42171 31815 42177
rect 31938 42168 31944 42183
rect 31996 42168 32002 42220
rect 32493 42211 32551 42217
rect 32493 42177 32505 42211
rect 32539 42177 32551 42211
rect 32493 42171 32551 42177
rect 32508 42140 32536 42171
rect 32674 42168 32680 42220
rect 32732 42208 32738 42220
rect 32769 42211 32827 42217
rect 32769 42208 32781 42211
rect 32732 42180 32781 42208
rect 32732 42168 32738 42180
rect 32769 42177 32781 42180
rect 32815 42177 32827 42211
rect 32769 42171 32827 42177
rect 28736 42112 32536 42140
rect 32876 42140 32904 42248
rect 33686 42236 33692 42288
rect 33744 42276 33750 42288
rect 33744 42248 34100 42276
rect 33744 42236 33750 42248
rect 33042 42168 33048 42220
rect 33100 42208 33106 42220
rect 34072 42217 34100 42248
rect 33873 42214 33931 42217
rect 33796 42211 33931 42214
rect 33796 42208 33885 42211
rect 33100 42186 33885 42208
rect 33100 42180 33824 42186
rect 33100 42168 33106 42180
rect 33873 42177 33885 42186
rect 33919 42177 33931 42211
rect 33873 42171 33931 42177
rect 33965 42211 34023 42217
rect 33965 42177 33977 42211
rect 34011 42177 34023 42211
rect 33965 42171 34023 42177
rect 34057 42211 34115 42217
rect 34057 42177 34069 42211
rect 34103 42177 34115 42211
rect 34057 42171 34115 42177
rect 34253 42211 34311 42217
rect 34253 42177 34265 42211
rect 34299 42208 34311 42211
rect 34348 42208 34376 42316
rect 34790 42208 34796 42220
rect 34299 42180 34796 42208
rect 34299 42177 34311 42180
rect 34253 42171 34311 42177
rect 33980 42140 34008 42171
rect 34790 42168 34796 42180
rect 34848 42168 34854 42220
rect 34698 42140 34704 42152
rect 32876 42112 34704 42140
rect 28169 42103 28227 42109
rect 34698 42100 34704 42112
rect 34756 42100 34762 42152
rect 24486 42072 24492 42084
rect 24320 42044 24492 42072
rect 24486 42032 24492 42044
rect 24544 42032 24550 42084
rect 25038 42032 25044 42084
rect 25096 42032 25102 42084
rect 26970 42072 26976 42084
rect 26068 42044 26976 42072
rect 19429 42007 19487 42013
rect 19429 41973 19441 42007
rect 19475 42004 19487 42007
rect 20070 42004 20076 42016
rect 19475 41976 20076 42004
rect 19475 41973 19487 41976
rect 19429 41967 19487 41973
rect 20070 41964 20076 41976
rect 20128 41964 20134 42016
rect 20809 42007 20867 42013
rect 20809 41973 20821 42007
rect 20855 42004 20867 42007
rect 21266 42004 21272 42016
rect 20855 41976 21272 42004
rect 20855 41973 20867 41976
rect 20809 41967 20867 41973
rect 21266 41964 21272 41976
rect 21324 41964 21330 42016
rect 21818 41964 21824 42016
rect 21876 42004 21882 42016
rect 24578 42004 24584 42016
rect 21876 41976 24584 42004
rect 21876 41964 21882 41976
rect 24578 41964 24584 41976
rect 24636 41964 24642 42016
rect 25133 42007 25191 42013
rect 25133 41973 25145 42007
rect 25179 42004 25191 42007
rect 25314 42004 25320 42016
rect 25179 41976 25320 42004
rect 25179 41973 25191 41976
rect 25133 41967 25191 41973
rect 25314 41964 25320 41976
rect 25372 41964 25378 42016
rect 25682 42004 25688 42016
rect 25643 41976 25688 42004
rect 25682 41964 25688 41976
rect 25740 41964 25746 42016
rect 26068 42013 26096 42044
rect 26970 42032 26976 42044
rect 27028 42032 27034 42084
rect 28077 42075 28135 42081
rect 28077 42041 28089 42075
rect 28123 42072 28135 42075
rect 29454 42072 29460 42084
rect 28123 42044 29460 42072
rect 28123 42041 28135 42044
rect 28077 42035 28135 42041
rect 29454 42032 29460 42044
rect 29512 42032 29518 42084
rect 30561 42075 30619 42081
rect 30561 42041 30573 42075
rect 30607 42072 30619 42075
rect 33597 42075 33655 42081
rect 33597 42072 33609 42075
rect 30607 42044 31340 42072
rect 30607 42041 30619 42044
rect 30561 42035 30619 42041
rect 26053 42007 26111 42013
rect 26053 41973 26065 42007
rect 26099 41973 26111 42007
rect 26602 42004 26608 42016
rect 26563 41976 26608 42004
rect 26053 41967 26111 41973
rect 26602 41964 26608 41976
rect 26660 41964 26666 42016
rect 26878 41964 26884 42016
rect 26936 42004 26942 42016
rect 27525 42007 27583 42013
rect 27525 42004 27537 42007
rect 26936 41976 27537 42004
rect 26936 41964 26942 41976
rect 27525 41973 27537 41976
rect 27571 41973 27583 42007
rect 27525 41967 27583 41973
rect 27982 41964 27988 42016
rect 28040 42004 28046 42016
rect 30193 42007 30251 42013
rect 30193 42004 30205 42007
rect 28040 41976 30205 42004
rect 28040 41964 28046 41976
rect 30193 41973 30205 41976
rect 30239 41973 30251 42007
rect 30193 41967 30251 41973
rect 30742 41964 30748 42016
rect 30800 42004 30806 42016
rect 31205 42007 31263 42013
rect 31205 42004 31217 42007
rect 30800 41976 31217 42004
rect 30800 41964 30806 41976
rect 31205 41973 31217 41976
rect 31251 41973 31263 42007
rect 31312 42004 31340 42044
rect 31496 42044 33609 42072
rect 31496 42004 31524 42044
rect 33597 42041 33609 42044
rect 33643 42041 33655 42075
rect 33597 42035 33655 42041
rect 31312 41976 31524 42004
rect 31205 41967 31263 41973
rect 32030 41964 32036 42016
rect 32088 42004 32094 42016
rect 32309 42007 32367 42013
rect 32309 42004 32321 42007
rect 32088 41976 32321 42004
rect 32088 41964 32094 41976
rect 32309 41973 32321 41976
rect 32355 41973 32367 42007
rect 32309 41967 32367 41973
rect 32582 41964 32588 42016
rect 32640 42004 32646 42016
rect 32677 42007 32735 42013
rect 32677 42004 32689 42007
rect 32640 41976 32689 42004
rect 32640 41964 32646 41976
rect 32677 41973 32689 41976
rect 32723 41973 32735 42007
rect 32677 41967 32735 41973
rect 33962 41964 33968 42016
rect 34020 42004 34026 42016
rect 34793 42007 34851 42013
rect 34793 42004 34805 42007
rect 34020 41976 34805 42004
rect 34020 41964 34026 41976
rect 34793 41973 34805 41976
rect 34839 41973 34851 42007
rect 34793 41967 34851 41973
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 21450 41760 21456 41812
rect 21508 41800 21514 41812
rect 23658 41800 23664 41812
rect 21508 41772 22416 41800
rect 23619 41772 23664 41800
rect 21508 41760 21514 41772
rect 21542 41692 21548 41744
rect 21600 41732 21606 41744
rect 21821 41735 21879 41741
rect 21821 41732 21833 41735
rect 21600 41704 21833 41732
rect 21600 41692 21606 41704
rect 21821 41701 21833 41704
rect 21867 41732 21879 41735
rect 22186 41732 22192 41744
rect 21867 41704 22192 41732
rect 21867 41701 21879 41704
rect 21821 41695 21879 41701
rect 22186 41692 22192 41704
rect 22244 41692 22250 41744
rect 20073 41667 20131 41673
rect 20073 41633 20085 41667
rect 20119 41664 20131 41667
rect 20346 41664 20352 41676
rect 20119 41636 20352 41664
rect 20119 41633 20131 41636
rect 20073 41627 20131 41633
rect 20346 41624 20352 41636
rect 20404 41664 20410 41676
rect 20404 41636 21680 41664
rect 20404 41624 20410 41636
rect 21652 41537 21680 41636
rect 21910 41556 21916 41608
rect 21968 41596 21974 41608
rect 22388 41605 22416 41772
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 23750 41760 23756 41812
rect 23808 41800 23814 41812
rect 23845 41803 23903 41809
rect 23845 41800 23857 41803
rect 23808 41772 23857 41800
rect 23808 41760 23814 41772
rect 23845 41769 23857 41772
rect 23891 41769 23903 41803
rect 23845 41763 23903 41769
rect 26789 41803 26847 41809
rect 26789 41769 26801 41803
rect 26835 41800 26847 41803
rect 26970 41800 26976 41812
rect 26835 41772 26976 41800
rect 26835 41769 26847 41772
rect 26789 41763 26847 41769
rect 26970 41760 26976 41772
rect 27028 41760 27034 41812
rect 30650 41800 30656 41812
rect 27080 41772 28994 41800
rect 30611 41772 30656 41800
rect 24673 41735 24731 41741
rect 24673 41732 24685 41735
rect 23584 41704 24685 41732
rect 23584 41664 23612 41704
rect 24673 41701 24685 41704
rect 24719 41732 24731 41735
rect 27080 41732 27108 41772
rect 24719 41704 27108 41732
rect 28966 41732 28994 41772
rect 30650 41760 30656 41772
rect 30708 41760 30714 41812
rect 31202 41760 31208 41812
rect 31260 41800 31266 41812
rect 33594 41800 33600 41812
rect 31260 41772 33600 41800
rect 31260 41760 31266 41772
rect 33594 41760 33600 41772
rect 33652 41760 33658 41812
rect 34698 41760 34704 41812
rect 34756 41800 34762 41812
rect 34977 41803 35035 41809
rect 34977 41800 34989 41803
rect 34756 41772 34989 41800
rect 34756 41760 34762 41772
rect 34977 41769 34989 41772
rect 35023 41769 35035 41803
rect 34977 41763 35035 41769
rect 31294 41732 31300 41744
rect 28966 41704 31300 41732
rect 24719 41701 24731 41704
rect 24673 41695 24731 41701
rect 31294 41692 31300 41704
rect 31352 41732 31358 41744
rect 31938 41732 31944 41744
rect 31352 41704 31944 41732
rect 31352 41692 31358 41704
rect 31938 41692 31944 41704
rect 31996 41692 32002 41744
rect 32493 41735 32551 41741
rect 32493 41701 32505 41735
rect 32539 41732 32551 41735
rect 32582 41732 32588 41744
rect 32539 41704 32588 41732
rect 32539 41701 32551 41704
rect 32493 41695 32551 41701
rect 32582 41692 32588 41704
rect 32640 41692 32646 41744
rect 35342 41732 35348 41744
rect 32692 41704 35348 41732
rect 22572 41636 23612 41664
rect 22373 41599 22431 41605
rect 21968 41568 22013 41596
rect 21968 41556 21974 41568
rect 22373 41565 22385 41599
rect 22419 41596 22431 41599
rect 22462 41596 22468 41608
rect 22419 41568 22468 41596
rect 22419 41565 22431 41568
rect 22373 41559 22431 41565
rect 22462 41556 22468 41568
rect 22520 41556 22526 41608
rect 21637 41531 21695 41537
rect 21637 41497 21649 41531
rect 21683 41528 21695 41531
rect 22572 41528 22600 41636
rect 24578 41624 24584 41676
rect 24636 41664 24642 41676
rect 27890 41664 27896 41676
rect 24636 41636 25452 41664
rect 24636 41624 24642 41636
rect 25038 41596 25044 41608
rect 23492 41568 25044 41596
rect 21683 41500 22600 41528
rect 21683 41497 21695 41500
rect 21637 41491 21695 41497
rect 22738 41488 22744 41540
rect 22796 41488 22802 41540
rect 23492 41537 23520 41568
rect 25038 41556 25044 41568
rect 25096 41556 25102 41608
rect 25314 41596 25320 41608
rect 25275 41568 25320 41596
rect 25314 41556 25320 41568
rect 25372 41556 25378 41608
rect 25424 41605 25452 41636
rect 27172 41636 27896 41664
rect 25409 41599 25467 41605
rect 25409 41565 25421 41599
rect 25455 41565 25467 41599
rect 25590 41596 25596 41608
rect 25551 41568 25596 41596
rect 25409 41559 25467 41565
rect 25590 41556 25596 41568
rect 25648 41556 25654 41608
rect 25685 41599 25743 41605
rect 25685 41565 25697 41599
rect 25731 41596 25743 41599
rect 25866 41596 25872 41608
rect 25731 41568 25872 41596
rect 25731 41565 25743 41568
rect 25685 41559 25743 41565
rect 25866 41556 25872 41568
rect 25924 41596 25930 41608
rect 27062 41596 27068 41608
rect 25924 41568 26372 41596
rect 27023 41568 27068 41596
rect 25924 41556 25930 41568
rect 23477 41531 23535 41537
rect 23477 41497 23489 41531
rect 23523 41497 23535 41531
rect 23477 41491 23535 41497
rect 23693 41531 23751 41537
rect 23693 41497 23705 41531
rect 23739 41528 23751 41531
rect 24302 41528 24308 41540
rect 23739 41500 24308 41528
rect 23739 41497 23751 41500
rect 23693 41491 23751 41497
rect 20438 41420 20444 41472
rect 20496 41460 20502 41472
rect 20533 41463 20591 41469
rect 20533 41460 20545 41463
rect 20496 41432 20545 41460
rect 20496 41420 20502 41432
rect 20533 41429 20545 41432
rect 20579 41429 20591 41463
rect 20533 41423 20591 41429
rect 20898 41420 20904 41472
rect 20956 41460 20962 41472
rect 21085 41463 21143 41469
rect 21085 41460 21097 41463
rect 20956 41432 21097 41460
rect 20956 41420 20962 41432
rect 21085 41429 21097 41432
rect 21131 41429 21143 41463
rect 21910 41460 21916 41472
rect 21871 41432 21916 41460
rect 21085 41423 21143 41429
rect 21910 41420 21916 41432
rect 21968 41420 21974 41472
rect 22557 41463 22615 41469
rect 22557 41429 22569 41463
rect 22603 41460 22615 41463
rect 22756 41460 22784 41488
rect 23492 41460 23520 41491
rect 24302 41488 24308 41500
rect 24360 41528 24366 41540
rect 26142 41528 26148 41540
rect 24360 41500 26148 41528
rect 24360 41488 24366 41500
rect 26142 41488 26148 41500
rect 26200 41488 26206 41540
rect 26344 41528 26372 41568
rect 27062 41556 27068 41568
rect 27120 41556 27126 41608
rect 27172 41605 27200 41636
rect 27890 41624 27896 41636
rect 27948 41624 27954 41676
rect 29270 41664 29276 41676
rect 28828 41636 29276 41664
rect 27157 41599 27215 41605
rect 27157 41565 27169 41599
rect 27203 41565 27215 41599
rect 27157 41559 27215 41565
rect 27249 41599 27307 41605
rect 27249 41565 27261 41599
rect 27295 41596 27307 41599
rect 27338 41596 27344 41608
rect 27295 41568 27344 41596
rect 27295 41565 27307 41568
rect 27249 41559 27307 41565
rect 27338 41556 27344 41568
rect 27396 41556 27402 41608
rect 27430 41556 27436 41608
rect 27488 41596 27494 41608
rect 27488 41568 27533 41596
rect 27488 41556 27494 41568
rect 27614 41556 27620 41608
rect 27672 41596 27678 41608
rect 28537 41599 28595 41605
rect 28537 41596 28549 41599
rect 27672 41568 28549 41596
rect 27672 41556 27678 41568
rect 28537 41565 28549 41568
rect 28583 41565 28595 41599
rect 28537 41559 28595 41565
rect 28629 41599 28687 41605
rect 28629 41565 28641 41599
rect 28675 41565 28687 41599
rect 28629 41559 28687 41565
rect 28644 41528 28672 41559
rect 28828 41540 28856 41636
rect 29270 41624 29276 41636
rect 29328 41624 29334 41676
rect 28997 41599 29055 41605
rect 28997 41565 29009 41599
rect 29043 41596 29055 41599
rect 29546 41596 29552 41608
rect 29043 41568 29552 41596
rect 29043 41565 29055 41568
rect 28997 41559 29055 41565
rect 29546 41556 29552 41568
rect 29604 41556 29610 41608
rect 29730 41596 29736 41608
rect 29691 41568 29736 41596
rect 29730 41556 29736 41568
rect 29788 41556 29794 41608
rect 29914 41596 29920 41608
rect 29875 41568 29920 41596
rect 29914 41556 29920 41568
rect 29972 41556 29978 41608
rect 30742 41596 30748 41608
rect 30703 41568 30748 41596
rect 30742 41556 30748 41568
rect 30800 41556 30806 41608
rect 30837 41599 30895 41605
rect 30837 41565 30849 41599
rect 30883 41596 30895 41599
rect 30926 41596 30932 41608
rect 30883 41568 30932 41596
rect 30883 41565 30895 41568
rect 30837 41559 30895 41565
rect 30926 41556 30932 41568
rect 30984 41556 30990 41608
rect 31386 41556 31392 41608
rect 31444 41596 31450 41608
rect 31570 41596 31576 41608
rect 31444 41568 31576 41596
rect 31444 41556 31450 41568
rect 31570 41556 31576 41568
rect 31628 41556 31634 41608
rect 32692 41605 32720 41704
rect 35342 41692 35348 41704
rect 35400 41692 35406 41744
rect 33042 41624 33048 41676
rect 33100 41664 33106 41676
rect 35161 41667 35219 41673
rect 35161 41664 35173 41667
rect 33100 41636 35173 41664
rect 33100 41624 33106 41636
rect 35161 41633 35173 41636
rect 35207 41633 35219 41667
rect 35161 41627 35219 41633
rect 32677 41599 32735 41605
rect 32677 41565 32689 41599
rect 32723 41565 32735 41599
rect 32677 41559 32735 41565
rect 32953 41599 33011 41605
rect 32953 41565 32965 41599
rect 32999 41565 33011 41599
rect 33594 41596 33600 41608
rect 33555 41568 33600 41596
rect 32953 41559 33011 41565
rect 28810 41528 28816 41540
rect 26344 41500 28672 41528
rect 28771 41500 28816 41528
rect 28810 41488 28816 41500
rect 28868 41488 28874 41540
rect 28905 41531 28963 41537
rect 28905 41497 28917 41531
rect 28951 41497 28963 41531
rect 30561 41531 30619 41537
rect 30561 41528 30573 41531
rect 28905 41491 28963 41497
rect 29196 41500 30573 41528
rect 25130 41460 25136 41472
rect 22603 41432 23520 41460
rect 25091 41432 25136 41460
rect 22603 41429 22615 41432
rect 22557 41423 22615 41429
rect 25130 41420 25136 41432
rect 25188 41420 25194 41472
rect 26329 41463 26387 41469
rect 26329 41429 26341 41463
rect 26375 41460 26387 41463
rect 26510 41460 26516 41472
rect 26375 41432 26516 41460
rect 26375 41429 26387 41432
rect 26329 41423 26387 41429
rect 26510 41420 26516 41432
rect 26568 41420 26574 41472
rect 26602 41420 26608 41472
rect 26660 41460 26666 41472
rect 27893 41463 27951 41469
rect 27893 41460 27905 41463
rect 26660 41432 27905 41460
rect 26660 41420 26666 41432
rect 27893 41429 27905 41432
rect 27939 41460 27951 41463
rect 28074 41460 28080 41472
rect 27939 41432 28080 41460
rect 27939 41429 27951 41432
rect 27893 41423 27951 41429
rect 28074 41420 28080 41432
rect 28132 41420 28138 41472
rect 28718 41420 28724 41472
rect 28776 41460 28782 41472
rect 28920 41460 28948 41491
rect 29196 41469 29224 41500
rect 30561 41497 30573 41500
rect 30607 41497 30619 41531
rect 32968 41528 32996 41559
rect 33594 41556 33600 41568
rect 33652 41556 33658 41608
rect 34790 41556 34796 41608
rect 34848 41596 34854 41608
rect 34885 41599 34943 41605
rect 34885 41596 34897 41599
rect 34848 41568 34897 41596
rect 34848 41556 34854 41568
rect 34885 41565 34897 41568
rect 34931 41565 34943 41599
rect 34885 41559 34943 41565
rect 35621 41599 35679 41605
rect 35621 41565 35633 41599
rect 35667 41596 35679 41599
rect 35894 41596 35900 41608
rect 35667 41568 35900 41596
rect 35667 41565 35679 41568
rect 35621 41559 35679 41565
rect 35894 41556 35900 41568
rect 35952 41596 35958 41608
rect 35952 41568 36400 41596
rect 35952 41556 35958 41568
rect 33413 41531 33471 41537
rect 33413 41528 33425 41531
rect 32968 41500 33425 41528
rect 30561 41491 30619 41497
rect 33413 41497 33425 41500
rect 33459 41497 33471 41531
rect 33778 41528 33784 41540
rect 33739 41500 33784 41528
rect 33413 41491 33471 41497
rect 28776 41432 28948 41460
rect 29181 41463 29239 41469
rect 28776 41420 28782 41432
rect 29181 41429 29193 41463
rect 29227 41429 29239 41463
rect 29181 41423 29239 41429
rect 29825 41463 29883 41469
rect 29825 41429 29837 41463
rect 29871 41460 29883 41463
rect 30006 41460 30012 41472
rect 29871 41432 30012 41460
rect 29871 41429 29883 41432
rect 29825 41423 29883 41429
rect 30006 41420 30012 41432
rect 30064 41420 30070 41472
rect 32766 41420 32772 41472
rect 32824 41460 32830 41472
rect 32861 41463 32919 41469
rect 32861 41460 32873 41463
rect 32824 41432 32873 41460
rect 32824 41420 32830 41432
rect 32861 41429 32873 41432
rect 32907 41429 32919 41463
rect 33428 41460 33456 41491
rect 33778 41488 33784 41500
rect 33836 41488 33842 41540
rect 33686 41460 33692 41472
rect 33428 41432 33692 41460
rect 32861 41423 32919 41429
rect 33686 41420 33692 41432
rect 33744 41420 33750 41472
rect 35158 41460 35164 41472
rect 35119 41432 35164 41460
rect 35158 41420 35164 41432
rect 35216 41420 35222 41472
rect 35710 41460 35716 41472
rect 35671 41432 35716 41460
rect 35710 41420 35716 41432
rect 35768 41420 35774 41472
rect 36372 41469 36400 41568
rect 36357 41463 36415 41469
rect 36357 41429 36369 41463
rect 36403 41460 36415 41463
rect 37458 41460 37464 41472
rect 36403 41432 37464 41460
rect 36403 41429 36415 41432
rect 36357 41423 36415 41429
rect 37458 41420 37464 41432
rect 37516 41420 37522 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 21174 41216 21180 41268
rect 21232 41256 21238 41268
rect 23017 41259 23075 41265
rect 23017 41256 23029 41259
rect 21232 41228 23029 41256
rect 21232 41216 21238 41228
rect 23017 41225 23029 41228
rect 23063 41225 23075 41259
rect 23017 41219 23075 41225
rect 23185 41259 23243 41265
rect 23185 41225 23197 41259
rect 23231 41256 23243 41259
rect 24762 41256 24768 41268
rect 23231 41228 24768 41256
rect 23231 41225 23243 41228
rect 23185 41219 23243 41225
rect 24762 41216 24768 41228
rect 24820 41216 24826 41268
rect 25590 41216 25596 41268
rect 25648 41256 25654 41268
rect 26234 41256 26240 41268
rect 25648 41228 26240 41256
rect 25648 41216 25654 41228
rect 26234 41216 26240 41228
rect 26292 41216 26298 41268
rect 26970 41216 26976 41268
rect 27028 41256 27034 41268
rect 27028 41228 27568 41256
rect 27028 41216 27034 41228
rect 20622 41188 20628 41200
rect 19904 41160 20628 41188
rect 19334 41080 19340 41132
rect 19392 41120 19398 41132
rect 19904 41120 19932 41160
rect 20622 41148 20628 41160
rect 20680 41148 20686 41200
rect 23382 41188 23388 41200
rect 23343 41160 23388 41188
rect 23382 41148 23388 41160
rect 23440 41148 23446 41200
rect 24486 41148 24492 41200
rect 24544 41188 24550 41200
rect 24544 41160 25452 41188
rect 24544 41148 24550 41160
rect 20070 41120 20076 41132
rect 19392 41092 19932 41120
rect 20031 41092 20076 41120
rect 19392 41080 19398 41092
rect 20070 41080 20076 41092
rect 20128 41080 20134 41132
rect 20165 41123 20223 41129
rect 20165 41089 20177 41123
rect 20211 41120 20223 41123
rect 20901 41123 20959 41129
rect 20901 41120 20913 41123
rect 20211 41092 20913 41120
rect 20211 41089 20223 41092
rect 20165 41083 20223 41089
rect 20901 41089 20913 41092
rect 20947 41089 20959 41123
rect 21082 41120 21088 41132
rect 21043 41092 21088 41120
rect 20901 41083 20959 41089
rect 21082 41080 21088 41092
rect 21140 41080 21146 41132
rect 21361 41123 21419 41129
rect 21361 41089 21373 41123
rect 21407 41120 21419 41123
rect 21450 41120 21456 41132
rect 21407 41092 21456 41120
rect 21407 41089 21419 41092
rect 21361 41083 21419 41089
rect 21450 41080 21456 41092
rect 21508 41080 21514 41132
rect 22186 41120 22192 41132
rect 22147 41092 22192 41120
rect 22186 41080 22192 41092
rect 22244 41080 22250 41132
rect 22462 41120 22468 41132
rect 22423 41092 22468 41120
rect 22462 41080 22468 41092
rect 22520 41080 22526 41132
rect 23290 41080 23296 41132
rect 23348 41120 23354 41132
rect 24029 41123 24087 41129
rect 24029 41120 24041 41123
rect 23348 41092 24041 41120
rect 23348 41080 23354 41092
rect 24029 41089 24041 41092
rect 24075 41089 24087 41123
rect 24029 41083 24087 41089
rect 24213 41123 24271 41129
rect 24213 41089 24225 41123
rect 24259 41120 24271 41123
rect 24854 41120 24860 41132
rect 24259 41092 24860 41120
rect 24259 41089 24271 41092
rect 24213 41083 24271 41089
rect 24854 41080 24860 41092
rect 24912 41080 24918 41132
rect 24949 41123 25007 41129
rect 24949 41089 24961 41123
rect 24995 41089 25007 41123
rect 25130 41120 25136 41132
rect 25091 41092 25136 41120
rect 24949 41083 25007 41089
rect 20441 41055 20499 41061
rect 20441 41052 20453 41055
rect 18708 41024 20453 41052
rect 18708 40928 18736 41024
rect 20441 41021 20453 41024
rect 20487 41052 20499 41055
rect 20714 41052 20720 41064
rect 20487 41024 20720 41052
rect 20487 41021 20499 41024
rect 20441 41015 20499 41021
rect 20714 41012 20720 41024
rect 20772 41012 20778 41064
rect 21177 41055 21235 41061
rect 21177 41021 21189 41055
rect 21223 41052 21235 41055
rect 21818 41052 21824 41064
rect 21223 41024 21824 41052
rect 21223 41021 21235 41024
rect 21177 41015 21235 41021
rect 21818 41012 21824 41024
rect 21876 41012 21882 41064
rect 22373 41055 22431 41061
rect 22373 41021 22385 41055
rect 22419 41021 22431 41055
rect 22373 41015 22431 41021
rect 20349 40987 20407 40993
rect 20349 40953 20361 40987
rect 20395 40984 20407 40987
rect 21269 40987 21327 40993
rect 20395 40956 21128 40984
rect 20395 40953 20407 40956
rect 20349 40947 20407 40953
rect 18690 40916 18696 40928
rect 18651 40888 18696 40916
rect 18690 40876 18696 40888
rect 18748 40876 18754 40928
rect 19889 40919 19947 40925
rect 19889 40885 19901 40919
rect 19935 40916 19947 40919
rect 20622 40916 20628 40928
rect 19935 40888 20628 40916
rect 19935 40885 19947 40888
rect 19889 40879 19947 40885
rect 20622 40876 20628 40888
rect 20680 40876 20686 40928
rect 21100 40916 21128 40956
rect 21269 40953 21281 40987
rect 21315 40984 21327 40987
rect 21358 40984 21364 40996
rect 21315 40956 21364 40984
rect 21315 40953 21327 40956
rect 21269 40947 21327 40953
rect 21358 40944 21364 40956
rect 21416 40944 21422 40996
rect 21542 40944 21548 40996
rect 21600 40984 21606 40996
rect 22281 40987 22339 40993
rect 22281 40984 22293 40987
rect 21600 40956 22293 40984
rect 21600 40944 21606 40956
rect 22281 40953 22293 40956
rect 22327 40953 22339 40987
rect 22281 40947 22339 40953
rect 22005 40919 22063 40925
rect 22005 40916 22017 40919
rect 21100 40888 22017 40916
rect 22005 40885 22017 40888
rect 22051 40885 22063 40919
rect 22388 40916 22416 41015
rect 22922 41012 22928 41064
rect 22980 41052 22986 41064
rect 23106 41052 23112 41064
rect 22980 41024 23112 41052
rect 22980 41012 22986 41024
rect 23106 41012 23112 41024
rect 23164 41012 23170 41064
rect 23934 41012 23940 41064
rect 23992 41052 23998 41064
rect 24121 41055 24179 41061
rect 24121 41052 24133 41055
rect 23992 41024 24133 41052
rect 23992 41012 23998 41024
rect 24121 41021 24133 41024
rect 24167 41021 24179 41055
rect 24121 41015 24179 41021
rect 24302 41012 24308 41064
rect 24360 41052 24366 41064
rect 24489 41055 24547 41061
rect 24360 41024 24405 41052
rect 24360 41012 24366 41024
rect 24489 41021 24501 41055
rect 24535 41052 24547 41055
rect 24964 41052 24992 41083
rect 25130 41080 25136 41092
rect 25188 41080 25194 41132
rect 25424 41129 25452 41160
rect 26142 41148 26148 41200
rect 26200 41188 26206 41200
rect 26389 41191 26447 41197
rect 26389 41188 26401 41191
rect 26200 41160 26401 41188
rect 26200 41148 26206 41160
rect 26389 41157 26401 41160
rect 26435 41188 26447 41191
rect 26435 41157 26448 41188
rect 26389 41151 26448 41157
rect 25409 41123 25467 41129
rect 25409 41089 25421 41123
rect 25455 41089 25467 41123
rect 25682 41120 25688 41132
rect 25643 41092 25688 41120
rect 25409 41083 25467 41089
rect 25682 41080 25688 41092
rect 25740 41080 25746 41132
rect 26420 41120 26448 41151
rect 26510 41148 26516 41200
rect 26568 41188 26574 41200
rect 26605 41191 26663 41197
rect 26605 41188 26617 41191
rect 26568 41160 26617 41188
rect 26568 41148 26574 41160
rect 26605 41157 26617 41160
rect 26651 41188 26663 41191
rect 27338 41188 27344 41200
rect 26651 41160 27344 41188
rect 26651 41157 26663 41160
rect 26605 41151 26663 41157
rect 27338 41148 27344 41160
rect 27396 41148 27402 41200
rect 27540 41188 27568 41228
rect 27798 41216 27804 41268
rect 27856 41256 27862 41268
rect 28810 41256 28816 41268
rect 27856 41228 28816 41256
rect 27856 41216 27862 41228
rect 28810 41216 28816 41228
rect 28868 41216 28874 41268
rect 31018 41256 31024 41268
rect 28966 41228 31024 41256
rect 28966 41188 28994 41228
rect 31018 41216 31024 41228
rect 31076 41216 31082 41268
rect 31478 41256 31484 41268
rect 31391 41228 31484 41256
rect 31478 41216 31484 41228
rect 31536 41256 31542 41268
rect 31754 41256 31760 41268
rect 31536 41228 31760 41256
rect 31536 41216 31542 41228
rect 31754 41216 31760 41228
rect 31812 41216 31818 41268
rect 32122 41216 32128 41268
rect 32180 41256 32186 41268
rect 32509 41259 32567 41265
rect 32509 41256 32521 41259
rect 32180 41228 32521 41256
rect 32180 41216 32186 41228
rect 32509 41225 32521 41228
rect 32555 41225 32567 41259
rect 32509 41219 32567 41225
rect 33778 41216 33784 41268
rect 33836 41216 33842 41268
rect 29549 41191 29607 41197
rect 27540 41160 28994 41188
rect 29196 41160 29500 41188
rect 27540 41129 27568 41160
rect 27433 41123 27491 41129
rect 27433 41120 27445 41123
rect 26420 41092 27445 41120
rect 27433 41089 27445 41092
rect 27479 41089 27491 41123
rect 27433 41083 27491 41089
rect 27525 41123 27583 41129
rect 27525 41089 27537 41123
rect 27571 41089 27583 41123
rect 27525 41083 27583 41089
rect 27614 41080 27620 41132
rect 27672 41120 27678 41132
rect 29196 41120 29224 41160
rect 27672 41092 29224 41120
rect 27672 41080 27678 41092
rect 29270 41080 29276 41132
rect 29328 41120 29334 41132
rect 29365 41123 29423 41129
rect 29365 41120 29377 41123
rect 29328 41092 29377 41120
rect 29328 41080 29334 41092
rect 29365 41089 29377 41092
rect 29411 41089 29423 41123
rect 29472 41120 29500 41160
rect 29549 41157 29561 41191
rect 29595 41188 29607 41191
rect 29914 41188 29920 41200
rect 29595 41160 29920 41188
rect 29595 41157 29607 41160
rect 29549 41151 29607 41157
rect 29914 41148 29920 41160
rect 29972 41148 29978 41200
rect 32309 41191 32367 41197
rect 32309 41157 32321 41191
rect 32355 41188 32367 41191
rect 32674 41188 32680 41200
rect 32355 41160 32680 41188
rect 32355 41157 32367 41160
rect 32309 41151 32367 41157
rect 32674 41148 32680 41160
rect 32732 41148 32738 41200
rect 33594 41188 33600 41200
rect 32876 41160 33600 41188
rect 29733 41123 29791 41129
rect 29733 41120 29745 41123
rect 29472 41092 29745 41120
rect 29365 41083 29423 41089
rect 29733 41089 29745 41092
rect 29779 41120 29791 41123
rect 30098 41120 30104 41132
rect 29779 41092 30104 41120
rect 29779 41089 29791 41092
rect 29733 41083 29791 41089
rect 30098 41080 30104 41092
rect 30156 41120 30162 41132
rect 30193 41123 30251 41129
rect 30193 41120 30205 41123
rect 30156 41092 30205 41120
rect 30156 41080 30162 41092
rect 30193 41089 30205 41092
rect 30239 41089 30251 41123
rect 30193 41083 30251 41089
rect 32214 41080 32220 41132
rect 32272 41120 32278 41132
rect 32876 41120 32904 41160
rect 33594 41148 33600 41160
rect 33652 41188 33658 41200
rect 33796 41188 33824 41216
rect 33652 41160 33824 41188
rect 33652 41148 33658 41160
rect 32272 41092 32904 41120
rect 32272 41080 32278 41092
rect 33134 41080 33140 41132
rect 33192 41120 33198 41132
rect 33505 41123 33563 41129
rect 33505 41120 33517 41123
rect 33192 41092 33517 41120
rect 33192 41080 33198 41092
rect 33505 41089 33517 41092
rect 33551 41089 33563 41123
rect 33686 41120 33692 41132
rect 33647 41092 33692 41120
rect 33505 41083 33563 41089
rect 33686 41080 33692 41092
rect 33744 41080 33750 41132
rect 33781 41123 33839 41129
rect 33781 41089 33793 41123
rect 33827 41089 33839 41123
rect 33962 41120 33968 41132
rect 33923 41092 33968 41120
rect 33781 41083 33839 41089
rect 24535 41024 24992 41052
rect 24535 41021 24547 41024
rect 24489 41015 24547 41021
rect 27154 41012 27160 41064
rect 27212 41052 27218 41064
rect 27249 41055 27307 41061
rect 27249 41052 27261 41055
rect 27212 41024 27261 41052
rect 27212 41012 27218 41024
rect 27249 41021 27261 41024
rect 27295 41021 27307 41055
rect 27249 41015 27307 41021
rect 27338 41012 27344 41064
rect 27396 41052 27402 41064
rect 32582 41052 32588 41064
rect 27396 41024 32588 41052
rect 27396 41012 27402 41024
rect 32582 41012 32588 41024
rect 32640 41012 32646 41064
rect 33796 41052 33824 41083
rect 33962 41080 33968 41092
rect 34020 41120 34026 41132
rect 34425 41123 34483 41129
rect 34425 41120 34437 41123
rect 34020 41092 34437 41120
rect 34020 41080 34026 41092
rect 34425 41089 34437 41092
rect 34471 41089 34483 41123
rect 34425 41083 34483 41089
rect 35158 41052 35164 41064
rect 32692 41024 33732 41052
rect 33796 41024 35164 41052
rect 25314 40984 25320 40996
rect 25275 40956 25320 40984
rect 25314 40944 25320 40956
rect 25372 40944 25378 40996
rect 28074 40984 28080 40996
rect 26436 40956 28080 40984
rect 26436 40928 26464 40956
rect 28074 40944 28080 40956
rect 28132 40944 28138 40996
rect 29914 40944 29920 40996
rect 29972 40984 29978 40996
rect 30745 40987 30803 40993
rect 30745 40984 30757 40987
rect 29972 40956 30757 40984
rect 29972 40944 29978 40956
rect 30745 40953 30757 40956
rect 30791 40984 30803 40987
rect 30926 40984 30932 40996
rect 30791 40956 30932 40984
rect 30791 40953 30803 40956
rect 30745 40947 30803 40953
rect 30926 40944 30932 40956
rect 30984 40984 30990 40996
rect 32122 40984 32128 40996
rect 30984 40956 32128 40984
rect 30984 40944 30990 40956
rect 32122 40944 32128 40956
rect 32180 40984 32186 40996
rect 32692 40984 32720 41024
rect 32180 40956 32720 40984
rect 32180 40944 32186 40956
rect 33042 40944 33048 40996
rect 33100 40984 33106 40996
rect 33597 40987 33655 40993
rect 33597 40984 33609 40987
rect 33100 40956 33609 40984
rect 33100 40944 33106 40956
rect 33597 40953 33609 40956
rect 33643 40953 33655 40987
rect 33704 40984 33732 41024
rect 35158 41012 35164 41024
rect 35216 41012 35222 41064
rect 33778 40984 33784 40996
rect 33704 40956 33784 40984
rect 33597 40947 33655 40953
rect 33778 40944 33784 40956
rect 33836 40944 33842 40996
rect 22922 40916 22928 40928
rect 22388 40888 22928 40916
rect 22005 40879 22063 40885
rect 22922 40876 22928 40888
rect 22980 40876 22986 40928
rect 23201 40919 23259 40925
rect 23201 40885 23213 40919
rect 23247 40916 23259 40919
rect 23474 40916 23480 40928
rect 23247 40888 23480 40916
rect 23247 40885 23259 40888
rect 23201 40879 23259 40885
rect 23474 40876 23480 40888
rect 23532 40876 23538 40928
rect 26418 40916 26424 40928
rect 26379 40888 26424 40916
rect 26418 40876 26424 40888
rect 26476 40876 26482 40928
rect 27062 40876 27068 40928
rect 27120 40916 27126 40928
rect 27341 40919 27399 40925
rect 27341 40916 27353 40919
rect 27120 40888 27353 40916
rect 27120 40876 27126 40888
rect 27341 40885 27353 40888
rect 27387 40885 27399 40919
rect 27341 40879 27399 40885
rect 27798 40876 27804 40928
rect 27856 40916 27862 40928
rect 28261 40919 28319 40925
rect 28261 40916 28273 40919
rect 27856 40888 28273 40916
rect 27856 40876 27862 40888
rect 28261 40885 28273 40888
rect 28307 40885 28319 40919
rect 28261 40879 28319 40885
rect 28810 40876 28816 40928
rect 28868 40916 28874 40928
rect 28905 40919 28963 40925
rect 28905 40916 28917 40919
rect 28868 40888 28917 40916
rect 28868 40876 28874 40888
rect 28905 40885 28917 40888
rect 28951 40916 28963 40919
rect 30282 40916 30288 40928
rect 28951 40888 30288 40916
rect 28951 40885 28963 40888
rect 28905 40879 28963 40885
rect 30282 40876 30288 40888
rect 30340 40876 30346 40928
rect 30374 40876 30380 40928
rect 30432 40916 30438 40928
rect 32306 40916 32312 40928
rect 30432 40888 32312 40916
rect 30432 40876 30438 40888
rect 32306 40876 32312 40888
rect 32364 40916 32370 40928
rect 32493 40919 32551 40925
rect 32493 40916 32505 40919
rect 32364 40888 32505 40916
rect 32364 40876 32370 40888
rect 32493 40885 32505 40888
rect 32539 40885 32551 40919
rect 32674 40916 32680 40928
rect 32635 40888 32680 40916
rect 32493 40879 32551 40885
rect 32674 40876 32680 40888
rect 32732 40876 32738 40928
rect 33226 40876 33232 40928
rect 33284 40916 33290 40928
rect 33321 40919 33379 40925
rect 33321 40916 33333 40919
rect 33284 40888 33333 40916
rect 33284 40876 33290 40888
rect 33321 40885 33333 40888
rect 33367 40885 33379 40919
rect 33321 40879 33379 40885
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 20165 40715 20223 40721
rect 20165 40681 20177 40715
rect 20211 40712 20223 40715
rect 20254 40712 20260 40724
rect 20211 40684 20260 40712
rect 20211 40681 20223 40684
rect 20165 40675 20223 40681
rect 20254 40672 20260 40684
rect 20312 40672 20318 40724
rect 21634 40672 21640 40724
rect 21692 40712 21698 40724
rect 23934 40712 23940 40724
rect 21692 40684 23940 40712
rect 21692 40672 21698 40684
rect 23934 40672 23940 40684
rect 23992 40672 23998 40724
rect 24302 40672 24308 40724
rect 24360 40712 24366 40724
rect 24673 40715 24731 40721
rect 24673 40712 24685 40715
rect 24360 40684 24685 40712
rect 24360 40672 24366 40684
rect 24673 40681 24685 40684
rect 24719 40681 24731 40715
rect 24673 40675 24731 40681
rect 26234 40672 26240 40724
rect 26292 40712 26298 40724
rect 26602 40712 26608 40724
rect 26292 40684 26608 40712
rect 26292 40672 26298 40684
rect 26602 40672 26608 40684
rect 26660 40672 26666 40724
rect 27246 40672 27252 40724
rect 27304 40672 27310 40724
rect 28166 40672 28172 40724
rect 28224 40712 28230 40724
rect 28537 40715 28595 40721
rect 28537 40712 28549 40715
rect 28224 40684 28549 40712
rect 28224 40672 28230 40684
rect 28537 40681 28549 40684
rect 28583 40681 28595 40715
rect 28537 40675 28595 40681
rect 31938 40672 31944 40724
rect 31996 40712 32002 40724
rect 32306 40712 32312 40724
rect 31996 40684 32312 40712
rect 31996 40672 32002 40684
rect 32306 40672 32312 40684
rect 32364 40712 32370 40724
rect 33873 40715 33931 40721
rect 33873 40712 33885 40715
rect 32364 40684 33885 40712
rect 32364 40672 32370 40684
rect 33873 40681 33885 40684
rect 33919 40681 33931 40715
rect 33873 40675 33931 40681
rect 23952 40644 23980 40672
rect 25225 40647 25283 40653
rect 25225 40644 25237 40647
rect 23952 40616 25237 40644
rect 25225 40613 25237 40616
rect 25271 40644 25283 40647
rect 25682 40644 25688 40656
rect 25271 40616 25688 40644
rect 25271 40613 25283 40616
rect 25225 40607 25283 40613
rect 25682 40604 25688 40616
rect 25740 40644 25746 40656
rect 25869 40647 25927 40653
rect 25869 40644 25881 40647
rect 25740 40616 25881 40644
rect 25740 40604 25746 40616
rect 25869 40613 25881 40616
rect 25915 40613 25927 40647
rect 25869 40607 25927 40613
rect 26510 40604 26516 40656
rect 26568 40644 26574 40656
rect 27264 40644 27292 40672
rect 30558 40644 30564 40656
rect 26568 40616 27200 40644
rect 27264 40616 30564 40644
rect 26568 40604 26574 40616
rect 18509 40579 18567 40585
rect 18509 40545 18521 40579
rect 18555 40576 18567 40579
rect 19426 40576 19432 40588
rect 18555 40548 19432 40576
rect 18555 40545 18567 40548
rect 18509 40539 18567 40545
rect 19426 40536 19432 40548
rect 19484 40536 19490 40588
rect 20257 40579 20315 40585
rect 20257 40545 20269 40579
rect 20303 40576 20315 40579
rect 21174 40576 21180 40588
rect 20303 40548 21180 40576
rect 20303 40545 20315 40548
rect 20257 40539 20315 40545
rect 21174 40536 21180 40548
rect 21232 40536 21238 40588
rect 23845 40579 23903 40585
rect 23845 40576 23857 40579
rect 22020 40548 23857 40576
rect 1857 40511 1915 40517
rect 1857 40477 1869 40511
rect 1903 40508 1915 40511
rect 1946 40508 1952 40520
rect 1903 40480 1952 40508
rect 1903 40477 1915 40480
rect 1857 40471 1915 40477
rect 1946 40468 1952 40480
rect 2004 40508 2010 40520
rect 2317 40511 2375 40517
rect 2317 40508 2329 40511
rect 2004 40480 2329 40508
rect 2004 40468 2010 40480
rect 2317 40477 2329 40480
rect 2363 40477 2375 40511
rect 2317 40471 2375 40477
rect 18233 40511 18291 40517
rect 18233 40477 18245 40511
rect 18279 40477 18291 40511
rect 18233 40471 18291 40477
rect 17773 40443 17831 40449
rect 17773 40409 17785 40443
rect 17819 40440 17831 40443
rect 18248 40440 18276 40471
rect 18322 40468 18328 40520
rect 18380 40508 18386 40520
rect 19795 40511 19853 40517
rect 18380 40480 18425 40508
rect 18380 40468 18386 40480
rect 19795 40477 19807 40511
rect 19841 40508 19853 40511
rect 21726 40508 21732 40520
rect 19841 40480 20208 40508
rect 21687 40480 21732 40508
rect 19841 40477 19853 40480
rect 19795 40471 19853 40477
rect 18874 40440 18880 40452
rect 17819 40412 18880 40440
rect 17819 40409 17831 40412
rect 17773 40403 17831 40409
rect 18874 40400 18880 40412
rect 18932 40400 18938 40452
rect 20180 40440 20208 40480
rect 21726 40468 21732 40480
rect 21784 40468 21790 40520
rect 22020 40517 22048 40548
rect 21821 40511 21879 40517
rect 21821 40477 21833 40511
rect 21867 40477 21879 40511
rect 21821 40471 21879 40477
rect 22005 40511 22063 40517
rect 22005 40477 22017 40511
rect 22051 40477 22063 40511
rect 22005 40471 22063 40477
rect 22097 40511 22155 40517
rect 22097 40477 22109 40511
rect 22143 40508 22155 40511
rect 22278 40508 22284 40520
rect 22143 40480 22284 40508
rect 22143 40477 22155 40480
rect 22097 40471 22155 40477
rect 21545 40443 21603 40449
rect 21545 40440 21557 40443
rect 20180 40412 21557 40440
rect 21545 40409 21557 40412
rect 21591 40409 21603 40443
rect 21836 40440 21864 40471
rect 22278 40468 22284 40480
rect 22336 40468 22342 40520
rect 22922 40508 22928 40520
rect 22883 40480 22928 40508
rect 22922 40468 22928 40480
rect 22980 40468 22986 40520
rect 23308 40517 23336 40548
rect 23845 40545 23857 40548
rect 23891 40545 23903 40579
rect 27062 40576 27068 40588
rect 27023 40548 27068 40576
rect 23845 40539 23903 40545
rect 27062 40536 27068 40548
rect 27120 40536 27126 40588
rect 27172 40576 27200 40616
rect 30558 40604 30564 40616
rect 30616 40604 30622 40656
rect 33686 40644 33692 40656
rect 30668 40616 33692 40644
rect 27249 40579 27307 40585
rect 27249 40576 27261 40579
rect 27172 40548 27261 40576
rect 27249 40545 27261 40548
rect 27295 40545 27307 40579
rect 27249 40539 27307 40545
rect 27338 40536 27344 40588
rect 27396 40576 27402 40588
rect 30668 40576 30696 40616
rect 33686 40604 33692 40616
rect 33744 40604 33750 40656
rect 27396 40548 27441 40576
rect 27540 40548 30696 40576
rect 27396 40536 27402 40548
rect 23017 40511 23075 40517
rect 23017 40477 23029 40511
rect 23063 40477 23075 40511
rect 23017 40471 23075 40477
rect 23201 40511 23259 40517
rect 23201 40477 23213 40511
rect 23247 40477 23259 40511
rect 23201 40471 23259 40477
rect 23293 40511 23351 40517
rect 23293 40477 23305 40511
rect 23339 40477 23351 40511
rect 23293 40471 23351 40477
rect 22830 40440 22836 40452
rect 21836 40412 22836 40440
rect 21545 40403 21603 40409
rect 22830 40400 22836 40412
rect 22888 40440 22894 40452
rect 23032 40440 23060 40471
rect 22888 40412 23060 40440
rect 23216 40440 23244 40471
rect 23658 40468 23664 40520
rect 23716 40508 23722 40520
rect 23753 40511 23811 40517
rect 23753 40508 23765 40511
rect 23716 40480 23765 40508
rect 23716 40468 23722 40480
rect 23753 40477 23765 40480
rect 23799 40477 23811 40511
rect 23753 40471 23811 40477
rect 23937 40511 23995 40517
rect 23937 40477 23949 40511
rect 23983 40508 23995 40511
rect 24026 40508 24032 40520
rect 23983 40480 24032 40508
rect 23983 40477 23995 40480
rect 23937 40471 23995 40477
rect 24026 40468 24032 40480
rect 24084 40508 24090 40520
rect 24210 40508 24216 40520
rect 24084 40480 24216 40508
rect 24084 40468 24090 40480
rect 24210 40468 24216 40480
rect 24268 40468 24274 40520
rect 24581 40511 24639 40517
rect 24581 40477 24593 40511
rect 24627 40477 24639 40511
rect 24762 40508 24768 40520
rect 24723 40480 24768 40508
rect 24581 40471 24639 40477
rect 23216 40412 23336 40440
rect 22888 40400 22894 40412
rect 1670 40372 1676 40384
rect 1631 40344 1676 40372
rect 1670 40332 1676 40344
rect 1728 40332 1734 40384
rect 18506 40372 18512 40384
rect 18467 40344 18512 40372
rect 18506 40332 18512 40344
rect 18564 40332 18570 40384
rect 18782 40332 18788 40384
rect 18840 40372 18846 40384
rect 19613 40375 19671 40381
rect 19613 40372 19625 40375
rect 18840 40344 19625 40372
rect 18840 40332 18846 40344
rect 19613 40341 19625 40344
rect 19659 40341 19671 40375
rect 19613 40335 19671 40341
rect 19797 40375 19855 40381
rect 19797 40341 19809 40375
rect 19843 40372 19855 40375
rect 19978 40372 19984 40384
rect 19843 40344 19984 40372
rect 19843 40341 19855 40344
rect 19797 40335 19855 40341
rect 19978 40332 19984 40344
rect 20036 40332 20042 40384
rect 21082 40372 21088 40384
rect 21043 40344 21088 40372
rect 21082 40332 21088 40344
rect 21140 40332 21146 40384
rect 21174 40332 21180 40384
rect 21232 40372 21238 40384
rect 21726 40372 21732 40384
rect 21232 40344 21732 40372
rect 21232 40332 21238 40344
rect 21726 40332 21732 40344
rect 21784 40332 21790 40384
rect 22741 40375 22799 40381
rect 22741 40341 22753 40375
rect 22787 40372 22799 40375
rect 23014 40372 23020 40384
rect 22787 40344 23020 40372
rect 22787 40341 22799 40344
rect 22741 40335 22799 40341
rect 23014 40332 23020 40344
rect 23072 40332 23078 40384
rect 23308 40372 23336 40412
rect 23382 40400 23388 40452
rect 23440 40440 23446 40452
rect 24596 40440 24624 40471
rect 24762 40468 24768 40480
rect 24820 40468 24826 40520
rect 27154 40508 27160 40520
rect 27115 40480 27160 40508
rect 27154 40468 27160 40480
rect 27212 40468 27218 40520
rect 25774 40440 25780 40452
rect 23440 40412 24624 40440
rect 24688 40412 25780 40440
rect 23440 40400 23446 40412
rect 24578 40372 24584 40384
rect 23308 40344 24584 40372
rect 24578 40332 24584 40344
rect 24636 40372 24642 40384
rect 24688 40372 24716 40412
rect 25774 40400 25780 40412
rect 25832 40400 25838 40452
rect 25958 40400 25964 40452
rect 26016 40440 26022 40452
rect 27540 40440 27568 40548
rect 27706 40468 27712 40520
rect 27764 40508 27770 40520
rect 28169 40511 28227 40517
rect 28169 40508 28181 40511
rect 27764 40480 28181 40508
rect 27764 40468 27770 40480
rect 28169 40477 28181 40480
rect 28215 40508 28227 40511
rect 28215 40480 28672 40508
rect 28215 40477 28227 40480
rect 28169 40471 28227 40477
rect 28534 40440 28540 40452
rect 26016 40412 27568 40440
rect 28495 40412 28540 40440
rect 26016 40400 26022 40412
rect 28534 40400 28540 40412
rect 28592 40400 28598 40452
rect 28644 40440 28672 40480
rect 28718 40468 28724 40520
rect 28776 40508 28782 40520
rect 29733 40511 29791 40517
rect 29733 40508 29745 40511
rect 28776 40480 29745 40508
rect 28776 40468 28782 40480
rect 29733 40477 29745 40480
rect 29779 40508 29791 40511
rect 29914 40508 29920 40520
rect 29779 40480 29920 40508
rect 29779 40477 29791 40480
rect 29733 40471 29791 40477
rect 29914 40468 29920 40480
rect 29972 40468 29978 40520
rect 30668 40517 30696 40548
rect 30929 40579 30987 40585
rect 30929 40545 30941 40579
rect 30975 40576 30987 40579
rect 31018 40576 31024 40588
rect 30975 40548 31024 40576
rect 30975 40545 30987 40548
rect 30929 40539 30987 40545
rect 31018 40536 31024 40548
rect 31076 40536 31082 40588
rect 31938 40576 31944 40588
rect 31772 40548 31944 40576
rect 31772 40517 31800 40548
rect 31938 40536 31944 40548
rect 31996 40536 32002 40588
rect 32600 40548 33272 40576
rect 30653 40511 30711 40517
rect 30653 40477 30665 40511
rect 30699 40477 30711 40511
rect 30653 40471 30711 40477
rect 31749 40511 31807 40517
rect 31749 40477 31761 40511
rect 31795 40477 31807 40511
rect 31749 40471 31807 40477
rect 31849 40511 31907 40517
rect 31849 40477 31861 40511
rect 31895 40477 31907 40511
rect 32030 40508 32036 40520
rect 31991 40480 32036 40508
rect 31849 40471 31907 40477
rect 31864 40440 31892 40471
rect 32030 40468 32036 40480
rect 32088 40468 32094 40520
rect 32125 40511 32183 40517
rect 32125 40477 32137 40511
rect 32171 40508 32183 40511
rect 32398 40508 32404 40520
rect 32171 40480 32404 40508
rect 32171 40477 32183 40480
rect 32125 40471 32183 40477
rect 32398 40468 32404 40480
rect 32456 40468 32462 40520
rect 32490 40468 32496 40520
rect 32548 40508 32554 40520
rect 32600 40517 32628 40548
rect 33244 40517 33272 40548
rect 32585 40511 32643 40517
rect 32585 40508 32597 40511
rect 32548 40480 32597 40508
rect 32548 40468 32554 40480
rect 32585 40477 32597 40480
rect 32631 40477 32643 40511
rect 32585 40471 32643 40477
rect 32769 40511 32827 40517
rect 32769 40477 32781 40511
rect 32815 40477 32827 40511
rect 32769 40471 32827 40477
rect 33229 40511 33287 40517
rect 33229 40477 33241 40511
rect 33275 40477 33287 40511
rect 33410 40508 33416 40520
rect 33371 40480 33416 40508
rect 33229 40471 33287 40477
rect 32677 40443 32735 40449
rect 32677 40440 32689 40443
rect 28644 40412 32689 40440
rect 32677 40409 32689 40412
rect 32723 40409 32735 40443
rect 32677 40403 32735 40409
rect 24636 40344 24716 40372
rect 24636 40332 24642 40344
rect 25498 40332 25504 40384
rect 25556 40372 25562 40384
rect 26421 40375 26479 40381
rect 26421 40372 26433 40375
rect 25556 40344 26433 40372
rect 25556 40332 25562 40344
rect 26421 40341 26433 40344
rect 26467 40372 26479 40375
rect 27154 40372 27160 40384
rect 26467 40344 27160 40372
rect 26467 40341 26479 40344
rect 26421 40335 26479 40341
rect 27154 40332 27160 40344
rect 27212 40332 27218 40384
rect 27430 40332 27436 40384
rect 27488 40372 27494 40384
rect 27525 40375 27583 40381
rect 27525 40372 27537 40375
rect 27488 40344 27537 40372
rect 27488 40332 27494 40344
rect 27525 40341 27537 40344
rect 27571 40341 27583 40375
rect 27525 40335 27583 40341
rect 28721 40375 28779 40381
rect 28721 40341 28733 40375
rect 28767 40372 28779 40375
rect 29178 40372 29184 40384
rect 28767 40344 29184 40372
rect 28767 40341 28779 40344
rect 28721 40335 28779 40341
rect 29178 40332 29184 40344
rect 29236 40332 29242 40384
rect 30282 40372 30288 40384
rect 30243 40344 30288 40372
rect 30282 40332 30288 40344
rect 30340 40332 30346 40384
rect 30558 40332 30564 40384
rect 30616 40372 30622 40384
rect 30745 40375 30803 40381
rect 30745 40372 30757 40375
rect 30616 40344 30757 40372
rect 30616 40332 30622 40344
rect 30745 40341 30757 40344
rect 30791 40341 30803 40375
rect 30745 40335 30803 40341
rect 31294 40332 31300 40384
rect 31352 40372 31358 40384
rect 31573 40375 31631 40381
rect 31573 40372 31585 40375
rect 31352 40344 31585 40372
rect 31352 40332 31358 40344
rect 31573 40341 31585 40344
rect 31619 40341 31631 40375
rect 31573 40335 31631 40341
rect 32490 40332 32496 40384
rect 32548 40372 32554 40384
rect 32784 40372 32812 40471
rect 33410 40468 33416 40480
rect 33468 40508 33474 40520
rect 33873 40511 33931 40517
rect 33873 40508 33885 40511
rect 33468 40480 33885 40508
rect 33468 40468 33474 40480
rect 33873 40477 33885 40480
rect 33919 40477 33931 40511
rect 33873 40471 33931 40477
rect 34057 40511 34115 40517
rect 34057 40477 34069 40511
rect 34103 40508 34115 40511
rect 35342 40508 35348 40520
rect 34103 40480 35348 40508
rect 34103 40477 34115 40480
rect 34057 40471 34115 40477
rect 35342 40468 35348 40480
rect 35400 40468 35406 40520
rect 58069 40511 58127 40517
rect 58069 40508 58081 40511
rect 57716 40480 58081 40508
rect 57716 40384 57744 40480
rect 58069 40477 58081 40480
rect 58115 40477 58127 40511
rect 58069 40471 58127 40477
rect 33318 40372 33324 40384
rect 32548 40344 32812 40372
rect 33279 40344 33324 40372
rect 32548 40332 32554 40344
rect 33318 40332 33324 40344
rect 33376 40332 33382 40384
rect 34977 40375 35035 40381
rect 34977 40341 34989 40375
rect 35023 40372 35035 40375
rect 35621 40375 35679 40381
rect 35621 40372 35633 40375
rect 35023 40344 35633 40372
rect 35023 40341 35035 40344
rect 34977 40335 35035 40341
rect 35621 40341 35633 40344
rect 35667 40372 35679 40375
rect 35802 40372 35808 40384
rect 35667 40344 35808 40372
rect 35667 40341 35679 40344
rect 35621 40335 35679 40341
rect 35802 40332 35808 40344
rect 35860 40332 35866 40384
rect 35894 40332 35900 40384
rect 35952 40372 35958 40384
rect 36081 40375 36139 40381
rect 36081 40372 36093 40375
rect 35952 40344 36093 40372
rect 35952 40332 35958 40344
rect 36081 40341 36093 40344
rect 36127 40341 36139 40375
rect 36081 40335 36139 40341
rect 57609 40375 57667 40381
rect 57609 40341 57621 40375
rect 57655 40372 57667 40375
rect 57698 40372 57704 40384
rect 57655 40344 57704 40372
rect 57655 40341 57667 40344
rect 57609 40335 57667 40341
rect 57698 40332 57704 40344
rect 57756 40332 57762 40384
rect 58250 40372 58256 40384
rect 58211 40344 58256 40372
rect 58250 40332 58256 40344
rect 58308 40332 58314 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 19886 40177 19892 40180
rect 19882 40168 19892 40177
rect 19847 40140 19892 40168
rect 19882 40131 19892 40140
rect 19886 40128 19892 40131
rect 19944 40128 19950 40180
rect 22094 40168 22100 40180
rect 19996 40140 22100 40168
rect 19996 40109 20024 40140
rect 22094 40128 22100 40140
rect 22152 40168 22158 40180
rect 22649 40171 22707 40177
rect 22152 40140 22600 40168
rect 22152 40128 22158 40140
rect 17313 40103 17371 40109
rect 17313 40069 17325 40103
rect 17359 40100 17371 40103
rect 19797 40103 19855 40109
rect 17359 40072 18644 40100
rect 17359 40069 17371 40072
rect 17313 40063 17371 40069
rect 17770 40032 17776 40044
rect 17731 40004 17776 40032
rect 17770 39992 17776 40004
rect 17828 39992 17834 40044
rect 17954 40032 17960 40044
rect 17915 40004 17960 40032
rect 17954 39992 17960 40004
rect 18012 39992 18018 40044
rect 18322 39992 18328 40044
rect 18380 40032 18386 40044
rect 18616 40041 18644 40072
rect 19797 40069 19809 40103
rect 19843 40100 19855 40103
rect 19981 40103 20039 40109
rect 19843 40072 19932 40100
rect 19843 40069 19855 40072
rect 19797 40063 19855 40069
rect 18417 40035 18475 40041
rect 18417 40032 18429 40035
rect 18380 40004 18429 40032
rect 18380 39992 18386 40004
rect 18417 40001 18429 40004
rect 18463 40001 18475 40035
rect 18417 39995 18475 40001
rect 18601 40035 18659 40041
rect 18601 40001 18613 40035
rect 18647 40032 18659 40035
rect 18874 40032 18880 40044
rect 18647 40004 18880 40032
rect 18647 40001 18659 40004
rect 18601 39995 18659 40001
rect 18874 39992 18880 40004
rect 18932 39992 18938 40044
rect 19334 39992 19340 40044
rect 19392 40032 19398 40044
rect 19705 40035 19763 40041
rect 19705 40032 19717 40035
rect 19392 40004 19717 40032
rect 19392 39992 19398 40004
rect 19705 40001 19717 40004
rect 19751 40001 19763 40035
rect 19904 40032 19932 40072
rect 19981 40069 19993 40103
rect 20027 40069 20039 40103
rect 20162 40100 20168 40112
rect 19981 40063 20039 40069
rect 20088 40072 20168 40100
rect 20088 40032 20116 40072
rect 20162 40060 20168 40072
rect 20220 40100 20226 40112
rect 20220 40072 22094 40100
rect 20220 40060 20226 40072
rect 22066 40044 22094 40072
rect 20898 40032 20904 40044
rect 19904 40004 20116 40032
rect 20859 40004 20904 40032
rect 19705 39995 19763 40001
rect 20898 39992 20904 40004
rect 20956 39992 20962 40044
rect 22066 40004 22100 40044
rect 22094 39992 22100 40004
rect 22152 39992 22158 40044
rect 22189 40035 22247 40041
rect 22189 40001 22201 40035
rect 22235 40032 22247 40035
rect 22278 40032 22284 40044
rect 22235 40004 22284 40032
rect 22235 40001 22247 40004
rect 22189 39995 22247 40001
rect 22278 39992 22284 40004
rect 22336 39992 22342 40044
rect 22572 40032 22600 40140
rect 22649 40137 22661 40171
rect 22695 40137 22707 40171
rect 22649 40131 22707 40137
rect 23293 40171 23351 40177
rect 23293 40137 23305 40171
rect 23339 40168 23351 40171
rect 23339 40140 27292 40168
rect 23339 40137 23351 40140
rect 23293 40131 23351 40137
rect 22664 40100 22692 40131
rect 23382 40100 23388 40112
rect 22664 40072 23388 40100
rect 23382 40060 23388 40072
rect 23440 40060 23446 40112
rect 27154 40100 27160 40112
rect 23998 40072 27160 40100
rect 22922 40032 22928 40044
rect 22572 40004 22928 40032
rect 22922 39992 22928 40004
rect 22980 39992 22986 40044
rect 23474 40032 23480 40044
rect 23387 40004 23480 40032
rect 23474 39992 23480 40004
rect 23532 40032 23538 40044
rect 23998 40032 24026 40072
rect 27154 40060 27160 40072
rect 27212 40060 27218 40112
rect 27264 40100 27292 40140
rect 27338 40128 27344 40180
rect 27396 40168 27402 40180
rect 29993 40171 30051 40177
rect 27396 40140 29316 40168
rect 27396 40128 27402 40140
rect 27614 40100 27620 40112
rect 27264 40072 27620 40100
rect 27614 40060 27620 40072
rect 27672 40060 27678 40112
rect 27982 40060 27988 40112
rect 28040 40100 28046 40112
rect 28534 40100 28540 40112
rect 28040 40072 28540 40100
rect 28040 40060 28046 40072
rect 28534 40060 28540 40072
rect 28592 40060 28598 40112
rect 28718 40100 28724 40112
rect 28690 40060 28724 40100
rect 28776 40060 28782 40112
rect 28905 40103 28963 40109
rect 28905 40069 28917 40103
rect 28951 40069 28963 40103
rect 29288 40100 29316 40140
rect 29993 40137 30005 40171
rect 30039 40168 30051 40171
rect 30282 40168 30288 40180
rect 30039 40140 30288 40168
rect 30039 40137 30051 40140
rect 29993 40131 30051 40137
rect 30282 40128 30288 40140
rect 30340 40128 30346 40180
rect 32214 40168 32220 40180
rect 30392 40140 32220 40168
rect 30193 40103 30251 40109
rect 30193 40100 30205 40103
rect 29288 40072 30205 40100
rect 28905 40063 28963 40069
rect 30193 40069 30205 40072
rect 30239 40100 30251 40103
rect 30392 40100 30420 40140
rect 32214 40128 32220 40140
rect 32272 40128 32278 40180
rect 32490 40128 32496 40180
rect 32548 40168 32554 40180
rect 35345 40171 35403 40177
rect 32548 40140 35296 40168
rect 32548 40128 32554 40140
rect 30239 40072 30420 40100
rect 30239 40069 30251 40072
rect 30193 40063 30251 40069
rect 24118 40032 24124 40044
rect 23532 40004 24026 40032
rect 24079 40004 24124 40032
rect 23532 39992 23538 40004
rect 24118 39992 24124 40004
rect 24176 39992 24182 40044
rect 24762 39992 24768 40044
rect 24820 40032 24826 40044
rect 25015 40035 25073 40041
rect 25015 40032 25027 40035
rect 24820 40004 25027 40032
rect 24820 39992 24826 40004
rect 25015 40001 25027 40004
rect 25061 40001 25073 40035
rect 25015 39995 25073 40001
rect 25225 40035 25283 40041
rect 25225 40001 25237 40035
rect 25271 40032 25283 40035
rect 25866 40032 25872 40044
rect 25271 40004 25872 40032
rect 25271 40001 25283 40004
rect 25225 39995 25283 40001
rect 25866 39992 25872 40004
rect 25924 39992 25930 40044
rect 26234 39992 26240 40044
rect 26292 40032 26298 40044
rect 26329 40035 26387 40041
rect 26329 40032 26341 40035
rect 26292 40004 26341 40032
rect 26292 39992 26298 40004
rect 26329 40001 26341 40004
rect 26375 40001 26387 40035
rect 26329 39995 26387 40001
rect 26513 40035 26571 40041
rect 26513 40001 26525 40035
rect 26559 40032 26571 40035
rect 27062 40032 27068 40044
rect 26559 40004 27068 40032
rect 26559 40001 26571 40004
rect 26513 39995 26571 40001
rect 27062 39992 27068 40004
rect 27120 39992 27126 40044
rect 27525 40035 27583 40041
rect 27525 40032 27537 40035
rect 27172 40004 27537 40032
rect 17865 39967 17923 39973
rect 17865 39933 17877 39967
rect 17911 39964 17923 39967
rect 18340 39964 18368 39992
rect 17911 39936 18368 39964
rect 20916 39964 20944 39992
rect 23109 39967 23167 39973
rect 23109 39964 23121 39967
rect 20916 39936 23121 39964
rect 17911 39933 17923 39936
rect 17865 39927 17923 39933
rect 23109 39933 23121 39936
rect 23155 39964 23167 39967
rect 23382 39964 23388 39976
rect 23155 39936 23388 39964
rect 23155 39933 23167 39936
rect 23109 39927 23167 39933
rect 23382 39924 23388 39936
rect 23440 39924 23446 39976
rect 24394 39964 24400 39976
rect 24355 39936 24400 39964
rect 24394 39924 24400 39936
rect 24452 39924 24458 39976
rect 25130 39964 25136 39976
rect 25091 39936 25136 39964
rect 25130 39924 25136 39936
rect 25188 39924 25194 39976
rect 25317 39967 25375 39973
rect 25317 39933 25329 39967
rect 25363 39933 25375 39967
rect 25317 39927 25375 39933
rect 19426 39896 19432 39908
rect 18524 39868 19432 39896
rect 18524 39837 18552 39868
rect 19426 39856 19432 39868
rect 19484 39856 19490 39908
rect 22094 39856 22100 39908
rect 22152 39896 22158 39908
rect 23474 39896 23480 39908
rect 22152 39868 23480 39896
rect 22152 39856 22158 39868
rect 23474 39856 23480 39868
rect 23532 39856 23538 39908
rect 25038 39856 25044 39908
rect 25096 39896 25102 39908
rect 25332 39896 25360 39927
rect 25682 39924 25688 39976
rect 25740 39964 25746 39976
rect 26605 39967 26663 39973
rect 25740 39936 26556 39964
rect 25740 39924 25746 39936
rect 25096 39868 25360 39896
rect 26528 39896 26556 39936
rect 26605 39933 26617 39967
rect 26651 39964 26663 39967
rect 26970 39964 26976 39976
rect 26651 39936 26976 39964
rect 26651 39933 26663 39936
rect 26605 39927 26663 39933
rect 26970 39924 26976 39936
rect 27028 39924 27034 39976
rect 27172 39964 27200 40004
rect 27525 40001 27537 40004
rect 27571 40032 27583 40035
rect 28690 40032 28718 40060
rect 28810 40032 28816 40044
rect 27571 40004 28718 40032
rect 28771 40004 28816 40032
rect 27571 40001 27583 40004
rect 27525 39995 27583 40001
rect 28810 39992 28816 40004
rect 28868 39992 28874 40044
rect 27338 39964 27344 39976
rect 27080 39936 27200 39964
rect 27299 39936 27344 39964
rect 27080 39896 27108 39936
rect 27338 39924 27344 39936
rect 27396 39924 27402 39976
rect 27430 39924 27436 39976
rect 27488 39964 27494 39976
rect 27488 39936 27533 39964
rect 27488 39924 27494 39936
rect 27614 39924 27620 39976
rect 27672 39964 27678 39976
rect 27672 39936 27717 39964
rect 27672 39924 27678 39936
rect 27798 39924 27804 39976
rect 27856 39964 27862 39976
rect 27982 39964 27988 39976
rect 27856 39936 27988 39964
rect 27856 39924 27862 39936
rect 27982 39924 27988 39936
rect 28040 39924 28046 39976
rect 28920 39964 28948 40063
rect 32122 40060 32128 40112
rect 32180 40100 32186 40112
rect 33318 40100 33324 40112
rect 32180 40072 32444 40100
rect 32180 40060 32186 40072
rect 28994 39992 29000 40044
rect 29052 40032 29058 40044
rect 29178 40032 29184 40044
rect 29052 40004 29097 40032
rect 29139 40004 29184 40032
rect 29052 39992 29058 40004
rect 29178 39992 29184 40004
rect 29236 39992 29242 40044
rect 29273 40035 29331 40041
rect 29273 40001 29285 40035
rect 29319 40032 29331 40035
rect 31297 40035 31355 40041
rect 29319 40004 29868 40032
rect 29319 40001 29331 40004
rect 29273 39995 29331 40001
rect 29730 39964 29736 39976
rect 28920 39936 29736 39964
rect 29730 39924 29736 39936
rect 29788 39924 29794 39976
rect 29840 39905 29868 40004
rect 31297 40001 31309 40035
rect 31343 40032 31355 40035
rect 31478 40032 31484 40044
rect 31343 40004 31484 40032
rect 31343 40001 31355 40004
rect 31297 39995 31355 40001
rect 31478 39992 31484 40004
rect 31536 39992 31542 40044
rect 31754 39992 31760 40044
rect 31812 40032 31818 40044
rect 32309 40035 32367 40041
rect 32309 40032 32321 40035
rect 31812 40004 32321 40032
rect 31812 39992 31818 40004
rect 32309 40001 32321 40004
rect 32355 40001 32367 40035
rect 32416 40032 32444 40072
rect 32692 40072 33324 40100
rect 32692 40041 32720 40072
rect 33318 40060 33324 40072
rect 33376 40060 33382 40112
rect 35268 40100 35296 40140
rect 35345 40137 35357 40171
rect 35391 40168 35403 40171
rect 35434 40168 35440 40180
rect 35391 40140 35440 40168
rect 35391 40137 35403 40140
rect 35345 40131 35403 40137
rect 35434 40128 35440 40140
rect 35492 40128 35498 40180
rect 35710 40100 35716 40112
rect 35268 40072 35716 40100
rect 35710 40060 35716 40072
rect 35768 40100 35774 40112
rect 35768 40072 36032 40100
rect 35768 40060 35774 40072
rect 32493 40035 32551 40041
rect 32493 40032 32505 40035
rect 32416 40004 32505 40032
rect 32309 39995 32367 40001
rect 32493 40001 32505 40004
rect 32539 40001 32551 40035
rect 32493 39995 32551 40001
rect 32585 40035 32643 40041
rect 32585 40001 32597 40035
rect 32631 40001 32643 40035
rect 32585 39995 32643 40001
rect 32677 40035 32735 40041
rect 32677 40001 32689 40035
rect 32723 40001 32735 40035
rect 35802 40032 35808 40044
rect 35006 40004 35808 40032
rect 32677 39995 32735 40001
rect 31205 39967 31263 39973
rect 31205 39933 31217 39967
rect 31251 39964 31263 39967
rect 31251 39936 31754 39964
rect 31251 39933 31263 39936
rect 31205 39927 31263 39933
rect 29825 39899 29883 39905
rect 26528 39868 27108 39896
rect 28552 39868 28948 39896
rect 25096 39856 25102 39868
rect 18509 39831 18567 39837
rect 18509 39797 18521 39831
rect 18555 39797 18567 39831
rect 18509 39791 18567 39797
rect 18598 39788 18604 39840
rect 18656 39828 18662 39840
rect 18785 39831 18843 39837
rect 18785 39828 18797 39831
rect 18656 39800 18797 39828
rect 18656 39788 18662 39800
rect 18785 39797 18797 39800
rect 18831 39797 18843 39831
rect 18785 39791 18843 39797
rect 20990 39788 20996 39840
rect 21048 39828 21054 39840
rect 21453 39831 21511 39837
rect 21453 39828 21465 39831
rect 21048 39800 21465 39828
rect 21048 39788 21054 39800
rect 21453 39797 21465 39800
rect 21499 39828 21511 39831
rect 21818 39828 21824 39840
rect 21499 39800 21824 39828
rect 21499 39797 21511 39800
rect 21453 39791 21511 39797
rect 21818 39788 21824 39800
rect 21876 39788 21882 39840
rect 22370 39828 22376 39840
rect 22331 39800 22376 39828
rect 22370 39788 22376 39800
rect 22428 39788 22434 39840
rect 22462 39788 22468 39840
rect 22520 39828 22526 39840
rect 23201 39831 23259 39837
rect 23201 39828 23213 39831
rect 22520 39800 23213 39828
rect 22520 39788 22526 39800
rect 23201 39797 23213 39800
rect 23247 39797 23259 39831
rect 23934 39828 23940 39840
rect 23895 39800 23940 39828
rect 23201 39791 23259 39797
rect 23934 39788 23940 39800
rect 23992 39788 23998 39840
rect 24305 39831 24363 39837
rect 24305 39797 24317 39831
rect 24351 39828 24363 39831
rect 24857 39831 24915 39837
rect 24857 39828 24869 39831
rect 24351 39800 24869 39828
rect 24351 39797 24363 39800
rect 24305 39791 24363 39797
rect 24857 39797 24869 39800
rect 24903 39797 24915 39831
rect 24857 39791 24915 39797
rect 24946 39788 24952 39840
rect 25004 39828 25010 39840
rect 26145 39831 26203 39837
rect 26145 39828 26157 39831
rect 25004 39800 26157 39828
rect 25004 39788 25010 39800
rect 26145 39797 26157 39800
rect 26191 39797 26203 39831
rect 26145 39791 26203 39797
rect 27157 39831 27215 39837
rect 27157 39797 27169 39831
rect 27203 39828 27215 39831
rect 27430 39828 27436 39840
rect 27203 39800 27436 39828
rect 27203 39797 27215 39800
rect 27157 39791 27215 39797
rect 27430 39788 27436 39800
rect 27488 39788 27494 39840
rect 27522 39788 27528 39840
rect 27580 39828 27586 39840
rect 28552 39828 28580 39868
rect 27580 39800 28580 39828
rect 27580 39788 27586 39800
rect 28626 39788 28632 39840
rect 28684 39828 28690 39840
rect 28920 39828 28948 39868
rect 29825 39865 29837 39899
rect 29871 39865 29883 39899
rect 31726 39896 31754 39936
rect 32122 39924 32128 39976
rect 32180 39964 32186 39976
rect 32600 39964 32628 39995
rect 35802 39992 35808 40004
rect 35860 39992 35866 40044
rect 36004 40041 36032 40072
rect 35989 40035 36047 40041
rect 35989 40001 36001 40035
rect 36035 40001 36047 40035
rect 35989 39995 36047 40001
rect 32180 39936 32628 39964
rect 33597 39967 33655 39973
rect 32180 39924 32186 39936
rect 33597 39933 33609 39967
rect 33643 39933 33655 39967
rect 33870 39964 33876 39976
rect 33831 39936 33876 39964
rect 33597 39927 33655 39933
rect 33502 39896 33508 39908
rect 31726 39868 33508 39896
rect 29825 39859 29883 39865
rect 33502 39856 33508 39868
rect 33560 39856 33566 39908
rect 29546 39828 29552 39840
rect 28684 39800 28729 39828
rect 28920 39800 29552 39828
rect 28684 39788 28690 39800
rect 29546 39788 29552 39800
rect 29604 39788 29610 39840
rect 30006 39828 30012 39840
rect 29967 39800 30012 39828
rect 30006 39788 30012 39800
rect 30064 39788 30070 39840
rect 30098 39788 30104 39840
rect 30156 39828 30162 39840
rect 30929 39831 30987 39837
rect 30929 39828 30941 39831
rect 30156 39800 30941 39828
rect 30156 39788 30162 39800
rect 30929 39797 30941 39800
rect 30975 39797 30987 39831
rect 30929 39791 30987 39797
rect 31297 39831 31355 39837
rect 31297 39797 31309 39831
rect 31343 39828 31355 39831
rect 31570 39828 31576 39840
rect 31343 39800 31576 39828
rect 31343 39797 31355 39800
rect 31297 39791 31355 39797
rect 31570 39788 31576 39800
rect 31628 39788 31634 39840
rect 32214 39788 32220 39840
rect 32272 39828 32278 39840
rect 32953 39831 33011 39837
rect 32953 39828 32965 39831
rect 32272 39800 32965 39828
rect 32272 39788 32278 39800
rect 32953 39797 32965 39800
rect 32999 39797 33011 39831
rect 33612 39828 33640 39927
rect 33870 39924 33876 39936
rect 33928 39924 33934 39976
rect 35894 39964 35900 39976
rect 35855 39936 35900 39964
rect 35894 39924 35900 39936
rect 35952 39924 35958 39976
rect 35710 39828 35716 39840
rect 33612 39800 35716 39828
rect 32953 39791 33011 39797
rect 35710 39788 35716 39800
rect 35768 39788 35774 39840
rect 36078 39788 36084 39840
rect 36136 39828 36142 39840
rect 36265 39831 36323 39837
rect 36265 39828 36277 39831
rect 36136 39800 36277 39828
rect 36136 39788 36142 39800
rect 36265 39797 36277 39800
rect 36311 39797 36323 39831
rect 36265 39791 36323 39797
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 18506 39624 18512 39636
rect 18467 39596 18512 39624
rect 18506 39584 18512 39596
rect 18564 39584 18570 39636
rect 18690 39584 18696 39636
rect 18748 39624 18754 39636
rect 18748 39596 19334 39624
rect 18748 39584 18754 39596
rect 19306 39556 19334 39596
rect 23382 39584 23388 39636
rect 23440 39624 23446 39636
rect 26050 39624 26056 39636
rect 23440 39596 26056 39624
rect 23440 39584 23446 39596
rect 26050 39584 26056 39596
rect 26108 39584 26114 39636
rect 26145 39627 26203 39633
rect 26145 39593 26157 39627
rect 26191 39624 26203 39627
rect 27338 39624 27344 39636
rect 26191 39596 27344 39624
rect 26191 39593 26203 39596
rect 26145 39587 26203 39593
rect 27338 39584 27344 39596
rect 27396 39584 27402 39636
rect 27525 39627 27583 39633
rect 27525 39593 27537 39627
rect 27571 39624 27583 39627
rect 27614 39624 27620 39636
rect 27571 39596 27620 39624
rect 27571 39593 27583 39596
rect 27525 39587 27583 39593
rect 27614 39584 27620 39596
rect 27672 39584 27678 39636
rect 28350 39624 28356 39636
rect 27816 39596 28356 39624
rect 20898 39556 20904 39568
rect 19306 39528 20904 39556
rect 20898 39516 20904 39528
rect 20956 39556 20962 39568
rect 21634 39556 21640 39568
rect 20956 39528 21640 39556
rect 20956 39516 20962 39528
rect 17773 39491 17831 39497
rect 17773 39457 17785 39491
rect 17819 39488 17831 39491
rect 20346 39488 20352 39500
rect 17819 39460 20352 39488
rect 17819 39457 17831 39460
rect 17773 39451 17831 39457
rect 20346 39448 20352 39460
rect 20404 39488 20410 39500
rect 21100 39497 21128 39528
rect 21634 39516 21640 39528
rect 21692 39516 21698 39568
rect 21818 39516 21824 39568
rect 21876 39556 21882 39568
rect 25130 39556 25136 39568
rect 21876 39528 24992 39556
rect 25091 39528 25136 39556
rect 21876 39516 21882 39528
rect 21085 39491 21143 39497
rect 20404 39460 20852 39488
rect 20404 39448 20410 39460
rect 20162 39420 20168 39432
rect 17328 39392 18736 39420
rect 20123 39392 20168 39420
rect 17328 39296 17356 39392
rect 18493 39355 18551 39361
rect 18493 39321 18505 39355
rect 18539 39352 18551 39355
rect 18598 39352 18604 39364
rect 18539 39324 18604 39352
rect 18539 39321 18551 39324
rect 18493 39315 18551 39321
rect 18598 39312 18604 39324
rect 18656 39312 18662 39364
rect 18708 39361 18736 39392
rect 20162 39380 20168 39392
rect 20220 39380 20226 39432
rect 20254 39380 20260 39432
rect 20312 39420 20318 39432
rect 20824 39429 20852 39460
rect 21085 39457 21097 39491
rect 21131 39457 21143 39491
rect 21085 39451 21143 39457
rect 22094 39448 22100 39500
rect 22152 39488 22158 39500
rect 22649 39491 22707 39497
rect 22649 39488 22661 39491
rect 22152 39460 22661 39488
rect 22152 39448 22158 39460
rect 22649 39457 22661 39460
rect 22695 39457 22707 39491
rect 22649 39451 22707 39457
rect 20717 39423 20775 39429
rect 20312 39392 20357 39420
rect 20312 39380 20318 39392
rect 20717 39389 20729 39423
rect 20763 39389 20775 39423
rect 20717 39383 20775 39389
rect 20809 39423 20867 39429
rect 20809 39389 20821 39423
rect 20855 39420 20867 39423
rect 21174 39420 21180 39432
rect 20855 39392 21180 39420
rect 20855 39389 20867 39392
rect 20809 39383 20867 39389
rect 18693 39355 18751 39361
rect 18693 39321 18705 39355
rect 18739 39321 18751 39355
rect 20732 39352 20760 39383
rect 21174 39380 21180 39392
rect 21232 39380 21238 39432
rect 21358 39420 21364 39432
rect 21319 39392 21364 39420
rect 21358 39380 21364 39392
rect 21416 39380 21422 39432
rect 21542 39380 21548 39432
rect 21600 39420 21606 39432
rect 22373 39423 22431 39429
rect 22373 39420 22385 39423
rect 21600 39392 22385 39420
rect 21600 39380 21606 39392
rect 22373 39389 22385 39392
rect 22419 39420 22431 39423
rect 22557 39423 22615 39429
rect 22419 39392 22508 39420
rect 22419 39389 22431 39392
rect 22373 39383 22431 39389
rect 22189 39355 22247 39361
rect 22189 39352 22201 39355
rect 20732 39324 22201 39352
rect 18693 39315 18751 39321
rect 22189 39321 22201 39324
rect 22235 39321 22247 39355
rect 22189 39315 22247 39321
rect 16485 39287 16543 39293
rect 16485 39253 16497 39287
rect 16531 39284 16543 39287
rect 16574 39284 16580 39296
rect 16531 39256 16580 39284
rect 16531 39253 16543 39256
rect 16485 39247 16543 39253
rect 16574 39244 16580 39256
rect 16632 39284 16638 39296
rect 17310 39284 17316 39296
rect 16632 39256 17316 39284
rect 16632 39244 16638 39256
rect 17310 39244 17316 39256
rect 17368 39244 17374 39296
rect 18046 39244 18052 39296
rect 18104 39284 18110 39296
rect 18325 39287 18383 39293
rect 18325 39284 18337 39287
rect 18104 39256 18337 39284
rect 18104 39244 18110 39256
rect 18325 39253 18337 39256
rect 18371 39253 18383 39287
rect 18325 39247 18383 39253
rect 20714 39244 20720 39296
rect 20772 39284 20778 39296
rect 21450 39284 21456 39296
rect 20772 39256 21456 39284
rect 20772 39244 20778 39256
rect 21450 39244 21456 39256
rect 21508 39244 21514 39296
rect 22480 39284 22508 39392
rect 22557 39389 22569 39423
rect 22603 39389 22615 39423
rect 22738 39420 22744 39432
rect 22699 39392 22744 39420
rect 22557 39383 22615 39389
rect 22572 39352 22600 39383
rect 22738 39380 22744 39392
rect 22796 39380 22802 39432
rect 22922 39420 22928 39432
rect 22883 39392 22928 39420
rect 22922 39380 22928 39392
rect 22980 39380 22986 39432
rect 23382 39380 23388 39432
rect 23440 39420 23446 39432
rect 23569 39423 23627 39429
rect 23569 39420 23581 39423
rect 23440 39392 23581 39420
rect 23440 39380 23446 39392
rect 23569 39389 23581 39392
rect 23615 39389 23627 39423
rect 23569 39383 23627 39389
rect 23753 39423 23811 39429
rect 23753 39389 23765 39423
rect 23799 39420 23811 39423
rect 24854 39420 24860 39432
rect 23799 39392 24860 39420
rect 23799 39389 23811 39392
rect 23753 39383 23811 39389
rect 24854 39380 24860 39392
rect 24912 39380 24918 39432
rect 24964 39420 24992 39528
rect 25130 39516 25136 39528
rect 25188 39516 25194 39568
rect 27816 39556 27844 39596
rect 28350 39584 28356 39596
rect 28408 39584 28414 39636
rect 28537 39627 28595 39633
rect 28537 39593 28549 39627
rect 28583 39624 28595 39627
rect 28810 39624 28816 39636
rect 28583 39596 28816 39624
rect 28583 39593 28595 39596
rect 28537 39587 28595 39593
rect 28810 39584 28816 39596
rect 28868 39584 28874 39636
rect 30558 39584 30564 39636
rect 30616 39624 30622 39636
rect 30926 39624 30932 39636
rect 30616 39596 30932 39624
rect 30616 39584 30622 39596
rect 30926 39584 30932 39596
rect 30984 39584 30990 39636
rect 32122 39584 32128 39636
rect 32180 39624 32186 39636
rect 32585 39627 32643 39633
rect 32585 39624 32597 39627
rect 32180 39596 32597 39624
rect 32180 39584 32186 39596
rect 32585 39593 32597 39596
rect 32631 39593 32643 39627
rect 32585 39587 32643 39593
rect 27893 39559 27951 39565
rect 27893 39556 27905 39559
rect 27816 39528 27905 39556
rect 27893 39525 27905 39528
rect 27939 39525 27951 39559
rect 27893 39519 27951 39525
rect 28166 39516 28172 39568
rect 28224 39516 28230 39568
rect 29822 39516 29828 39568
rect 29880 39556 29886 39568
rect 32490 39556 32496 39568
rect 29880 39528 32496 39556
rect 29880 39516 29886 39528
rect 32490 39516 32496 39528
rect 32548 39516 32554 39568
rect 32950 39556 32956 39568
rect 32600 39528 32956 39556
rect 27062 39448 27068 39500
rect 27120 39488 27126 39500
rect 28184 39488 28212 39516
rect 30282 39488 30288 39500
rect 27120 39460 27936 39488
rect 27120 39448 27126 39460
rect 24964 39392 25176 39420
rect 23842 39352 23848 39364
rect 22572 39324 23848 39352
rect 23842 39312 23848 39324
rect 23900 39312 23906 39364
rect 25148 39361 25176 39392
rect 25222 39380 25228 39432
rect 25280 39420 25286 39432
rect 25869 39423 25927 39429
rect 25869 39420 25881 39423
rect 25280 39392 25881 39420
rect 25280 39380 25286 39392
rect 25869 39389 25881 39392
rect 25915 39389 25927 39423
rect 26142 39420 26148 39432
rect 26103 39392 26148 39420
rect 25869 39383 25927 39389
rect 26142 39380 26148 39392
rect 26200 39380 26206 39432
rect 26605 39423 26663 39429
rect 26605 39420 26617 39423
rect 26344 39392 26617 39420
rect 25133 39355 25191 39361
rect 25133 39321 25145 39355
rect 25179 39352 25191 39355
rect 25406 39352 25412 39364
rect 25179 39324 25412 39352
rect 25179 39321 25191 39324
rect 25133 39315 25191 39321
rect 25406 39312 25412 39324
rect 25464 39312 25470 39364
rect 25682 39312 25688 39364
rect 25740 39352 25746 39364
rect 26053 39355 26111 39361
rect 26053 39352 26065 39355
rect 25740 39324 26065 39352
rect 25740 39312 25746 39324
rect 26053 39321 26065 39324
rect 26099 39321 26111 39355
rect 26053 39315 26111 39321
rect 22830 39284 22836 39296
rect 22480 39256 22836 39284
rect 22830 39244 22836 39256
rect 22888 39244 22894 39296
rect 23382 39284 23388 39296
rect 23343 39256 23388 39284
rect 23382 39244 23388 39256
rect 23440 39244 23446 39296
rect 23750 39244 23756 39296
rect 23808 39284 23814 39296
rect 24026 39284 24032 39296
rect 23808 39256 24032 39284
rect 23808 39244 23814 39256
rect 24026 39244 24032 39256
rect 24084 39284 24090 39296
rect 24949 39287 25007 39293
rect 24949 39284 24961 39287
rect 24084 39256 24961 39284
rect 24084 39244 24090 39256
rect 24949 39253 24961 39256
rect 24995 39284 25007 39287
rect 26344 39284 26372 39392
rect 26605 39389 26617 39392
rect 26651 39389 26663 39423
rect 26605 39383 26663 39389
rect 26789 39423 26847 39429
rect 26789 39389 26801 39423
rect 26835 39389 26847 39423
rect 26789 39383 26847 39389
rect 26510 39312 26516 39364
rect 26568 39352 26574 39364
rect 26804 39352 26832 39383
rect 27614 39380 27620 39432
rect 27672 39420 27678 39432
rect 27709 39423 27767 39429
rect 27709 39420 27721 39423
rect 27672 39392 27721 39420
rect 27672 39380 27678 39392
rect 27709 39389 27721 39392
rect 27755 39389 27767 39423
rect 27709 39383 27767 39389
rect 27801 39423 27859 39429
rect 27801 39389 27813 39423
rect 27847 39389 27859 39423
rect 27908 39418 27936 39460
rect 28092 39460 28212 39488
rect 28920 39460 30288 39488
rect 27985 39423 28043 39429
rect 27985 39418 27997 39423
rect 27908 39390 27997 39418
rect 27801 39383 27859 39389
rect 27985 39389 27997 39390
rect 28031 39420 28043 39423
rect 28092 39420 28120 39460
rect 28031 39392 28120 39420
rect 28031 39389 28043 39392
rect 27985 39383 28043 39389
rect 27816 39352 27844 39383
rect 28166 39380 28172 39432
rect 28224 39420 28230 39432
rect 28920 39429 28948 39460
rect 30282 39448 30288 39460
rect 30340 39488 30346 39500
rect 30653 39491 30711 39497
rect 30653 39488 30665 39491
rect 30340 39460 30665 39488
rect 30340 39448 30346 39460
rect 30653 39457 30665 39460
rect 30699 39457 30711 39491
rect 30653 39451 30711 39457
rect 30926 39448 30932 39500
rect 30984 39488 30990 39500
rect 32600 39488 32628 39528
rect 32766 39488 32772 39500
rect 30984 39460 32628 39488
rect 32727 39460 32772 39488
rect 30984 39448 30990 39460
rect 32766 39448 32772 39460
rect 32824 39448 32830 39500
rect 32876 39497 32904 39528
rect 32950 39516 32956 39528
rect 33008 39516 33014 39568
rect 32861 39491 32919 39497
rect 32861 39457 32873 39491
rect 32907 39457 32919 39491
rect 32861 39451 32919 39457
rect 35434 39448 35440 39500
rect 35492 39488 35498 39500
rect 35710 39488 35716 39500
rect 35492 39460 35716 39488
rect 35492 39448 35498 39460
rect 35710 39448 35716 39460
rect 35768 39448 35774 39500
rect 35894 39488 35900 39500
rect 35866 39448 35900 39488
rect 35952 39448 35958 39500
rect 36078 39488 36084 39500
rect 36039 39460 36084 39488
rect 36078 39448 36084 39460
rect 36136 39448 36142 39500
rect 37458 39488 37464 39500
rect 37419 39460 37464 39488
rect 37458 39448 37464 39460
rect 37516 39448 37522 39500
rect 28675 39423 28733 39429
rect 28675 39420 28687 39423
rect 28224 39392 28687 39420
rect 28224 39380 28230 39392
rect 28675 39389 28687 39392
rect 28721 39389 28733 39423
rect 28675 39383 28733 39389
rect 28905 39423 28963 39429
rect 28905 39389 28917 39423
rect 28951 39389 28963 39423
rect 29086 39420 29092 39432
rect 29047 39392 29092 39420
rect 28905 39383 28963 39389
rect 29086 39380 29092 39392
rect 29144 39380 29150 39432
rect 29181 39423 29239 39429
rect 29181 39389 29193 39423
rect 29227 39420 29239 39423
rect 29270 39420 29276 39432
rect 29227 39392 29276 39420
rect 29227 39389 29239 39392
rect 29181 39383 29239 39389
rect 29270 39380 29276 39392
rect 29328 39380 29334 39432
rect 29730 39420 29736 39432
rect 29691 39392 29736 39420
rect 29730 39380 29736 39392
rect 29788 39380 29794 39432
rect 29822 39380 29828 39432
rect 29880 39420 29886 39432
rect 29917 39423 29975 39429
rect 29917 39420 29929 39423
rect 29880 39392 29929 39420
rect 29880 39380 29886 39392
rect 29917 39389 29929 39392
rect 29963 39389 29975 39423
rect 30374 39420 30380 39432
rect 29917 39383 29975 39389
rect 30024 39392 30380 39420
rect 26568 39324 26832 39352
rect 27724 39324 27844 39352
rect 28813 39355 28871 39361
rect 26568 39312 26574 39324
rect 27724 39296 27752 39324
rect 28813 39321 28825 39355
rect 28859 39352 28871 39355
rect 30024 39352 30052 39392
rect 30374 39380 30380 39392
rect 30432 39420 30438 39432
rect 30561 39423 30619 39429
rect 30561 39420 30573 39423
rect 30432 39392 30573 39420
rect 30432 39380 30438 39392
rect 30561 39389 30573 39392
rect 30607 39389 30619 39423
rect 30561 39383 30619 39389
rect 30745 39423 30803 39429
rect 30745 39389 30757 39423
rect 30791 39420 30803 39423
rect 31202 39420 31208 39432
rect 30791 39392 31208 39420
rect 30791 39389 30803 39392
rect 30745 39383 30803 39389
rect 28859 39324 30052 39352
rect 28859 39321 28871 39324
rect 28813 39315 28871 39321
rect 30098 39312 30104 39364
rect 30156 39352 30162 39364
rect 30576 39352 30604 39383
rect 31202 39380 31208 39392
rect 31260 39380 31266 39432
rect 31297 39423 31355 39429
rect 31297 39389 31309 39423
rect 31343 39420 31355 39423
rect 32490 39420 32496 39432
rect 31343 39392 32496 39420
rect 31343 39389 31355 39392
rect 31297 39383 31355 39389
rect 31312 39352 31340 39383
rect 32490 39380 32496 39392
rect 32548 39380 32554 39432
rect 32953 39423 33011 39429
rect 32953 39420 32965 39423
rect 32876 39392 32965 39420
rect 32876 39364 32904 39392
rect 32953 39389 32965 39392
rect 32999 39389 33011 39423
rect 32953 39383 33011 39389
rect 33045 39423 33103 39429
rect 33045 39389 33057 39423
rect 33091 39420 33103 39423
rect 33502 39420 33508 39432
rect 33091 39392 33508 39420
rect 33091 39389 33103 39392
rect 33045 39383 33103 39389
rect 33502 39380 33508 39392
rect 33560 39380 33566 39432
rect 34054 39380 34060 39432
rect 34112 39420 34118 39432
rect 34885 39423 34943 39429
rect 34885 39420 34897 39423
rect 34112 39392 34897 39420
rect 34112 39380 34118 39392
rect 34885 39389 34897 39392
rect 34931 39420 34943 39423
rect 35866 39420 35894 39448
rect 34931 39392 35894 39420
rect 34931 39389 34943 39392
rect 34885 39383 34943 39389
rect 32858 39352 32864 39364
rect 30156 39324 30201 39352
rect 30576 39324 31340 39352
rect 31404 39324 32864 39352
rect 30156 39312 30162 39324
rect 26694 39284 26700 39296
rect 24995 39256 26372 39284
rect 26655 39256 26700 39284
rect 24995 39253 25007 39256
rect 24949 39247 25007 39253
rect 26694 39244 26700 39256
rect 26752 39244 26758 39296
rect 26786 39244 26792 39296
rect 26844 39284 26850 39296
rect 26970 39284 26976 39296
rect 26844 39256 26976 39284
rect 26844 39244 26850 39256
rect 26970 39244 26976 39256
rect 27028 39244 27034 39296
rect 27706 39244 27712 39296
rect 27764 39244 27770 39296
rect 27798 39244 27804 39296
rect 27856 39284 27862 39296
rect 29086 39284 29092 39296
rect 27856 39256 29092 39284
rect 27856 39244 27862 39256
rect 29086 39244 29092 39256
rect 29144 39284 29150 39296
rect 31404 39284 31432 39324
rect 32858 39312 32864 39324
rect 32916 39312 32922 39364
rect 34514 39352 34520 39364
rect 32968 39324 34520 39352
rect 32122 39284 32128 39296
rect 29144 39256 31432 39284
rect 32083 39256 32128 39284
rect 29144 39244 29150 39256
rect 32122 39244 32128 39256
rect 32180 39244 32186 39296
rect 32490 39244 32496 39296
rect 32548 39284 32554 39296
rect 32968 39284 32996 39324
rect 34514 39312 34520 39324
rect 34572 39312 34578 39364
rect 36372 39324 36478 39352
rect 33686 39284 33692 39296
rect 32548 39256 32996 39284
rect 33647 39256 33692 39284
rect 32548 39244 32554 39256
rect 33686 39244 33692 39256
rect 33744 39244 33750 39296
rect 34238 39284 34244 39296
rect 34199 39256 34244 39284
rect 34238 39244 34244 39256
rect 34296 39244 34302 39296
rect 35802 39244 35808 39296
rect 35860 39284 35866 39296
rect 36170 39284 36176 39296
rect 35860 39256 36176 39284
rect 35860 39244 35866 39256
rect 36170 39244 36176 39256
rect 36228 39284 36234 39296
rect 36372 39284 36400 39324
rect 36228 39256 36400 39284
rect 36228 39244 36234 39256
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 17954 39040 17960 39092
rect 18012 39080 18018 39092
rect 18141 39083 18199 39089
rect 18141 39080 18153 39083
rect 18012 39052 18153 39080
rect 18012 39040 18018 39052
rect 18141 39049 18153 39052
rect 18187 39080 18199 39083
rect 18506 39080 18512 39092
rect 18187 39052 18512 39080
rect 18187 39049 18199 39052
rect 18141 39043 18199 39049
rect 18506 39040 18512 39052
rect 18564 39040 18570 39092
rect 18690 39080 18696 39092
rect 18651 39052 18696 39080
rect 18690 39040 18696 39052
rect 18748 39040 18754 39092
rect 20162 39040 20168 39092
rect 20220 39080 20226 39092
rect 20257 39083 20315 39089
rect 20257 39080 20269 39083
rect 20220 39052 20269 39080
rect 20220 39040 20226 39052
rect 20257 39049 20269 39052
rect 20303 39049 20315 39083
rect 20438 39080 20444 39092
rect 20257 39043 20315 39049
rect 20364 39052 20444 39080
rect 16853 39015 16911 39021
rect 16853 39012 16865 39015
rect 16132 38984 16865 39012
rect 16132 38953 16160 38984
rect 16853 38981 16865 38984
rect 16899 38981 16911 39015
rect 19245 39015 19303 39021
rect 16853 38975 16911 38981
rect 17328 38984 18000 39012
rect 16117 38947 16175 38953
rect 16117 38913 16129 38947
rect 16163 38913 16175 38947
rect 16117 38907 16175 38913
rect 16301 38947 16359 38953
rect 16301 38913 16313 38947
rect 16347 38944 16359 38947
rect 16574 38944 16580 38956
rect 16347 38916 16580 38944
rect 16347 38913 16359 38916
rect 16301 38907 16359 38913
rect 16574 38904 16580 38916
rect 16632 38904 16638 38956
rect 17034 38904 17040 38956
rect 17092 38953 17098 38956
rect 17092 38947 17114 38953
rect 17102 38913 17114 38947
rect 17218 38944 17224 38956
rect 17179 38916 17224 38944
rect 17092 38907 17114 38913
rect 17092 38904 17098 38907
rect 17218 38904 17224 38916
rect 17276 38904 17282 38956
rect 17328 38953 17356 38984
rect 17972 38953 18000 38984
rect 19245 38981 19257 39015
rect 19291 39012 19303 39015
rect 20364 39012 20392 39052
rect 20438 39040 20444 39052
rect 20496 39080 20502 39092
rect 21361 39083 21419 39089
rect 21361 39080 21373 39083
rect 20496 39052 21373 39080
rect 20496 39040 20502 39052
rect 21361 39049 21373 39052
rect 21407 39080 21419 39083
rect 22094 39080 22100 39092
rect 21407 39052 22100 39080
rect 21407 39049 21419 39052
rect 21361 39043 21419 39049
rect 22094 39040 22100 39052
rect 22152 39080 22158 39092
rect 22152 39052 24164 39080
rect 22152 39040 22158 39052
rect 20806 39012 20812 39024
rect 19291 38984 20392 39012
rect 20456 38984 20812 39012
rect 19291 38981 19303 38984
rect 19245 38975 19303 38981
rect 20456 38953 20484 38984
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 21174 38972 21180 39024
rect 21232 39012 21238 39024
rect 21634 39012 21640 39024
rect 21232 38984 21640 39012
rect 21232 38972 21238 38984
rect 21634 38972 21640 38984
rect 21692 39012 21698 39024
rect 22373 39015 22431 39021
rect 22373 39012 22385 39015
rect 21692 38984 22385 39012
rect 21692 38972 21698 38984
rect 22373 38981 22385 38984
rect 22419 38981 22431 39015
rect 23290 39012 23296 39024
rect 22373 38975 22431 38981
rect 22572 38984 23296 39012
rect 17313 38947 17371 38953
rect 17313 38913 17325 38947
rect 17359 38913 17371 38947
rect 17313 38907 17371 38913
rect 17773 38947 17831 38953
rect 17773 38913 17785 38947
rect 17819 38913 17831 38947
rect 17773 38907 17831 38913
rect 17957 38947 18015 38953
rect 17957 38913 17969 38947
rect 18003 38913 18015 38947
rect 17957 38907 18015 38913
rect 20441 38947 20499 38953
rect 20441 38913 20453 38947
rect 20487 38913 20499 38947
rect 20441 38907 20499 38913
rect 20533 38947 20591 38953
rect 20533 38913 20545 38947
rect 20579 38944 20591 38947
rect 22002 38944 22008 38956
rect 20579 38916 22008 38944
rect 20579 38913 20591 38916
rect 20533 38907 20591 38913
rect 17328 38876 17356 38907
rect 17144 38848 17356 38876
rect 17144 38820 17172 38848
rect 17126 38768 17132 38820
rect 17184 38768 17190 38820
rect 16209 38743 16267 38749
rect 16209 38709 16221 38743
rect 16255 38740 16267 38743
rect 16574 38740 16580 38752
rect 16255 38712 16580 38740
rect 16255 38709 16267 38712
rect 16209 38703 16267 38709
rect 16574 38700 16580 38712
rect 16632 38700 16638 38752
rect 17034 38700 17040 38752
rect 17092 38740 17098 38752
rect 17788 38740 17816 38907
rect 22002 38904 22008 38916
rect 22060 38904 22066 38956
rect 22189 38947 22247 38953
rect 22189 38913 22201 38947
rect 22235 38913 22247 38947
rect 22189 38907 22247 38913
rect 22281 38947 22339 38953
rect 22281 38913 22293 38947
rect 22327 38944 22339 38947
rect 22462 38944 22468 38956
rect 22327 38916 22468 38944
rect 22327 38913 22339 38916
rect 22281 38907 22339 38913
rect 20625 38879 20683 38885
rect 20625 38876 20637 38879
rect 20456 38848 20637 38876
rect 20456 38820 20484 38848
rect 20625 38845 20637 38848
rect 20671 38845 20683 38879
rect 20625 38839 20683 38845
rect 20714 38836 20720 38888
rect 20772 38876 20778 38888
rect 20772 38848 20817 38876
rect 20772 38836 20778 38848
rect 22204 38820 22232 38907
rect 22462 38904 22468 38916
rect 22520 38904 22526 38956
rect 22572 38953 22600 38984
rect 23290 38972 23296 38984
rect 23348 38972 23354 39024
rect 23382 38972 23388 39024
rect 23440 39012 23446 39024
rect 23440 38984 23613 39012
rect 23440 38972 23446 38984
rect 22557 38947 22615 38953
rect 22557 38913 22569 38947
rect 22603 38913 22615 38947
rect 22557 38907 22615 38913
rect 22649 38947 22707 38953
rect 22649 38913 22661 38947
rect 22695 38913 22707 38947
rect 23474 38944 23480 38956
rect 23435 38916 23480 38944
rect 22649 38907 22707 38913
rect 22664 38876 22692 38907
rect 23474 38904 23480 38916
rect 23532 38904 23538 38956
rect 23585 38953 23613 38984
rect 24026 38953 24032 38956
rect 23570 38947 23628 38953
rect 23570 38913 23582 38947
rect 23616 38913 23628 38947
rect 23570 38907 23628 38913
rect 23753 38947 23811 38953
rect 23753 38913 23765 38947
rect 23799 38913 23811 38947
rect 23753 38907 23811 38913
rect 23845 38947 23903 38953
rect 23845 38913 23857 38947
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 23983 38947 24032 38953
rect 23983 38913 23995 38947
rect 24029 38913 24032 38947
rect 23983 38907 24032 38913
rect 23382 38876 23388 38888
rect 22664 38848 23388 38876
rect 23382 38836 23388 38848
rect 23440 38836 23446 38888
rect 23658 38876 23664 38888
rect 23571 38848 23664 38876
rect 20438 38768 20444 38820
rect 20496 38768 20502 38820
rect 21836 38780 22140 38808
rect 17862 38740 17868 38752
rect 17092 38712 17868 38740
rect 17092 38700 17098 38712
rect 17862 38700 17868 38712
rect 17920 38700 17926 38752
rect 19797 38743 19855 38749
rect 19797 38709 19809 38743
rect 19843 38740 19855 38743
rect 21836 38740 21864 38780
rect 22002 38740 22008 38752
rect 19843 38712 21864 38740
rect 21963 38712 22008 38740
rect 19843 38709 19855 38712
rect 19797 38703 19855 38709
rect 22002 38700 22008 38712
rect 22060 38700 22066 38752
rect 22112 38740 22140 38780
rect 22186 38768 22192 38820
rect 22244 38768 22250 38820
rect 23585 38740 23613 38848
rect 23658 38836 23664 38848
rect 23716 38876 23722 38888
rect 23768 38876 23796 38907
rect 23716 38848 23796 38876
rect 23716 38836 23722 38848
rect 22112 38712 23613 38740
rect 23658 38700 23664 38752
rect 23716 38740 23722 38752
rect 23860 38740 23888 38907
rect 24026 38904 24032 38907
rect 24084 38904 24090 38956
rect 24136 38808 24164 39052
rect 24486 39040 24492 39092
rect 24544 39080 24550 39092
rect 26326 39080 26332 39092
rect 24544 39052 26332 39080
rect 24544 39040 24550 39052
rect 26326 39040 26332 39052
rect 26384 39080 26390 39092
rect 26786 39080 26792 39092
rect 26384 39052 26792 39080
rect 26384 39040 26390 39052
rect 26786 39040 26792 39052
rect 26844 39080 26850 39092
rect 27430 39080 27436 39092
rect 26844 39052 27436 39080
rect 26844 39040 26850 39052
rect 27430 39040 27436 39052
rect 27488 39040 27494 39092
rect 27614 39040 27620 39092
rect 27672 39080 27678 39092
rect 30190 39080 30196 39092
rect 27672 39052 30196 39080
rect 27672 39040 27678 39052
rect 30190 39040 30196 39052
rect 30248 39080 30254 39092
rect 30374 39080 30380 39092
rect 30248 39052 30380 39080
rect 30248 39040 30254 39052
rect 30374 39040 30380 39052
rect 30432 39040 30438 39092
rect 30466 39040 30472 39092
rect 30524 39080 30530 39092
rect 32309 39083 32367 39089
rect 32309 39080 32321 39083
rect 30524 39052 31432 39080
rect 30524 39040 30530 39052
rect 26694 39012 26700 39024
rect 25056 38984 26700 39012
rect 25056 38953 25084 38984
rect 26694 38972 26700 38984
rect 26752 38972 26758 39024
rect 27338 38972 27344 39024
rect 27396 39012 27402 39024
rect 27798 39012 27804 39024
rect 27396 38984 27804 39012
rect 27396 38972 27402 38984
rect 27798 38972 27804 38984
rect 27856 39012 27862 39024
rect 28169 39015 28227 39021
rect 28169 39012 28181 39015
rect 27856 38984 28181 39012
rect 27856 38972 27862 38984
rect 28169 38981 28181 38984
rect 28215 38981 28227 39015
rect 28169 38975 28227 38981
rect 28353 39015 28411 39021
rect 28353 38981 28365 39015
rect 28399 38981 28411 39015
rect 28353 38975 28411 38981
rect 25041 38947 25099 38953
rect 25041 38913 25053 38947
rect 25087 38913 25099 38947
rect 25041 38907 25099 38913
rect 25225 38947 25283 38953
rect 25225 38913 25237 38947
rect 25271 38913 25283 38947
rect 25225 38907 25283 38913
rect 25409 38947 25467 38953
rect 25409 38913 25421 38947
rect 25455 38944 25467 38947
rect 26237 38947 26295 38953
rect 26237 38944 26249 38947
rect 25455 38916 26249 38944
rect 25455 38913 25467 38916
rect 25409 38907 25467 38913
rect 26237 38913 26249 38916
rect 26283 38913 26295 38947
rect 26237 38907 26295 38913
rect 26329 38947 26387 38953
rect 26329 38913 26341 38947
rect 26375 38913 26387 38947
rect 26329 38907 26387 38913
rect 26605 38947 26663 38953
rect 26605 38913 26617 38947
rect 26651 38944 26663 38947
rect 26878 38944 26884 38956
rect 26651 38916 26884 38944
rect 26651 38913 26663 38916
rect 26605 38907 26663 38913
rect 24949 38879 25007 38885
rect 24949 38845 24961 38879
rect 24995 38876 25007 38879
rect 25130 38876 25136 38888
rect 24995 38848 25136 38876
rect 24995 38845 25007 38848
rect 24949 38839 25007 38845
rect 25130 38836 25136 38848
rect 25188 38836 25194 38888
rect 25240 38808 25268 38907
rect 26344 38876 26372 38907
rect 26878 38904 26884 38916
rect 26936 38904 26942 38956
rect 27430 38944 27436 38956
rect 27391 38916 27436 38944
rect 27430 38904 27436 38916
rect 27488 38904 27494 38956
rect 28368 38888 28396 38975
rect 28994 38972 29000 39024
rect 29052 39012 29058 39024
rect 29730 39012 29736 39024
rect 29052 38984 29736 39012
rect 29052 38972 29058 38984
rect 29730 38972 29736 38984
rect 29788 38972 29794 39024
rect 31404 39021 31432 39052
rect 31496 39052 32321 39080
rect 31496 39021 31524 39052
rect 32309 39049 32321 39052
rect 32355 39049 32367 39083
rect 32309 39043 32367 39049
rect 32950 39040 32956 39092
rect 33008 39040 33014 39092
rect 33870 39080 33876 39092
rect 33831 39052 33876 39080
rect 33870 39040 33876 39052
rect 33928 39040 33934 39092
rect 34514 39040 34520 39092
rect 34572 39080 34578 39092
rect 36265 39083 36323 39089
rect 36265 39080 36277 39083
rect 34572 39052 36277 39080
rect 34572 39040 34578 39052
rect 36265 39049 36277 39052
rect 36311 39049 36323 39083
rect 36265 39043 36323 39049
rect 31389 39015 31447 39021
rect 31389 38981 31401 39015
rect 31435 38981 31447 39015
rect 31389 38975 31447 38981
rect 31481 39015 31539 39021
rect 31481 38981 31493 39015
rect 31527 38981 31539 39015
rect 32398 39012 32404 39024
rect 31481 38975 31539 38981
rect 31956 38984 32404 39012
rect 28442 38904 28448 38956
rect 28500 38944 28506 38956
rect 28500 38916 28994 38944
rect 28500 38904 28506 38916
rect 27154 38876 27160 38888
rect 26344 38848 27160 38876
rect 27154 38836 27160 38848
rect 27212 38836 27218 38888
rect 27246 38836 27252 38888
rect 27304 38876 27310 38888
rect 27341 38879 27399 38885
rect 27341 38876 27353 38879
rect 27304 38848 27353 38876
rect 27304 38836 27310 38848
rect 27341 38845 27353 38848
rect 27387 38845 27399 38879
rect 27341 38839 27399 38845
rect 27525 38879 27583 38885
rect 27525 38845 27537 38879
rect 27571 38845 27583 38879
rect 27525 38839 27583 38845
rect 27617 38879 27675 38885
rect 27617 38845 27629 38879
rect 27663 38876 27675 38879
rect 27798 38876 27804 38888
rect 27663 38848 27804 38876
rect 27663 38845 27675 38848
rect 27617 38839 27675 38845
rect 24136 38780 25268 38808
rect 26142 38768 26148 38820
rect 26200 38808 26206 38820
rect 27540 38808 27568 38839
rect 27798 38836 27804 38848
rect 27856 38836 27862 38888
rect 28350 38836 28356 38888
rect 28408 38836 28414 38888
rect 28966 38876 28994 38916
rect 29178 38904 29184 38956
rect 29236 38944 29242 38956
rect 29638 38944 29644 38956
rect 29236 38916 29644 38944
rect 29236 38904 29242 38916
rect 29638 38904 29644 38916
rect 29696 38904 29702 38956
rect 29914 38904 29920 38956
rect 29972 38944 29978 38956
rect 30009 38947 30067 38953
rect 30009 38944 30021 38947
rect 29972 38916 30021 38944
rect 29972 38904 29978 38916
rect 30009 38913 30021 38916
rect 30055 38913 30067 38947
rect 30190 38944 30196 38956
rect 30151 38916 30196 38944
rect 30009 38907 30067 38913
rect 30190 38904 30196 38916
rect 30248 38904 30254 38956
rect 30282 38904 30288 38956
rect 30340 38944 30346 38956
rect 30469 38947 30527 38953
rect 30340 38916 30385 38944
rect 30340 38904 30346 38916
rect 30469 38913 30481 38947
rect 30515 38913 30527 38947
rect 31294 38944 31300 38956
rect 31255 38916 31300 38944
rect 30469 38907 30527 38913
rect 29822 38876 29828 38888
rect 28966 38848 29828 38876
rect 29822 38836 29828 38848
rect 29880 38836 29886 38888
rect 27706 38808 27712 38820
rect 26200 38780 27712 38808
rect 26200 38768 26206 38780
rect 27706 38768 27712 38780
rect 27764 38768 27770 38820
rect 28169 38811 28227 38817
rect 28169 38808 28181 38811
rect 27908 38780 28181 38808
rect 24118 38740 24124 38752
rect 23716 38712 23888 38740
rect 24079 38712 24124 38740
rect 23716 38700 23722 38712
rect 24118 38700 24124 38712
rect 24176 38700 24182 38752
rect 26050 38740 26056 38752
rect 26011 38712 26056 38740
rect 26050 38700 26056 38712
rect 26108 38700 26114 38752
rect 26513 38743 26571 38749
rect 26513 38709 26525 38743
rect 26559 38740 26571 38743
rect 26602 38740 26608 38752
rect 26559 38712 26608 38740
rect 26559 38709 26571 38712
rect 26513 38703 26571 38709
rect 26602 38700 26608 38712
rect 26660 38700 26666 38752
rect 27154 38740 27160 38752
rect 27067 38712 27160 38740
rect 27154 38700 27160 38712
rect 27212 38740 27218 38752
rect 27338 38740 27344 38752
rect 27212 38712 27344 38740
rect 27212 38700 27218 38712
rect 27338 38700 27344 38712
rect 27396 38700 27402 38752
rect 27614 38700 27620 38752
rect 27672 38740 27678 38752
rect 27908 38740 27936 38780
rect 28169 38777 28181 38780
rect 28215 38777 28227 38811
rect 28169 38771 28227 38777
rect 28997 38811 29055 38817
rect 28997 38777 29009 38811
rect 29043 38808 29055 38811
rect 29730 38808 29736 38820
rect 29043 38780 29736 38808
rect 29043 38777 29055 38780
rect 28997 38771 29055 38777
rect 29730 38768 29736 38780
rect 29788 38768 29794 38820
rect 30377 38811 30435 38817
rect 30377 38777 30389 38811
rect 30423 38777 30435 38811
rect 30484 38808 30512 38907
rect 31294 38904 31300 38916
rect 31352 38904 31358 38956
rect 31665 38947 31723 38953
rect 31665 38913 31677 38947
rect 31711 38913 31723 38947
rect 31665 38907 31723 38913
rect 30653 38879 30711 38885
rect 30653 38845 30665 38879
rect 30699 38876 30711 38879
rect 31680 38876 31708 38907
rect 31956 38876 31984 38984
rect 32398 38972 32404 38984
rect 32456 39012 32462 39024
rect 32677 39015 32735 39021
rect 32677 39012 32689 39015
rect 32456 38984 32689 39012
rect 32456 38972 32462 38984
rect 32677 38981 32689 38984
rect 32723 38981 32735 39015
rect 32968 39012 32996 39040
rect 36354 39012 36360 39024
rect 32677 38975 32735 38981
rect 32876 38984 32996 39012
rect 33244 38984 36360 39012
rect 32122 38904 32128 38956
rect 32180 38944 32186 38956
rect 32493 38947 32551 38953
rect 32493 38944 32505 38947
rect 32180 38916 32505 38944
rect 32180 38904 32186 38916
rect 32493 38913 32505 38916
rect 32539 38913 32551 38947
rect 32493 38907 32551 38913
rect 32582 38904 32588 38956
rect 32640 38944 32646 38956
rect 32876 38953 32904 38984
rect 32861 38947 32919 38953
rect 32640 38916 32685 38944
rect 32640 38904 32646 38916
rect 32861 38913 32873 38947
rect 32907 38913 32919 38947
rect 32861 38907 32919 38913
rect 32953 38947 33011 38953
rect 32953 38913 32965 38947
rect 32999 38944 33011 38947
rect 33134 38944 33140 38956
rect 32999 38916 33140 38944
rect 32999 38913 33011 38916
rect 32953 38907 33011 38913
rect 33134 38904 33140 38916
rect 33192 38904 33198 38956
rect 30699 38848 31708 38876
rect 31864 38848 31984 38876
rect 30699 38845 30711 38848
rect 30653 38839 30711 38845
rect 31864 38808 31892 38848
rect 30484 38780 31892 38808
rect 30377 38771 30435 38777
rect 27672 38712 27936 38740
rect 27672 38700 27678 38712
rect 27982 38700 27988 38752
rect 28040 38740 28046 38752
rect 28626 38740 28632 38752
rect 28040 38712 28632 38740
rect 28040 38700 28046 38712
rect 28626 38700 28632 38712
rect 28684 38700 28690 38752
rect 29454 38740 29460 38752
rect 29415 38712 29460 38740
rect 29454 38700 29460 38712
rect 29512 38700 29518 38752
rect 29638 38700 29644 38752
rect 29696 38740 29702 38752
rect 30006 38740 30012 38752
rect 29696 38712 30012 38740
rect 29696 38700 29702 38712
rect 30006 38700 30012 38712
rect 30064 38700 30070 38752
rect 30392 38740 30420 38771
rect 31938 38768 31944 38820
rect 31996 38808 32002 38820
rect 33244 38808 33272 38984
rect 36354 38972 36360 38984
rect 36412 38972 36418 39024
rect 34149 38947 34207 38953
rect 34149 38913 34161 38947
rect 34195 38944 34207 38947
rect 34514 38944 34520 38956
rect 34195 38916 34520 38944
rect 34195 38913 34207 38916
rect 34149 38907 34207 38913
rect 34514 38904 34520 38916
rect 34572 38904 34578 38956
rect 34790 38904 34796 38956
rect 34848 38944 34854 38956
rect 35253 38947 35311 38953
rect 35253 38944 35265 38947
rect 34848 38916 35265 38944
rect 34848 38904 34854 38916
rect 35253 38913 35265 38916
rect 35299 38913 35311 38947
rect 35253 38907 35311 38913
rect 33594 38836 33600 38888
rect 33652 38876 33658 38888
rect 34054 38876 34060 38888
rect 33652 38848 34060 38876
rect 33652 38836 33658 38848
rect 34054 38836 34060 38848
rect 34112 38836 34118 38888
rect 34238 38876 34244 38888
rect 34151 38848 34244 38876
rect 34238 38836 34244 38848
rect 34296 38836 34302 38888
rect 34330 38836 34336 38888
rect 34388 38876 34394 38888
rect 34388 38848 34433 38876
rect 34388 38836 34394 38848
rect 34606 38836 34612 38888
rect 34664 38876 34670 38888
rect 35066 38876 35072 38888
rect 34664 38848 35072 38876
rect 34664 38836 34670 38848
rect 35066 38836 35072 38848
rect 35124 38836 35130 38888
rect 35161 38879 35219 38885
rect 35161 38845 35173 38879
rect 35207 38876 35219 38879
rect 35342 38876 35348 38888
rect 35207 38848 35348 38876
rect 35207 38845 35219 38848
rect 35161 38839 35219 38845
rect 31996 38780 33272 38808
rect 34256 38808 34284 38836
rect 34256 38780 34376 38808
rect 31996 38768 32002 38780
rect 30650 38740 30656 38752
rect 30392 38712 30656 38740
rect 30650 38700 30656 38712
rect 30708 38700 30714 38752
rect 31110 38740 31116 38752
rect 31071 38712 31116 38740
rect 31110 38700 31116 38712
rect 31168 38700 31174 38752
rect 34348 38740 34376 38780
rect 34422 38768 34428 38820
rect 34480 38808 34486 38820
rect 35176 38808 35204 38839
rect 35342 38836 35348 38848
rect 35400 38836 35406 38888
rect 34480 38780 35204 38808
rect 34480 38768 34486 38780
rect 34514 38740 34520 38752
rect 34348 38712 34520 38740
rect 34514 38700 34520 38712
rect 34572 38700 34578 38752
rect 34698 38700 34704 38752
rect 34756 38740 34762 38752
rect 34885 38743 34943 38749
rect 34885 38740 34897 38743
rect 34756 38712 34897 38740
rect 34756 38700 34762 38712
rect 34885 38709 34897 38712
rect 34931 38709 34943 38743
rect 35066 38740 35072 38752
rect 35027 38712 35072 38740
rect 34885 38703 34943 38709
rect 35066 38700 35072 38712
rect 35124 38700 35130 38752
rect 35805 38743 35863 38749
rect 35805 38709 35817 38743
rect 35851 38740 35863 38743
rect 36170 38740 36176 38752
rect 35851 38712 36176 38740
rect 35851 38709 35863 38712
rect 35805 38703 35863 38709
rect 36170 38700 36176 38712
rect 36228 38700 36234 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 17126 38536 17132 38548
rect 16316 38508 17132 38536
rect 16316 38400 16344 38508
rect 17126 38496 17132 38508
rect 17184 38496 17190 38548
rect 17773 38539 17831 38545
rect 17773 38505 17785 38539
rect 17819 38536 17831 38539
rect 18325 38539 18383 38545
rect 18325 38536 18337 38539
rect 17819 38508 18337 38536
rect 17819 38505 17831 38508
rect 17773 38499 17831 38505
rect 18325 38505 18337 38508
rect 18371 38505 18383 38539
rect 18506 38536 18512 38548
rect 18467 38508 18512 38536
rect 18325 38499 18383 38505
rect 18506 38496 18512 38508
rect 18564 38496 18570 38548
rect 18598 38496 18604 38548
rect 18656 38536 18662 38548
rect 18656 38508 20760 38536
rect 18656 38496 18662 38508
rect 17862 38428 17868 38480
rect 17920 38468 17926 38480
rect 20732 38468 20760 38508
rect 20806 38496 20812 38548
rect 20864 38536 20870 38548
rect 22005 38539 22063 38545
rect 22005 38536 22017 38539
rect 20864 38508 22017 38536
rect 20864 38496 20870 38508
rect 22005 38505 22017 38508
rect 22051 38505 22063 38539
rect 22005 38499 22063 38505
rect 22738 38496 22744 38548
rect 22796 38536 22802 38548
rect 28629 38539 28687 38545
rect 28629 38536 28641 38539
rect 22796 38508 28641 38536
rect 22796 38496 22802 38508
rect 28629 38505 28641 38508
rect 28675 38505 28687 38539
rect 28629 38499 28687 38505
rect 28828 38508 29500 38536
rect 17920 38440 20668 38468
rect 20732 38440 24072 38468
rect 17920 38428 17926 38440
rect 16393 38403 16451 38409
rect 16393 38400 16405 38403
rect 16316 38372 16405 38400
rect 16393 38369 16405 38372
rect 16439 38369 16451 38403
rect 16574 38400 16580 38412
rect 16535 38372 16580 38400
rect 16393 38363 16451 38369
rect 16574 38360 16580 38372
rect 16632 38360 16638 38412
rect 19242 38360 19248 38412
rect 19300 38400 19306 38412
rect 19300 38372 19932 38400
rect 19300 38360 19306 38372
rect 16301 38335 16359 38341
rect 16301 38301 16313 38335
rect 16347 38301 16359 38335
rect 16301 38295 16359 38301
rect 16485 38335 16543 38341
rect 16485 38301 16497 38335
rect 16531 38332 16543 38335
rect 17218 38332 17224 38344
rect 16531 38304 17224 38332
rect 16531 38301 16543 38304
rect 16485 38295 16543 38301
rect 16316 38264 16344 38295
rect 17218 38292 17224 38304
rect 17276 38292 17282 38344
rect 17589 38335 17647 38341
rect 17589 38301 17601 38335
rect 17635 38332 17647 38335
rect 17678 38332 17684 38344
rect 17635 38304 17684 38332
rect 17635 38301 17647 38304
rect 17589 38295 17647 38301
rect 17678 38292 17684 38304
rect 17736 38292 17742 38344
rect 17862 38332 17868 38344
rect 17823 38304 17868 38332
rect 17862 38292 17868 38304
rect 17920 38292 17926 38344
rect 19904 38341 19932 38372
rect 19978 38360 19984 38412
rect 20036 38400 20042 38412
rect 20640 38400 20668 38440
rect 20036 38372 20081 38400
rect 20640 38372 20944 38400
rect 20036 38360 20042 38372
rect 19429 38335 19487 38341
rect 19429 38301 19441 38335
rect 19475 38301 19487 38335
rect 19429 38295 19487 38301
rect 19889 38335 19947 38341
rect 19889 38301 19901 38335
rect 19935 38301 19947 38335
rect 20530 38332 20536 38344
rect 20491 38304 20536 38332
rect 19889 38295 19947 38301
rect 17034 38264 17040 38276
rect 16316 38236 17040 38264
rect 17034 38224 17040 38236
rect 17092 38224 17098 38276
rect 18690 38264 18696 38276
rect 18651 38236 18696 38264
rect 18690 38224 18696 38236
rect 18748 38264 18754 38276
rect 19444 38264 19472 38295
rect 20530 38292 20536 38304
rect 20588 38292 20594 38344
rect 20916 38341 20944 38372
rect 20901 38335 20959 38341
rect 20901 38301 20913 38335
rect 20947 38332 20959 38335
rect 21174 38332 21180 38344
rect 20947 38304 21180 38332
rect 20947 38301 20959 38304
rect 20901 38295 20959 38301
rect 21174 38292 21180 38304
rect 21232 38292 21238 38344
rect 21361 38335 21419 38341
rect 21361 38301 21373 38335
rect 21407 38332 21419 38335
rect 21468 38332 21496 38440
rect 21542 38360 21548 38412
rect 21600 38360 21606 38412
rect 21913 38403 21971 38409
rect 21913 38369 21925 38403
rect 21959 38400 21971 38403
rect 22462 38400 22468 38412
rect 21959 38372 22468 38400
rect 21959 38369 21971 38372
rect 21913 38363 21971 38369
rect 22462 38360 22468 38372
rect 22520 38360 22526 38412
rect 23106 38400 23112 38412
rect 22756 38372 23112 38400
rect 21407 38304 21496 38332
rect 21560 38332 21588 38360
rect 21821 38335 21879 38341
rect 21821 38332 21833 38335
rect 21560 38304 21833 38332
rect 21407 38301 21419 38304
rect 21361 38295 21419 38301
rect 21821 38301 21833 38304
rect 21867 38301 21879 38335
rect 22143 38335 22201 38341
rect 22143 38332 22155 38335
rect 21821 38295 21879 38301
rect 22066 38304 22155 38332
rect 18748 38236 19472 38264
rect 18748 38224 18754 38236
rect 16117 38199 16175 38205
rect 16117 38165 16129 38199
rect 16163 38196 16175 38199
rect 16298 38196 16304 38208
rect 16163 38168 16304 38196
rect 16163 38165 16175 38168
rect 16117 38159 16175 38165
rect 16298 38156 16304 38168
rect 16356 38156 16362 38208
rect 16390 38156 16396 38208
rect 16448 38196 16454 38208
rect 17313 38199 17371 38205
rect 17313 38196 17325 38199
rect 16448 38168 17325 38196
rect 16448 38156 16454 38168
rect 17313 38165 17325 38168
rect 17359 38165 17371 38199
rect 17313 38159 17371 38165
rect 17770 38156 17776 38208
rect 17828 38196 17834 38208
rect 18493 38199 18551 38205
rect 18493 38196 18505 38199
rect 17828 38168 18505 38196
rect 17828 38156 17834 38168
rect 18493 38165 18505 38168
rect 18539 38196 18551 38199
rect 20530 38196 20536 38208
rect 18539 38168 20536 38196
rect 18539 38165 18551 38168
rect 18493 38159 18551 38165
rect 20530 38156 20536 38168
rect 20588 38156 20594 38208
rect 21910 38156 21916 38208
rect 21968 38196 21974 38208
rect 22066 38196 22094 38304
rect 22143 38301 22155 38304
rect 22189 38301 22201 38335
rect 22143 38295 22201 38301
rect 22278 38292 22284 38344
rect 22336 38332 22342 38344
rect 22756 38341 22784 38372
rect 23106 38360 23112 38372
rect 23164 38360 23170 38412
rect 24044 38400 24072 38440
rect 24118 38428 24124 38480
rect 24176 38468 24182 38480
rect 24857 38471 24915 38477
rect 24857 38468 24869 38471
rect 24176 38440 24869 38468
rect 24176 38428 24182 38440
rect 24857 38437 24869 38440
rect 24903 38437 24915 38471
rect 24857 38431 24915 38437
rect 25130 38428 25136 38480
rect 25188 38468 25194 38480
rect 25958 38468 25964 38480
rect 25188 38440 25964 38468
rect 25188 38428 25194 38440
rect 25958 38428 25964 38440
rect 26016 38468 26022 38480
rect 26016 38440 27292 38468
rect 26016 38428 26022 38440
rect 26145 38403 26203 38409
rect 26145 38400 26157 38403
rect 24044 38372 26157 38400
rect 26145 38369 26157 38372
rect 26191 38369 26203 38403
rect 26145 38363 26203 38369
rect 26234 38360 26240 38412
rect 26292 38400 26298 38412
rect 26602 38400 26608 38412
rect 26292 38372 26608 38400
rect 26292 38360 26298 38372
rect 26602 38360 26608 38372
rect 26660 38360 26666 38412
rect 26789 38403 26847 38409
rect 26789 38369 26801 38403
rect 26835 38400 26847 38403
rect 27062 38400 27068 38412
rect 26835 38372 27068 38400
rect 26835 38369 26847 38372
rect 26789 38363 26847 38369
rect 22741 38335 22799 38341
rect 22336 38304 22429 38332
rect 22336 38292 22342 38304
rect 22741 38301 22753 38335
rect 22787 38301 22799 38335
rect 22741 38295 22799 38301
rect 22925 38335 22983 38341
rect 22925 38301 22937 38335
rect 22971 38332 22983 38335
rect 23566 38332 23572 38344
rect 22971 38304 23572 38332
rect 22971 38301 22983 38304
rect 22925 38295 22983 38301
rect 23566 38292 23572 38304
rect 23624 38292 23630 38344
rect 23661 38335 23719 38341
rect 23661 38301 23673 38335
rect 23707 38332 23719 38335
rect 24578 38332 24584 38344
rect 23707 38304 24584 38332
rect 23707 38301 23719 38304
rect 23661 38295 23719 38301
rect 24578 38292 24584 38304
rect 24636 38292 24642 38344
rect 26050 38332 26056 38344
rect 26011 38304 26056 38332
rect 26050 38292 26056 38304
rect 26108 38292 26114 38344
rect 22296 38264 22324 38292
rect 23290 38264 23296 38276
rect 22296 38236 23296 38264
rect 23290 38224 23296 38236
rect 23348 38224 23354 38276
rect 23845 38267 23903 38273
rect 23845 38233 23857 38267
rect 23891 38264 23903 38267
rect 26252 38264 26280 38360
rect 26326 38292 26332 38344
rect 26384 38332 26390 38344
rect 26804 38332 26832 38363
rect 27062 38360 27068 38372
rect 27120 38360 27126 38412
rect 27264 38409 27292 38440
rect 27890 38428 27896 38480
rect 27948 38468 27954 38480
rect 28828 38468 28856 38508
rect 27948 38440 28856 38468
rect 27948 38428 27954 38440
rect 28902 38428 28908 38480
rect 28960 38468 28966 38480
rect 28960 38440 29224 38468
rect 28960 38428 28966 38440
rect 27249 38403 27307 38409
rect 27249 38369 27261 38403
rect 27295 38369 27307 38403
rect 27249 38363 27307 38369
rect 28718 38360 28724 38412
rect 28776 38400 28782 38412
rect 28776 38372 28948 38400
rect 28776 38360 28782 38372
rect 26384 38304 26832 38332
rect 26973 38335 27031 38341
rect 26384 38292 26390 38304
rect 26973 38301 26985 38335
rect 27019 38332 27031 38335
rect 27430 38332 27436 38344
rect 27019 38304 27313 38332
rect 27391 38304 27436 38332
rect 27019 38301 27031 38304
rect 26973 38295 27031 38301
rect 23891 38236 26280 38264
rect 23891 38233 23903 38236
rect 23845 38227 23903 38233
rect 21968 38168 22094 38196
rect 21968 38156 21974 38168
rect 22646 38156 22652 38208
rect 22704 38196 22710 38208
rect 22741 38199 22799 38205
rect 22741 38196 22753 38199
rect 22704 38168 22753 38196
rect 22704 38156 22710 38168
rect 22741 38165 22753 38168
rect 22787 38165 22799 38199
rect 22741 38159 22799 38165
rect 22922 38156 22928 38208
rect 22980 38196 22986 38208
rect 23106 38196 23112 38208
rect 22980 38168 23112 38196
rect 22980 38156 22986 38168
rect 23106 38156 23112 38168
rect 23164 38196 23170 38208
rect 23860 38196 23888 38227
rect 24026 38196 24032 38208
rect 23164 38168 23888 38196
rect 23987 38168 24032 38196
rect 23164 38156 23170 38168
rect 24026 38156 24032 38168
rect 24084 38156 24090 38208
rect 25041 38199 25099 38205
rect 25041 38165 25053 38199
rect 25087 38196 25099 38199
rect 25130 38196 25136 38208
rect 25087 38168 25136 38196
rect 25087 38165 25099 38168
rect 25041 38159 25099 38165
rect 25130 38156 25136 38168
rect 25188 38156 25194 38208
rect 25590 38196 25596 38208
rect 25503 38168 25596 38196
rect 25590 38156 25596 38168
rect 25648 38196 25654 38208
rect 26142 38196 26148 38208
rect 25648 38168 26148 38196
rect 25648 38156 25654 38168
rect 26142 38156 26148 38168
rect 26200 38156 26206 38208
rect 27285 38196 27313 38304
rect 27430 38292 27436 38304
rect 27488 38292 27494 38344
rect 28920 38341 28948 38372
rect 28813 38335 28871 38341
rect 28813 38301 28825 38335
rect 28859 38301 28871 38335
rect 28813 38295 28871 38301
rect 28905 38335 28963 38341
rect 28905 38301 28917 38335
rect 28951 38301 28963 38335
rect 29086 38332 29092 38344
rect 29047 38304 29092 38332
rect 28905 38295 28963 38301
rect 28828 38264 28856 38295
rect 29086 38292 29092 38304
rect 29144 38292 29150 38344
rect 29196 38341 29224 38440
rect 29472 38400 29500 38508
rect 30558 38496 30564 38548
rect 30616 38536 30622 38548
rect 30745 38539 30803 38545
rect 30745 38536 30757 38539
rect 30616 38508 30757 38536
rect 30616 38496 30622 38508
rect 30745 38505 30757 38508
rect 30791 38505 30803 38539
rect 32582 38536 32588 38548
rect 30745 38499 30803 38505
rect 31726 38508 32588 38536
rect 30190 38428 30196 38480
rect 30248 38468 30254 38480
rect 30285 38471 30343 38477
rect 30285 38468 30297 38471
rect 30248 38440 30297 38468
rect 30248 38428 30254 38440
rect 30285 38437 30297 38440
rect 30331 38437 30343 38471
rect 30285 38431 30343 38437
rect 30561 38403 30619 38409
rect 30561 38400 30573 38403
rect 29472 38372 30573 38400
rect 30561 38369 30573 38372
rect 30607 38400 30619 38403
rect 31726 38400 31754 38508
rect 32582 38496 32588 38508
rect 32640 38496 32646 38548
rect 34606 38536 34612 38548
rect 33060 38508 34612 38536
rect 32858 38428 32864 38480
rect 32916 38468 32922 38480
rect 32953 38471 33011 38477
rect 32953 38468 32965 38471
rect 32916 38440 32965 38468
rect 32916 38428 32922 38440
rect 32953 38437 32965 38440
rect 32999 38437 33011 38471
rect 32953 38431 33011 38437
rect 32306 38400 32312 38412
rect 30607 38372 31754 38400
rect 32267 38372 32312 38400
rect 30607 38369 30619 38372
rect 30561 38363 30619 38369
rect 32306 38360 32312 38372
rect 32364 38360 32370 38412
rect 32582 38360 32588 38412
rect 32640 38400 32646 38412
rect 33060 38400 33088 38508
rect 34606 38496 34612 38508
rect 34664 38496 34670 38548
rect 33229 38403 33287 38409
rect 33229 38400 33241 38403
rect 32640 38372 33241 38400
rect 32640 38360 32646 38372
rect 33229 38369 33241 38372
rect 33275 38369 33287 38403
rect 33229 38363 33287 38369
rect 33318 38360 33324 38412
rect 33376 38409 33382 38412
rect 33376 38403 33404 38409
rect 33392 38369 33404 38403
rect 33502 38400 33508 38412
rect 33463 38372 33508 38400
rect 33376 38363 33404 38369
rect 33376 38360 33382 38363
rect 33502 38360 33508 38372
rect 33560 38360 33566 38412
rect 35161 38403 35219 38409
rect 35161 38369 35173 38403
rect 35207 38400 35219 38403
rect 35434 38400 35440 38412
rect 35207 38372 35440 38400
rect 35207 38369 35219 38372
rect 35161 38363 35219 38369
rect 35434 38360 35440 38372
rect 35492 38360 35498 38412
rect 29181 38335 29239 38341
rect 29181 38301 29193 38335
rect 29227 38301 29239 38335
rect 30374 38332 30380 38344
rect 30335 38304 30380 38332
rect 29181 38295 29239 38301
rect 30374 38292 30380 38304
rect 30432 38332 30438 38344
rect 30742 38332 30748 38344
rect 30432 38304 30748 38332
rect 30432 38292 30438 38304
rect 30742 38292 30748 38304
rect 30800 38292 30806 38344
rect 30837 38335 30895 38341
rect 30837 38301 30849 38335
rect 30883 38332 30895 38335
rect 31294 38332 31300 38344
rect 30883 38304 31300 38332
rect 30883 38301 30895 38304
rect 30837 38295 30895 38301
rect 28994 38264 29000 38276
rect 28828 38236 29000 38264
rect 28994 38224 29000 38236
rect 29052 38224 29058 38276
rect 29454 38224 29460 38276
rect 29512 38264 29518 38276
rect 30852 38264 30880 38295
rect 31294 38292 31300 38304
rect 31352 38332 31358 38344
rect 31938 38332 31944 38344
rect 31352 38304 31944 38332
rect 31352 38292 31358 38304
rect 31938 38292 31944 38304
rect 31996 38292 32002 38344
rect 32490 38332 32496 38344
rect 32451 38304 32496 38332
rect 32490 38292 32496 38304
rect 32548 38292 32554 38344
rect 29512 38236 30880 38264
rect 29512 38224 29518 38236
rect 35342 38224 35348 38276
rect 35400 38264 35406 38276
rect 35437 38267 35495 38273
rect 35437 38264 35449 38267
rect 35400 38236 35449 38264
rect 35400 38224 35406 38236
rect 35437 38233 35449 38236
rect 35483 38233 35495 38267
rect 35437 38227 35495 38233
rect 36170 38224 36176 38276
rect 36228 38224 36234 38276
rect 37090 38224 37096 38276
rect 37148 38264 37154 38276
rect 37185 38267 37243 38273
rect 37185 38264 37197 38267
rect 37148 38236 37197 38264
rect 37148 38224 37154 38236
rect 37185 38233 37197 38236
rect 37231 38233 37243 38267
rect 37185 38227 37243 38233
rect 28810 38196 28816 38208
rect 27285 38168 28816 38196
rect 28810 38156 28816 38168
rect 28868 38156 28874 38208
rect 29730 38196 29736 38208
rect 29691 38168 29736 38196
rect 29730 38156 29736 38168
rect 29788 38156 29794 38208
rect 30006 38156 30012 38208
rect 30064 38196 30070 38208
rect 30469 38199 30527 38205
rect 30469 38196 30481 38199
rect 30064 38168 30481 38196
rect 30064 38156 30070 38168
rect 30469 38165 30481 38168
rect 30515 38196 30527 38199
rect 31202 38196 31208 38208
rect 30515 38168 31208 38196
rect 30515 38165 30527 38168
rect 30469 38159 30527 38165
rect 31202 38156 31208 38168
rect 31260 38196 31266 38208
rect 31297 38199 31355 38205
rect 31297 38196 31309 38199
rect 31260 38168 31309 38196
rect 31260 38156 31266 38168
rect 31297 38165 31309 38168
rect 31343 38165 31355 38199
rect 34146 38196 34152 38208
rect 34107 38168 34152 38196
rect 31297 38159 31355 38165
rect 34146 38156 34152 38168
rect 34204 38156 34210 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 17218 37952 17224 38004
rect 17276 37992 17282 38004
rect 17865 37995 17923 38001
rect 17865 37992 17877 37995
rect 17276 37964 17877 37992
rect 17276 37952 17282 37964
rect 17865 37961 17877 37964
rect 17911 37992 17923 37995
rect 18690 37992 18696 38004
rect 17911 37964 18696 37992
rect 17911 37961 17923 37964
rect 17865 37955 17923 37961
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 19613 37995 19671 38001
rect 19613 37961 19625 37995
rect 19659 37992 19671 37995
rect 20714 37992 20720 38004
rect 19659 37964 20720 37992
rect 19659 37961 19671 37964
rect 19613 37955 19671 37961
rect 20714 37952 20720 37964
rect 20772 37952 20778 38004
rect 21082 37952 21088 38004
rect 21140 37992 21146 38004
rect 21361 37995 21419 38001
rect 21361 37992 21373 37995
rect 21140 37964 21373 37992
rect 21140 37952 21146 37964
rect 21361 37961 21373 37964
rect 21407 37961 21419 37995
rect 21361 37955 21419 37961
rect 22940 37964 23428 37992
rect 17681 37927 17739 37933
rect 17681 37893 17693 37927
rect 17727 37924 17739 37927
rect 17770 37924 17776 37936
rect 17727 37896 17776 37924
rect 17727 37893 17739 37896
rect 17681 37887 17739 37893
rect 17770 37884 17776 37896
rect 17828 37884 17834 37936
rect 22094 37924 22100 37936
rect 20456 37896 22100 37924
rect 15473 37859 15531 37865
rect 15473 37825 15485 37859
rect 15519 37856 15531 37859
rect 15562 37856 15568 37868
rect 15519 37828 15568 37856
rect 15519 37825 15531 37828
rect 15473 37819 15531 37825
rect 15562 37816 15568 37828
rect 15620 37816 15626 37868
rect 15657 37859 15715 37865
rect 15657 37825 15669 37859
rect 15703 37856 15715 37859
rect 16574 37856 16580 37868
rect 15703 37828 16580 37856
rect 15703 37825 15715 37828
rect 15657 37819 15715 37825
rect 16574 37816 16580 37828
rect 16632 37816 16638 37868
rect 17954 37816 17960 37868
rect 18012 37856 18018 37868
rect 18785 37859 18843 37865
rect 18012 37828 18057 37856
rect 18012 37816 18018 37828
rect 18785 37825 18797 37859
rect 18831 37856 18843 37859
rect 18874 37856 18880 37868
rect 18831 37828 18880 37856
rect 18831 37825 18843 37828
rect 18785 37819 18843 37825
rect 18874 37816 18880 37828
rect 18932 37816 18938 37868
rect 19794 37856 19800 37868
rect 19755 37828 19800 37856
rect 19794 37816 19800 37828
rect 19852 37816 19858 37868
rect 20456 37865 20484 37896
rect 22094 37884 22100 37896
rect 22152 37884 22158 37936
rect 22940 37924 22968 37964
rect 23400 37933 23428 37964
rect 23474 37952 23480 38004
rect 23532 37992 23538 38004
rect 28537 37995 28595 38001
rect 28537 37992 28549 37995
rect 23532 37964 28549 37992
rect 23532 37952 23538 37964
rect 28537 37961 28549 37964
rect 28583 37961 28595 37995
rect 31478 37992 31484 38004
rect 28537 37955 28595 37961
rect 28736 37964 31484 37992
rect 23169 37927 23227 37933
rect 23169 37924 23181 37927
rect 22204 37896 22968 37924
rect 23032 37896 23181 37924
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37825 20039 37859
rect 19981 37819 20039 37825
rect 20441 37859 20499 37865
rect 20441 37825 20453 37859
rect 20487 37825 20499 37859
rect 20441 37819 20499 37825
rect 20717 37859 20775 37865
rect 20717 37825 20729 37859
rect 20763 37856 20775 37859
rect 20898 37856 20904 37868
rect 20763 37828 20904 37856
rect 20763 37825 20775 37828
rect 20717 37819 20775 37825
rect 19996 37788 20024 37819
rect 20898 37816 20904 37828
rect 20956 37816 20962 37868
rect 21266 37816 21272 37868
rect 21324 37856 21330 37868
rect 22204 37865 22232 37896
rect 22189 37859 22247 37865
rect 22189 37856 22201 37859
rect 21324 37828 22201 37856
rect 21324 37816 21330 37828
rect 22189 37825 22201 37828
rect 22235 37825 22247 37859
rect 22189 37819 22247 37825
rect 22373 37859 22431 37865
rect 22373 37825 22385 37859
rect 22419 37856 22431 37859
rect 22554 37856 22560 37868
rect 22419 37828 22560 37856
rect 22419 37825 22431 37828
rect 22373 37819 22431 37825
rect 22554 37816 22560 37828
rect 22612 37856 22618 37868
rect 23032 37856 23060 37896
rect 23169 37893 23181 37896
rect 23215 37893 23227 37927
rect 23169 37887 23227 37893
rect 23385 37927 23443 37933
rect 23385 37893 23397 37927
rect 23431 37893 23443 37927
rect 23385 37887 23443 37893
rect 24026 37884 24032 37936
rect 24084 37924 24090 37936
rect 25406 37924 25412 37936
rect 24084 37896 25412 37924
rect 24084 37884 24090 37896
rect 25406 37884 25412 37896
rect 25464 37924 25470 37936
rect 26142 37924 26148 37936
rect 25464 37896 25682 37924
rect 26103 37896 26148 37924
rect 25464 37884 25470 37896
rect 22612 37828 23060 37856
rect 22612 37816 22618 37828
rect 23750 37816 23756 37868
rect 23808 37856 23814 37868
rect 23845 37859 23903 37865
rect 23845 37856 23857 37859
rect 23808 37828 23857 37856
rect 23808 37816 23814 37828
rect 23845 37825 23857 37828
rect 23891 37825 23903 37859
rect 23845 37819 23903 37825
rect 24486 37816 24492 37868
rect 24544 37856 24550 37868
rect 24581 37859 24639 37865
rect 24581 37856 24593 37859
rect 24544 37828 24593 37856
rect 24544 37816 24550 37828
rect 24581 37825 24593 37828
rect 24627 37825 24639 37859
rect 24581 37819 24639 37825
rect 24670 37816 24676 37868
rect 24728 37856 24734 37868
rect 25654 37865 25682 37896
rect 26142 37884 26148 37896
rect 26200 37884 26206 37936
rect 27798 37924 27804 37936
rect 27448 37896 27804 37924
rect 24765 37859 24823 37865
rect 24765 37856 24777 37859
rect 24728 37828 24777 37856
rect 24728 37816 24734 37828
rect 24765 37825 24777 37828
rect 24811 37825 24823 37859
rect 24765 37819 24823 37825
rect 25639 37859 25697 37865
rect 25639 37825 25651 37859
rect 25685 37825 25697 37859
rect 25639 37819 25697 37825
rect 25777 37859 25835 37865
rect 25777 37825 25789 37859
rect 25823 37856 25835 37859
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 25823 37828 27169 37856
rect 25823 37825 25835 37828
rect 25777 37819 25835 37825
rect 27157 37825 27169 37828
rect 27203 37825 27215 37859
rect 27157 37819 27215 37825
rect 27246 37816 27252 37868
rect 27304 37856 27310 37868
rect 27448 37865 27476 37896
rect 27798 37884 27804 37896
rect 27856 37924 27862 37936
rect 28258 37924 28264 37936
rect 27856 37896 28264 37924
rect 27856 37884 27862 37896
rect 28258 37884 28264 37896
rect 28316 37884 28322 37936
rect 27341 37859 27399 37865
rect 27341 37856 27353 37859
rect 27304 37828 27353 37856
rect 27304 37816 27310 37828
rect 27341 37825 27353 37828
rect 27387 37825 27399 37859
rect 27341 37819 27399 37825
rect 27433 37859 27491 37865
rect 27433 37825 27445 37859
rect 27479 37825 27491 37859
rect 27709 37859 27767 37865
rect 27709 37856 27721 37859
rect 27433 37819 27491 37825
rect 27540 37828 27721 37856
rect 21726 37788 21732 37800
rect 19996 37760 21732 37788
rect 21726 37748 21732 37760
rect 21784 37788 21790 37800
rect 21910 37788 21916 37800
rect 21784 37760 21916 37788
rect 21784 37748 21790 37760
rect 21910 37748 21916 37760
rect 21968 37748 21974 37800
rect 22097 37791 22155 37797
rect 22097 37757 22109 37791
rect 22143 37757 22155 37791
rect 22097 37751 22155 37757
rect 22281 37791 22339 37797
rect 22281 37757 22293 37791
rect 22327 37788 22339 37791
rect 22646 37788 22652 37800
rect 22327 37760 22652 37788
rect 22327 37757 22339 37760
rect 22281 37751 22339 37757
rect 17678 37720 17684 37732
rect 17639 37692 17684 37720
rect 17678 37680 17684 37692
rect 17736 37680 17742 37732
rect 15473 37655 15531 37661
rect 15473 37621 15485 37655
rect 15519 37652 15531 37655
rect 16390 37652 16396 37664
rect 15519 37624 16396 37652
rect 15519 37621 15531 37624
rect 15473 37615 15531 37621
rect 16390 37612 16396 37624
rect 16448 37612 16454 37664
rect 17218 37652 17224 37664
rect 17179 37624 17224 37652
rect 17218 37612 17224 37624
rect 17276 37612 17282 37664
rect 22112 37652 22140 37751
rect 22646 37748 22652 37760
rect 22704 37748 22710 37800
rect 26053 37791 26111 37797
rect 26053 37757 26065 37791
rect 26099 37757 26111 37791
rect 26053 37751 26111 37757
rect 22664 37720 22692 37748
rect 22664 37692 23244 37720
rect 22278 37652 22284 37664
rect 22112 37624 22284 37652
rect 22278 37612 22284 37624
rect 22336 37612 22342 37664
rect 22554 37652 22560 37664
rect 22515 37624 22560 37652
rect 22554 37612 22560 37624
rect 22612 37612 22618 37664
rect 22646 37612 22652 37664
rect 22704 37652 22710 37664
rect 23216 37661 23244 37692
rect 23290 37680 23296 37732
rect 23348 37720 23354 37732
rect 23348 37692 25084 37720
rect 23348 37680 23354 37692
rect 25056 37664 25084 37692
rect 25222 37680 25228 37732
rect 25280 37720 25286 37732
rect 25501 37723 25559 37729
rect 25501 37720 25513 37723
rect 25280 37692 25513 37720
rect 25280 37680 25286 37692
rect 25501 37689 25513 37692
rect 25547 37689 25559 37723
rect 25501 37683 25559 37689
rect 25774 37680 25780 37732
rect 25832 37720 25838 37732
rect 26068 37720 26096 37751
rect 26142 37748 26148 37800
rect 26200 37788 26206 37800
rect 27540 37788 27568 37828
rect 27709 37825 27721 37828
rect 27755 37856 27767 37859
rect 27755 37828 28396 37856
rect 27755 37825 27767 37828
rect 27709 37819 27767 37825
rect 26200 37760 27568 37788
rect 27617 37791 27675 37797
rect 26200 37748 26206 37760
rect 27617 37757 27629 37791
rect 27663 37788 27675 37791
rect 27890 37788 27896 37800
rect 27663 37760 27896 37788
rect 27663 37757 27675 37760
rect 27617 37751 27675 37757
rect 27890 37748 27896 37760
rect 27948 37748 27954 37800
rect 28368 37788 28396 37828
rect 28442 37816 28448 37868
rect 28500 37856 28506 37868
rect 28626 37856 28632 37868
rect 28500 37828 28632 37856
rect 28500 37816 28506 37828
rect 28626 37816 28632 37828
rect 28684 37856 28690 37868
rect 28736 37865 28764 37964
rect 31478 37952 31484 37964
rect 31536 37952 31542 38004
rect 31938 37952 31944 38004
rect 31996 37992 32002 38004
rect 33229 37995 33287 38001
rect 33229 37992 33241 37995
rect 31996 37964 33241 37992
rect 31996 37952 32002 37964
rect 33229 37961 33241 37964
rect 33275 37961 33287 37995
rect 33229 37955 33287 37961
rect 34241 37995 34299 38001
rect 34241 37961 34253 37995
rect 34287 37992 34299 37995
rect 34330 37992 34336 38004
rect 34287 37964 34336 37992
rect 34287 37961 34299 37964
rect 34241 37955 34299 37961
rect 34330 37952 34336 37964
rect 34388 37952 34394 38004
rect 34698 37992 34704 38004
rect 34659 37964 34704 37992
rect 34698 37952 34704 37964
rect 34756 37952 34762 38004
rect 35342 37992 35348 38004
rect 35303 37964 35348 37992
rect 35342 37952 35348 37964
rect 35400 37952 35406 38004
rect 31662 37924 31668 37936
rect 28920 37896 31668 37924
rect 28920 37865 28948 37896
rect 31662 37884 31668 37896
rect 31720 37884 31726 37936
rect 28721 37859 28779 37865
rect 28721 37856 28733 37859
rect 28684 37828 28733 37856
rect 28684 37816 28690 37828
rect 28721 37825 28733 37828
rect 28767 37825 28779 37859
rect 28721 37819 28779 37825
rect 28905 37859 28963 37865
rect 28905 37825 28917 37859
rect 28951 37825 28963 37859
rect 28905 37819 28963 37825
rect 29270 37816 29276 37868
rect 29328 37856 29334 37868
rect 29549 37859 29607 37865
rect 29549 37856 29561 37859
rect 29328 37828 29561 37856
rect 29328 37816 29334 37828
rect 29549 37825 29561 37828
rect 29595 37825 29607 37859
rect 29549 37819 29607 37825
rect 29687 37859 29745 37865
rect 29687 37825 29699 37859
rect 29733 37856 29745 37859
rect 30466 37856 30472 37868
rect 29733 37828 30472 37856
rect 29733 37825 29745 37828
rect 29687 37819 29745 37825
rect 30466 37816 30472 37828
rect 30524 37856 30530 37868
rect 31386 37856 31392 37868
rect 30524 37828 31392 37856
rect 30524 37816 30530 37828
rect 31386 37816 31392 37828
rect 31444 37816 31450 37868
rect 32490 37816 32496 37868
rect 32548 37856 32554 37868
rect 33042 37856 33048 37868
rect 32548 37828 33048 37856
rect 32548 37816 32554 37828
rect 33042 37816 33048 37828
rect 33100 37856 33106 37868
rect 34057 37859 34115 37865
rect 33100 37828 34008 37856
rect 33100 37816 33106 37828
rect 29454 37788 29460 37800
rect 28368 37760 29460 37788
rect 29454 37748 29460 37760
rect 29512 37748 29518 37800
rect 29917 37791 29975 37797
rect 29917 37757 29929 37791
rect 29963 37757 29975 37791
rect 33778 37788 33784 37800
rect 29917 37751 29975 37757
rect 30392 37760 33784 37788
rect 25832 37692 26096 37720
rect 25832 37680 25838 37692
rect 28442 37680 28448 37732
rect 28500 37720 28506 37732
rect 28718 37720 28724 37732
rect 28500 37692 28724 37720
rect 28500 37680 28506 37692
rect 28718 37680 28724 37692
rect 28776 37680 28782 37732
rect 29822 37720 29828 37732
rect 29783 37692 29828 37720
rect 29822 37680 29828 37692
rect 29880 37680 29886 37732
rect 23017 37655 23075 37661
rect 23017 37652 23029 37655
rect 22704 37624 23029 37652
rect 22704 37612 22710 37624
rect 23017 37621 23029 37624
rect 23063 37621 23075 37655
rect 23017 37615 23075 37621
rect 23201 37655 23259 37661
rect 23201 37621 23213 37655
rect 23247 37621 23259 37655
rect 23201 37615 23259 37621
rect 23658 37612 23664 37664
rect 23716 37652 23722 37664
rect 24029 37655 24087 37661
rect 24029 37652 24041 37655
rect 23716 37624 24041 37652
rect 23716 37612 23722 37624
rect 24029 37621 24041 37624
rect 24075 37652 24087 37655
rect 24118 37652 24124 37664
rect 24075 37624 24124 37652
rect 24075 37621 24087 37624
rect 24029 37615 24087 37621
rect 24118 37612 24124 37624
rect 24176 37612 24182 37664
rect 24210 37612 24216 37664
rect 24268 37652 24274 37664
rect 24673 37655 24731 37661
rect 24673 37652 24685 37655
rect 24268 37624 24685 37652
rect 24268 37612 24274 37624
rect 24673 37621 24685 37624
rect 24719 37621 24731 37655
rect 24673 37615 24731 37621
rect 25038 37612 25044 37664
rect 25096 37652 25102 37664
rect 27798 37652 27804 37664
rect 25096 37624 27804 37652
rect 25096 37612 25102 37624
rect 27798 37612 27804 37624
rect 27856 37612 27862 37664
rect 28902 37652 28908 37664
rect 28863 37624 28908 37652
rect 28902 37612 28908 37624
rect 28960 37612 28966 37664
rect 29178 37612 29184 37664
rect 29236 37652 29242 37664
rect 29932 37652 29960 37751
rect 30392 37664 30420 37760
rect 33778 37748 33784 37760
rect 33836 37788 33842 37800
rect 33873 37791 33931 37797
rect 33873 37788 33885 37791
rect 33836 37760 33885 37788
rect 33836 37748 33842 37760
rect 33873 37757 33885 37760
rect 33919 37757 33931 37791
rect 33980 37788 34008 37828
rect 34057 37825 34069 37859
rect 34103 37856 34115 37859
rect 34698 37856 34704 37868
rect 34103 37828 34704 37856
rect 34103 37825 34115 37828
rect 34057 37819 34115 37825
rect 34698 37816 34704 37828
rect 34756 37856 34762 37868
rect 35161 37859 35219 37865
rect 35161 37856 35173 37859
rect 34756 37828 35173 37856
rect 34756 37816 34762 37828
rect 35161 37825 35173 37828
rect 35207 37825 35219 37859
rect 35161 37819 35219 37825
rect 35069 37791 35127 37797
rect 35069 37788 35081 37791
rect 33980 37760 35081 37788
rect 33873 37751 33931 37757
rect 35069 37757 35081 37760
rect 35115 37757 35127 37791
rect 35069 37751 35127 37757
rect 32122 37720 32128 37732
rect 31404 37692 32128 37720
rect 31404 37664 31432 37692
rect 32122 37680 32128 37692
rect 32180 37680 32186 37732
rect 33888 37720 33916 37751
rect 35805 37723 35863 37729
rect 35805 37720 35817 37723
rect 32232 37692 33732 37720
rect 33888 37692 35817 37720
rect 30374 37652 30380 37664
rect 29236 37624 29960 37652
rect 30335 37624 30380 37652
rect 29236 37612 29242 37624
rect 30374 37612 30380 37624
rect 30432 37612 30438 37664
rect 31021 37655 31079 37661
rect 31021 37621 31033 37655
rect 31067 37652 31079 37655
rect 31202 37652 31208 37664
rect 31067 37624 31208 37652
rect 31067 37621 31079 37624
rect 31021 37615 31079 37621
rect 31202 37612 31208 37624
rect 31260 37652 31266 37664
rect 31386 37652 31392 37664
rect 31260 37624 31392 37652
rect 31260 37612 31266 37624
rect 31386 37612 31392 37624
rect 31444 37612 31450 37664
rect 31478 37612 31484 37664
rect 31536 37652 31542 37664
rect 32030 37652 32036 37664
rect 31536 37624 32036 37652
rect 31536 37612 31542 37624
rect 32030 37612 32036 37624
rect 32088 37652 32094 37664
rect 32232 37652 32260 37692
rect 32088 37624 32260 37652
rect 32769 37655 32827 37661
rect 32088 37612 32094 37624
rect 32769 37621 32781 37655
rect 32815 37652 32827 37655
rect 33594 37652 33600 37664
rect 32815 37624 33600 37652
rect 32815 37621 32827 37624
rect 32769 37615 32827 37621
rect 33594 37612 33600 37624
rect 33652 37612 33658 37664
rect 33704 37652 33732 37692
rect 35805 37689 35817 37692
rect 35851 37689 35863 37723
rect 35805 37683 35863 37689
rect 35986 37652 35992 37664
rect 33704 37624 35992 37652
rect 35986 37612 35992 37624
rect 36044 37612 36050 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 18877 37451 18935 37457
rect 18877 37417 18889 37451
rect 18923 37448 18935 37451
rect 19794 37448 19800 37460
rect 18923 37420 19800 37448
rect 18923 37417 18935 37420
rect 18877 37411 18935 37417
rect 19794 37408 19800 37420
rect 19852 37448 19858 37460
rect 20990 37448 20996 37460
rect 19852 37420 20996 37448
rect 19852 37408 19858 37420
rect 20990 37408 20996 37420
rect 21048 37408 21054 37460
rect 21082 37408 21088 37460
rect 21140 37448 21146 37460
rect 23658 37448 23664 37460
rect 21140 37420 23664 37448
rect 21140 37408 21146 37420
rect 23658 37408 23664 37420
rect 23716 37408 23722 37460
rect 23842 37408 23848 37460
rect 23900 37448 23906 37460
rect 23900 37420 23993 37448
rect 23900 37408 23906 37420
rect 24118 37408 24124 37460
rect 24176 37448 24182 37460
rect 25498 37448 25504 37460
rect 24176 37420 25504 37448
rect 24176 37408 24182 37420
rect 25498 37408 25504 37420
rect 25556 37448 25562 37460
rect 25774 37448 25780 37460
rect 25556 37420 25780 37448
rect 25556 37408 25562 37420
rect 25774 37408 25780 37420
rect 25832 37448 25838 37460
rect 26142 37448 26148 37460
rect 25832 37420 26148 37448
rect 25832 37408 25838 37420
rect 26142 37408 26148 37420
rect 26200 37408 26206 37460
rect 26878 37408 26884 37460
rect 26936 37448 26942 37460
rect 28077 37451 28135 37457
rect 28077 37448 28089 37451
rect 26936 37420 28089 37448
rect 26936 37408 26942 37420
rect 28077 37417 28089 37420
rect 28123 37448 28135 37451
rect 28350 37448 28356 37460
rect 28123 37420 28356 37448
rect 28123 37417 28135 37420
rect 28077 37411 28135 37417
rect 28350 37408 28356 37420
rect 28408 37408 28414 37460
rect 30190 37408 30196 37460
rect 30248 37448 30254 37460
rect 30745 37451 30803 37457
rect 30248 37420 30512 37448
rect 30248 37408 30254 37420
rect 22094 37340 22100 37392
rect 22152 37380 22158 37392
rect 23106 37380 23112 37392
rect 22152 37352 23112 37380
rect 22152 37340 22158 37352
rect 23106 37340 23112 37352
rect 23164 37340 23170 37392
rect 23860 37380 23888 37408
rect 26234 37380 26240 37392
rect 23860 37352 26240 37380
rect 15749 37315 15807 37321
rect 15749 37281 15761 37315
rect 15795 37312 15807 37315
rect 16574 37312 16580 37324
rect 15795 37284 16580 37312
rect 15795 37281 15807 37284
rect 15749 37275 15807 37281
rect 16574 37272 16580 37284
rect 16632 37312 16638 37324
rect 17586 37312 17592 37324
rect 16632 37284 17592 37312
rect 16632 37272 16638 37284
rect 17586 37272 17592 37284
rect 17644 37272 17650 37324
rect 18325 37315 18383 37321
rect 18325 37281 18337 37315
rect 18371 37312 18383 37315
rect 18874 37312 18880 37324
rect 18371 37284 18880 37312
rect 18371 37281 18383 37284
rect 18325 37275 18383 37281
rect 18874 37272 18880 37284
rect 18932 37312 18938 37324
rect 21542 37312 21548 37324
rect 18932 37284 21548 37312
rect 18932 37272 18938 37284
rect 21542 37272 21548 37284
rect 21600 37272 21606 37324
rect 22186 37272 22192 37324
rect 22244 37312 22250 37324
rect 23382 37312 23388 37324
rect 22244 37284 22692 37312
rect 22244 37272 22250 37284
rect 15562 37244 15568 37256
rect 15523 37216 15568 37244
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 16209 37247 16267 37253
rect 16209 37213 16221 37247
rect 16255 37213 16267 37247
rect 16390 37244 16396 37256
rect 16351 37216 16396 37244
rect 16209 37207 16267 37213
rect 15378 37176 15384 37188
rect 15291 37148 15384 37176
rect 15378 37136 15384 37148
rect 15436 37176 15442 37188
rect 16224 37176 16252 37207
rect 16390 37204 16396 37216
rect 16448 37204 16454 37256
rect 17037 37247 17095 37253
rect 17037 37213 17049 37247
rect 17083 37244 17095 37247
rect 17126 37244 17132 37256
rect 17083 37216 17132 37244
rect 17083 37213 17095 37216
rect 17037 37207 17095 37213
rect 17126 37204 17132 37216
rect 17184 37204 17190 37256
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 17276 37216 17816 37244
rect 17276 37204 17282 37216
rect 15436 37148 16252 37176
rect 15436 37136 15442 37148
rect 17788 37120 17816 37216
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20625 37247 20683 37253
rect 20625 37244 20637 37247
rect 20220 37216 20637 37244
rect 20220 37204 20226 37216
rect 20625 37213 20637 37216
rect 20671 37213 20683 37247
rect 20625 37207 20683 37213
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 21358 37244 21364 37256
rect 20947 37216 21364 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 21358 37204 21364 37216
rect 21416 37244 21422 37256
rect 22002 37244 22008 37256
rect 21416 37216 22008 37244
rect 21416 37204 21422 37216
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 22278 37204 22284 37256
rect 22336 37244 22342 37256
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 22336 37216 22385 37244
rect 22336 37204 22342 37216
rect 22373 37213 22385 37216
rect 22419 37213 22431 37247
rect 22373 37207 22431 37213
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22520 37216 22565 37244
rect 22520 37204 22526 37216
rect 21726 37136 21732 37188
rect 21784 37176 21790 37188
rect 22664 37185 22692 37284
rect 22756 37284 23388 37312
rect 22756 37253 22784 37284
rect 23124 37256 23152 37284
rect 23382 37272 23388 37284
rect 23440 37272 23446 37324
rect 23750 37312 23756 37324
rect 23711 37284 23756 37312
rect 23750 37272 23756 37284
rect 23808 37272 23814 37324
rect 22741 37247 22799 37253
rect 22741 37213 22753 37247
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 22830 37204 22836 37256
rect 22888 37253 22894 37256
rect 22888 37244 22896 37253
rect 22888 37216 22933 37244
rect 22888 37207 22896 37216
rect 22888 37204 22894 37207
rect 23106 37204 23112 37256
rect 23164 37204 23170 37256
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37213 23719 37247
rect 24762 37244 24768 37256
rect 24723 37216 24768 37244
rect 23661 37207 23719 37213
rect 21913 37179 21971 37185
rect 21913 37176 21925 37179
rect 21784 37148 21925 37176
rect 21784 37136 21790 37148
rect 21913 37145 21925 37148
rect 21959 37176 21971 37179
rect 22649 37179 22707 37185
rect 21959 37148 22600 37176
rect 21959 37145 21971 37148
rect 21913 37139 21971 37145
rect 16482 37108 16488 37120
rect 16443 37080 16488 37108
rect 16482 37068 16488 37080
rect 16540 37068 16546 37120
rect 17221 37111 17279 37117
rect 17221 37077 17233 37111
rect 17267 37108 17279 37111
rect 17494 37108 17500 37120
rect 17267 37080 17500 37108
rect 17267 37077 17279 37080
rect 17221 37071 17279 37077
rect 17494 37068 17500 37080
rect 17552 37068 17558 37120
rect 17770 37108 17776 37120
rect 17731 37080 17776 37108
rect 17770 37068 17776 37080
rect 17828 37068 17834 37120
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19705 37111 19763 37117
rect 19705 37108 19717 37111
rect 19484 37080 19717 37108
rect 19484 37068 19490 37080
rect 19705 37077 19717 37080
rect 19751 37077 19763 37111
rect 19705 37071 19763 37077
rect 20441 37111 20499 37117
rect 20441 37077 20453 37111
rect 20487 37108 20499 37111
rect 20530 37108 20536 37120
rect 20487 37080 20536 37108
rect 20487 37077 20499 37080
rect 20441 37071 20499 37077
rect 20530 37068 20536 37080
rect 20588 37068 20594 37120
rect 20809 37111 20867 37117
rect 20809 37077 20821 37111
rect 20855 37108 20867 37111
rect 21542 37108 21548 37120
rect 20855 37080 21548 37108
rect 20855 37077 20867 37080
rect 20809 37071 20867 37077
rect 21542 37068 21548 37080
rect 21600 37068 21606 37120
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 22462 37108 22468 37120
rect 22152 37080 22468 37108
rect 22152 37068 22158 37080
rect 22462 37068 22468 37080
rect 22520 37068 22526 37120
rect 22572 37108 22600 37148
rect 22649 37145 22661 37179
rect 22695 37176 22707 37179
rect 23474 37176 23480 37188
rect 22695 37148 23480 37176
rect 22695 37145 22707 37148
rect 22649 37139 22707 37145
rect 23474 37136 23480 37148
rect 23532 37136 23538 37188
rect 23676 37176 23704 37207
rect 24762 37204 24768 37216
rect 24820 37204 24826 37256
rect 24872 37253 24900 37352
rect 26234 37340 26240 37352
rect 26292 37340 26298 37392
rect 27540 37352 27936 37380
rect 25317 37315 25375 37321
rect 25317 37281 25329 37315
rect 25363 37312 25375 37315
rect 27540 37312 27568 37352
rect 27798 37312 27804 37324
rect 25363 37284 27568 37312
rect 27632 37284 27804 37312
rect 25363 37281 25375 37284
rect 25317 37275 25375 37281
rect 24857 37247 24915 37253
rect 24857 37213 24869 37247
rect 24903 37213 24915 37247
rect 25038 37244 25044 37256
rect 24999 37216 25044 37244
rect 24857 37207 24915 37213
rect 25038 37204 25044 37216
rect 25096 37204 25102 37256
rect 25133 37247 25191 37253
rect 25133 37213 25145 37247
rect 25179 37213 25191 37247
rect 25133 37207 25191 37213
rect 25777 37247 25835 37253
rect 25777 37213 25789 37247
rect 25823 37213 25835 37247
rect 25958 37244 25964 37256
rect 25919 37216 25964 37244
rect 25777 37207 25835 37213
rect 24670 37176 24676 37188
rect 23676 37148 24676 37176
rect 24670 37136 24676 37148
rect 24728 37176 24734 37188
rect 25148 37176 25176 37207
rect 24728 37148 25176 37176
rect 25792 37176 25820 37207
rect 25958 37204 25964 37216
rect 26016 37204 26022 37256
rect 26234 37204 26240 37256
rect 26292 37244 26298 37256
rect 26513 37247 26571 37253
rect 26513 37244 26525 37247
rect 26292 37216 26525 37244
rect 26292 37204 26298 37216
rect 26513 37213 26525 37216
rect 26559 37213 26571 37247
rect 26513 37207 26571 37213
rect 26697 37247 26755 37253
rect 26697 37213 26709 37247
rect 26743 37244 26755 37247
rect 26786 37244 26792 37256
rect 26743 37216 26792 37244
rect 26743 37213 26755 37216
rect 26697 37207 26755 37213
rect 26786 37204 26792 37216
rect 26844 37204 26850 37256
rect 27632 37253 27660 37284
rect 27798 37272 27804 37284
rect 27856 37272 27862 37324
rect 27908 37312 27936 37352
rect 28902 37340 28908 37392
rect 28960 37380 28966 37392
rect 30282 37380 30288 37392
rect 28960 37352 30288 37380
rect 28960 37340 28966 37352
rect 30282 37340 30288 37352
rect 30340 37340 30346 37392
rect 30190 37312 30196 37324
rect 27908 37284 30196 37312
rect 30190 37272 30196 37284
rect 30248 37272 30254 37324
rect 30484 37312 30512 37420
rect 30745 37417 30757 37451
rect 30791 37448 30803 37451
rect 30926 37448 30932 37460
rect 30791 37420 30932 37448
rect 30791 37417 30803 37420
rect 30745 37411 30803 37417
rect 30926 37408 30932 37420
rect 30984 37448 30990 37460
rect 32582 37448 32588 37460
rect 30984 37420 32588 37448
rect 30984 37408 30990 37420
rect 32582 37408 32588 37420
rect 32640 37408 32646 37460
rect 33870 37408 33876 37460
rect 33928 37448 33934 37460
rect 33965 37451 34023 37457
rect 33965 37448 33977 37451
rect 33928 37420 33977 37448
rect 33928 37408 33934 37420
rect 33965 37417 33977 37420
rect 34011 37448 34023 37451
rect 34422 37448 34428 37460
rect 34011 37420 34428 37448
rect 34011 37417 34023 37420
rect 33965 37411 34023 37417
rect 34422 37408 34428 37420
rect 34480 37408 34486 37460
rect 31662 37380 31668 37392
rect 31623 37352 31668 37380
rect 31662 37340 31668 37352
rect 31720 37340 31726 37392
rect 33594 37340 33600 37392
rect 33652 37380 33658 37392
rect 35529 37383 35587 37389
rect 35529 37380 35541 37383
rect 33652 37352 35541 37380
rect 33652 37340 33658 37352
rect 35529 37349 35541 37352
rect 35575 37349 35587 37383
rect 35529 37343 35587 37349
rect 31849 37315 31907 37321
rect 31849 37312 31861 37315
rect 30484 37284 31861 37312
rect 31849 37281 31861 37284
rect 31895 37281 31907 37315
rect 33318 37312 33324 37324
rect 31849 37275 31907 37281
rect 32692 37284 33324 37312
rect 27617 37247 27675 37253
rect 27617 37213 27629 37247
rect 27663 37213 27675 37247
rect 27617 37207 27675 37213
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 27893 37247 27951 37253
rect 27764 37216 27809 37244
rect 27764 37204 27770 37216
rect 27893 37213 27905 37247
rect 27939 37244 27951 37247
rect 28258 37244 28264 37256
rect 27939 37216 28264 37244
rect 27939 37213 27951 37216
rect 27893 37207 27951 37213
rect 28258 37204 28264 37216
rect 28316 37204 28322 37256
rect 28442 37204 28448 37256
rect 28500 37244 28506 37256
rect 28537 37247 28595 37253
rect 28537 37244 28549 37247
rect 28500 37216 28549 37244
rect 28500 37204 28506 37216
rect 28537 37213 28549 37216
rect 28583 37213 28595 37247
rect 30837 37247 30895 37253
rect 28537 37207 28595 37213
rect 28644 37216 30236 37244
rect 26418 37176 26424 37188
rect 25792 37148 26424 37176
rect 24728 37136 24734 37148
rect 26418 37136 26424 37148
rect 26476 37136 26482 37188
rect 26605 37179 26663 37185
rect 26605 37145 26617 37179
rect 26651 37176 26663 37179
rect 27246 37176 27252 37188
rect 26651 37148 27252 37176
rect 26651 37145 26663 37148
rect 26605 37139 26663 37145
rect 27246 37136 27252 37148
rect 27304 37176 27310 37188
rect 28644 37176 28672 37216
rect 27304 37148 28672 37176
rect 28721 37179 28779 37185
rect 27304 37136 27310 37148
rect 28721 37145 28733 37179
rect 28767 37145 28779 37179
rect 28721 37139 28779 37145
rect 22830 37108 22836 37120
rect 22572 37080 22836 37108
rect 22830 37068 22836 37080
rect 22888 37068 22894 37120
rect 23017 37111 23075 37117
rect 23017 37077 23029 37111
rect 23063 37108 23075 37111
rect 23658 37108 23664 37120
rect 23063 37080 23664 37108
rect 23063 37077 23075 37080
rect 23017 37071 23075 37077
rect 23658 37068 23664 37080
rect 23716 37068 23722 37120
rect 24029 37111 24087 37117
rect 24029 37077 24041 37111
rect 24075 37108 24087 37111
rect 24118 37108 24124 37120
rect 24075 37080 24124 37108
rect 24075 37077 24087 37080
rect 24029 37071 24087 37077
rect 24118 37068 24124 37080
rect 24176 37068 24182 37120
rect 25866 37108 25872 37120
rect 25827 37080 25872 37108
rect 25866 37068 25872 37080
rect 25924 37068 25930 37120
rect 26786 37068 26792 37120
rect 26844 37108 26850 37120
rect 28736 37108 28764 37139
rect 28810 37136 28816 37188
rect 28868 37176 28874 37188
rect 28905 37179 28963 37185
rect 28905 37176 28917 37179
rect 28868 37148 28917 37176
rect 28868 37136 28874 37148
rect 28905 37145 28917 37148
rect 28951 37145 28963 37179
rect 30208 37176 30236 37216
rect 30837 37213 30849 37247
rect 30883 37244 30895 37247
rect 30926 37244 30932 37256
rect 30883 37216 30932 37244
rect 30883 37213 30895 37216
rect 30837 37207 30895 37213
rect 30926 37204 30932 37216
rect 30984 37204 30990 37256
rect 31573 37247 31631 37253
rect 31573 37213 31585 37247
rect 31619 37213 31631 37247
rect 31573 37207 31631 37213
rect 31018 37176 31024 37188
rect 30208 37148 31024 37176
rect 28905 37139 28963 37145
rect 30098 37108 30104 37120
rect 26844 37080 28764 37108
rect 30059 37080 30104 37108
rect 26844 37068 26850 37080
rect 30098 37068 30104 37080
rect 30156 37068 30162 37120
rect 30282 37068 30288 37120
rect 30340 37108 30346 37120
rect 30484 37117 30512 37148
rect 31018 37136 31024 37148
rect 31076 37136 31082 37188
rect 31588 37176 31616 37207
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32033 37247 32091 37253
rect 31812 37216 31857 37244
rect 31812 37204 31818 37216
rect 32033 37213 32045 37247
rect 32079 37244 32091 37247
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32079 37216 32505 37244
rect 32079 37213 32091 37216
rect 32033 37207 32091 37213
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 32582 37204 32588 37256
rect 32640 37244 32646 37256
rect 32692 37253 32720 37284
rect 33318 37272 33324 37284
rect 33376 37272 33382 37324
rect 32677 37247 32735 37253
rect 32677 37244 32689 37247
rect 32640 37216 32689 37244
rect 32640 37204 32646 37216
rect 32677 37213 32689 37216
rect 32723 37213 32735 37247
rect 32677 37207 32735 37213
rect 32861 37247 32919 37253
rect 32861 37213 32873 37247
rect 32907 37244 32919 37247
rect 33134 37244 33140 37256
rect 32907 37216 33140 37244
rect 32907 37213 32919 37216
rect 32861 37207 32919 37213
rect 33134 37204 33140 37216
rect 33192 37244 33198 37256
rect 33962 37244 33968 37256
rect 33192 37216 33968 37244
rect 33192 37204 33198 37216
rect 33962 37204 33968 37216
rect 34020 37204 34026 37256
rect 34054 37204 34060 37256
rect 34112 37244 34118 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34112 37216 34897 37244
rect 34112 37204 34118 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 35069 37247 35127 37253
rect 35069 37213 35081 37247
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 33502 37176 33508 37188
rect 31588 37148 33508 37176
rect 33502 37136 33508 37148
rect 33560 37136 33566 37188
rect 33781 37179 33839 37185
rect 33781 37145 33793 37179
rect 33827 37176 33839 37179
rect 33980 37176 34008 37204
rect 34330 37176 34336 37188
rect 33827 37148 34008 37176
rect 34164 37148 34336 37176
rect 33827 37145 33839 37148
rect 33781 37139 33839 37145
rect 30383 37111 30441 37117
rect 30383 37108 30395 37111
rect 30340 37080 30395 37108
rect 30340 37068 30346 37080
rect 30383 37077 30395 37080
rect 30429 37077 30441 37111
rect 30383 37071 30441 37077
rect 30469 37111 30527 37117
rect 30469 37077 30481 37111
rect 30515 37077 30527 37111
rect 30469 37071 30527 37077
rect 30561 37111 30619 37117
rect 30561 37077 30573 37111
rect 30607 37108 30619 37111
rect 30926 37108 30932 37120
rect 30607 37080 30932 37108
rect 30607 37077 30619 37080
rect 30561 37071 30619 37077
rect 30926 37068 30932 37080
rect 30984 37068 30990 37120
rect 31202 37068 31208 37120
rect 31260 37108 31266 37120
rect 31389 37111 31447 37117
rect 31389 37108 31401 37111
rect 31260 37080 31401 37108
rect 31260 37068 31266 37080
rect 31389 37077 31401 37080
rect 31435 37077 31447 37111
rect 31389 37071 31447 37077
rect 33594 37068 33600 37120
rect 33652 37108 33658 37120
rect 34164 37117 34192 37148
rect 34330 37136 34336 37148
rect 34388 37176 34394 37188
rect 35084 37176 35112 37207
rect 34388 37148 35112 37176
rect 34388 37136 34394 37148
rect 33981 37111 34039 37117
rect 33981 37108 33993 37111
rect 33652 37080 33993 37108
rect 33652 37068 33658 37080
rect 33981 37077 33993 37080
rect 34027 37077 34039 37111
rect 33981 37071 34039 37077
rect 34149 37111 34207 37117
rect 34149 37077 34161 37111
rect 34195 37077 34207 37111
rect 34974 37108 34980 37120
rect 34935 37080 34980 37108
rect 34149 37071 34207 37077
rect 34974 37068 34980 37080
rect 35032 37068 35038 37120
rect 36170 37108 36176 37120
rect 36131 37080 36176 37108
rect 36170 37068 36176 37080
rect 36228 37068 36234 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 22462 36864 22468 36916
rect 22520 36904 22526 36916
rect 22738 36904 22744 36916
rect 22520 36876 22744 36904
rect 22520 36864 22526 36876
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 24118 36904 24124 36916
rect 24079 36876 24124 36904
rect 24118 36864 24124 36876
rect 24176 36864 24182 36916
rect 25406 36864 25412 36916
rect 25464 36904 25470 36916
rect 25464 36876 26004 36904
rect 25464 36864 25470 36876
rect 16298 36836 16304 36848
rect 15212 36808 16304 36836
rect 15105 36771 15163 36777
rect 15105 36737 15117 36771
rect 15151 36737 15163 36771
rect 15105 36731 15163 36737
rect 15120 36632 15148 36731
rect 15212 36709 15240 36808
rect 16298 36796 16304 36808
rect 16356 36796 16362 36848
rect 22094 36836 22100 36848
rect 19628 36808 20668 36836
rect 22055 36808 22100 36836
rect 19628 36780 19656 36808
rect 16114 36768 16120 36780
rect 16075 36740 16120 36768
rect 16114 36728 16120 36740
rect 16172 36728 16178 36780
rect 17494 36768 17500 36780
rect 17455 36740 17500 36768
rect 17494 36728 17500 36740
rect 17552 36728 17558 36780
rect 18782 36768 18788 36780
rect 18743 36740 18788 36768
rect 18782 36728 18788 36740
rect 18840 36728 18846 36780
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 19610 36768 19616 36780
rect 19571 36740 19616 36768
rect 19610 36728 19616 36740
rect 19668 36728 19674 36780
rect 20162 36728 20168 36780
rect 20220 36768 20226 36780
rect 20640 36777 20668 36808
rect 22094 36796 22100 36808
rect 22152 36796 22158 36848
rect 22186 36796 22192 36848
rect 22244 36836 22250 36848
rect 22281 36839 22339 36845
rect 22281 36836 22293 36839
rect 22244 36808 22293 36836
rect 22244 36796 22250 36808
rect 22281 36805 22293 36808
rect 22327 36805 22339 36839
rect 24394 36836 24400 36848
rect 22281 36799 22339 36805
rect 23860 36808 24400 36836
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 20220 36740 20361 36768
rect 20220 36728 20226 36740
rect 20349 36737 20361 36740
rect 20395 36737 20407 36771
rect 20349 36731 20407 36737
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 20625 36771 20683 36777
rect 20625 36737 20637 36771
rect 20671 36737 20683 36771
rect 20625 36731 20683 36737
rect 15197 36703 15255 36709
rect 15197 36669 15209 36703
rect 15243 36669 15255 36703
rect 15197 36663 15255 36669
rect 15473 36703 15531 36709
rect 15473 36669 15485 36703
rect 15519 36700 15531 36703
rect 15562 36700 15568 36712
rect 15519 36672 15568 36700
rect 15519 36669 15531 36672
rect 15473 36663 15531 36669
rect 15562 36660 15568 36672
rect 15620 36660 15626 36712
rect 16850 36700 16856 36712
rect 16811 36672 16856 36700
rect 16850 36660 16856 36672
rect 16908 36660 16914 36712
rect 17773 36703 17831 36709
rect 17773 36669 17785 36703
rect 17819 36669 17831 36703
rect 17773 36663 17831 36669
rect 18877 36703 18935 36709
rect 18877 36669 18889 36703
rect 18923 36700 18935 36703
rect 19521 36703 19579 36709
rect 19521 36700 19533 36703
rect 18923 36672 19533 36700
rect 18923 36669 18935 36672
rect 18877 36663 18935 36669
rect 19521 36669 19533 36672
rect 19567 36669 19579 36703
rect 20456 36700 20484 36731
rect 20714 36728 20720 36780
rect 20772 36768 20778 36780
rect 22373 36771 22431 36777
rect 20772 36740 20817 36768
rect 20772 36728 20778 36740
rect 22373 36737 22385 36771
rect 22419 36737 22431 36771
rect 22373 36731 22431 36737
rect 22189 36703 22247 36709
rect 22189 36700 22201 36703
rect 20456 36672 22201 36700
rect 19521 36663 19579 36669
rect 16114 36632 16120 36644
rect 15120 36604 16120 36632
rect 16114 36592 16120 36604
rect 16172 36592 16178 36644
rect 17218 36592 17224 36644
rect 17276 36632 17282 36644
rect 17788 36632 17816 36663
rect 20640 36644 20668 36672
rect 22189 36669 22201 36672
rect 22235 36669 22247 36703
rect 22388 36700 22416 36731
rect 22462 36728 22468 36780
rect 22520 36777 22526 36780
rect 22520 36768 22528 36777
rect 23382 36768 23388 36780
rect 22520 36740 22565 36768
rect 22756 36740 23388 36768
rect 22520 36731 22528 36740
rect 22520 36728 22526 36731
rect 22756 36700 22784 36740
rect 23382 36728 23388 36740
rect 23440 36768 23446 36780
rect 23860 36768 23888 36808
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 25866 36836 25872 36848
rect 25516 36808 25872 36836
rect 23440 36740 23888 36768
rect 23937 36771 23995 36777
rect 23440 36728 23446 36740
rect 23937 36737 23949 36771
rect 23983 36768 23995 36771
rect 24026 36768 24032 36780
rect 23983 36740 24032 36768
rect 23983 36737 23995 36740
rect 23937 36731 23995 36737
rect 24026 36728 24032 36740
rect 24084 36728 24090 36780
rect 24210 36768 24216 36780
rect 24171 36740 24216 36768
rect 24210 36728 24216 36740
rect 24268 36728 24274 36780
rect 25317 36771 25375 36777
rect 25317 36737 25329 36771
rect 25363 36768 25375 36771
rect 25406 36768 25412 36780
rect 25363 36740 25412 36768
rect 25363 36737 25375 36740
rect 25317 36731 25375 36737
rect 25406 36728 25412 36740
rect 25464 36728 25470 36780
rect 25516 36777 25544 36808
rect 25866 36796 25872 36808
rect 25924 36796 25930 36848
rect 25501 36771 25559 36777
rect 25501 36737 25513 36771
rect 25547 36737 25559 36771
rect 25501 36731 25559 36737
rect 25777 36771 25835 36777
rect 25777 36737 25789 36771
rect 25823 36768 25835 36771
rect 25976 36768 26004 36876
rect 28994 36864 29000 36916
rect 29052 36904 29058 36916
rect 29914 36904 29920 36916
rect 29052 36876 29920 36904
rect 29052 36864 29058 36876
rect 29914 36864 29920 36876
rect 29972 36904 29978 36916
rect 31662 36904 31668 36916
rect 29972 36876 30880 36904
rect 31623 36876 31668 36904
rect 29972 36864 29978 36876
rect 26602 36796 26608 36848
rect 26660 36836 26666 36848
rect 27617 36839 27675 36845
rect 27617 36836 27629 36839
rect 26660 36808 27629 36836
rect 26660 36796 26666 36808
rect 27617 36805 27629 36808
rect 27663 36805 27675 36839
rect 28626 36836 28632 36848
rect 27617 36799 27675 36805
rect 27816 36808 28632 36836
rect 25823 36740 26004 36768
rect 26237 36771 26295 36777
rect 25823 36737 25835 36740
rect 25777 36731 25835 36737
rect 26237 36737 26249 36771
rect 26283 36768 26295 36771
rect 26510 36768 26516 36780
rect 26283 36740 26516 36768
rect 26283 36737 26295 36740
rect 26237 36731 26295 36737
rect 26510 36728 26516 36740
rect 26568 36728 26574 36780
rect 26970 36728 26976 36780
rect 27028 36768 27034 36780
rect 27816 36768 27844 36808
rect 28626 36796 28632 36808
rect 28684 36796 28690 36848
rect 28718 36796 28724 36848
rect 28776 36836 28782 36848
rect 29089 36839 29147 36845
rect 29089 36836 29101 36839
rect 28776 36808 29101 36836
rect 28776 36796 28782 36808
rect 29089 36805 29101 36808
rect 29135 36805 29147 36839
rect 30006 36836 30012 36848
rect 29089 36799 29147 36805
rect 29932 36808 30012 36836
rect 27028 36740 27844 36768
rect 27893 36771 27951 36777
rect 27028 36728 27034 36740
rect 27893 36737 27905 36771
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 22388 36672 22784 36700
rect 22189 36663 22247 36669
rect 22830 36660 22836 36712
rect 22888 36700 22894 36712
rect 23293 36703 23351 36709
rect 23293 36700 23305 36703
rect 22888 36672 23305 36700
rect 22888 36660 22894 36672
rect 23293 36669 23305 36672
rect 23339 36700 23351 36703
rect 24762 36700 24768 36712
rect 23339 36672 24768 36700
rect 23339 36669 23351 36672
rect 23293 36663 23351 36669
rect 24762 36660 24768 36672
rect 24820 36660 24826 36712
rect 25593 36703 25651 36709
rect 25593 36669 25605 36703
rect 25639 36669 25651 36703
rect 27908 36700 27936 36731
rect 28166 36728 28172 36780
rect 28224 36768 28230 36780
rect 28353 36771 28411 36777
rect 28353 36768 28365 36771
rect 28224 36740 28365 36768
rect 28224 36728 28230 36740
rect 28353 36737 28365 36740
rect 28399 36737 28411 36771
rect 28353 36731 28411 36737
rect 28537 36771 28595 36777
rect 28537 36737 28549 36771
rect 28583 36768 28595 36771
rect 28994 36768 29000 36780
rect 28583 36740 29000 36768
rect 28583 36737 28595 36740
rect 28537 36731 28595 36737
rect 28994 36728 29000 36740
rect 29052 36728 29058 36780
rect 29638 36728 29644 36780
rect 29696 36768 29702 36780
rect 29932 36777 29960 36808
rect 30006 36796 30012 36808
rect 30064 36796 30070 36848
rect 29825 36771 29883 36777
rect 29825 36768 29837 36771
rect 29696 36740 29837 36768
rect 29696 36728 29702 36740
rect 29825 36737 29837 36740
rect 29871 36737 29883 36771
rect 29825 36731 29883 36737
rect 29917 36771 29975 36777
rect 29917 36737 29929 36771
rect 29963 36737 29975 36771
rect 30466 36768 30472 36780
rect 29917 36731 29975 36737
rect 30024 36740 30472 36768
rect 28718 36700 28724 36712
rect 27908 36672 28724 36700
rect 25593 36663 25651 36669
rect 18417 36635 18475 36641
rect 18417 36632 18429 36635
rect 17276 36604 18429 36632
rect 17276 36592 17282 36604
rect 18417 36601 18429 36604
rect 18463 36601 18475 36635
rect 18417 36595 18475 36601
rect 20622 36592 20628 36644
rect 20680 36592 20686 36644
rect 21818 36592 21824 36644
rect 21876 36632 21882 36644
rect 25409 36635 25467 36641
rect 25409 36632 25421 36635
rect 21876 36604 25421 36632
rect 21876 36592 21882 36604
rect 25409 36601 25421 36604
rect 25455 36601 25467 36635
rect 25608 36632 25636 36663
rect 28718 36660 28724 36672
rect 28776 36700 28782 36712
rect 29730 36700 29736 36712
rect 28776 36672 29736 36700
rect 28776 36660 28782 36672
rect 29730 36660 29736 36672
rect 29788 36660 29794 36712
rect 30024 36709 30052 36740
rect 30466 36728 30472 36740
rect 30524 36728 30530 36780
rect 30653 36771 30711 36777
rect 30653 36737 30665 36771
rect 30699 36768 30711 36771
rect 30742 36768 30748 36780
rect 30699 36740 30748 36768
rect 30699 36737 30711 36740
rect 30653 36731 30711 36737
rect 30742 36728 30748 36740
rect 30800 36728 30806 36780
rect 30852 36777 30880 36876
rect 31662 36864 31668 36876
rect 31720 36904 31726 36916
rect 33870 36904 33876 36916
rect 31720 36864 31754 36904
rect 33831 36876 33876 36904
rect 33870 36864 33876 36876
rect 33928 36864 33934 36916
rect 31726 36836 31754 36864
rect 36170 36836 36176 36848
rect 31726 36808 32812 36836
rect 36018 36808 36176 36836
rect 30837 36771 30895 36777
rect 30837 36737 30849 36771
rect 30883 36737 30895 36771
rect 30837 36731 30895 36737
rect 31110 36728 31116 36780
rect 31168 36768 31174 36780
rect 31478 36768 31484 36780
rect 31168 36740 31484 36768
rect 31168 36728 31174 36740
rect 31478 36728 31484 36740
rect 31536 36728 31542 36780
rect 32490 36768 32496 36780
rect 32451 36740 32496 36768
rect 32490 36728 32496 36740
rect 32548 36728 32554 36780
rect 32674 36768 32680 36780
rect 32635 36740 32680 36768
rect 32674 36728 32680 36740
rect 32732 36728 32738 36780
rect 32784 36777 32812 36808
rect 36170 36796 36176 36808
rect 36228 36796 36234 36848
rect 32769 36771 32827 36777
rect 32769 36737 32781 36771
rect 32815 36737 32827 36771
rect 32769 36731 32827 36737
rect 33594 36728 33600 36780
rect 33652 36768 33658 36780
rect 33778 36768 33784 36780
rect 33652 36740 33784 36768
rect 33652 36728 33658 36740
rect 33778 36728 33784 36740
rect 33836 36728 33842 36780
rect 33870 36728 33876 36780
rect 33928 36768 33934 36780
rect 34057 36771 34115 36777
rect 34057 36768 34069 36771
rect 33928 36740 34069 36768
rect 33928 36728 33934 36740
rect 34057 36737 34069 36740
rect 34103 36737 34115 36771
rect 34974 36768 34980 36780
rect 34935 36740 34980 36768
rect 34057 36731 34115 36737
rect 34974 36728 34980 36740
rect 35032 36728 35038 36780
rect 30009 36703 30067 36709
rect 30009 36669 30021 36703
rect 30055 36669 30067 36703
rect 30009 36663 30067 36669
rect 30098 36660 30104 36712
rect 30156 36700 30162 36712
rect 31294 36700 31300 36712
rect 30156 36672 30201 36700
rect 31255 36672 31300 36700
rect 30156 36660 30162 36672
rect 31294 36660 31300 36672
rect 31352 36660 31358 36712
rect 34609 36703 34667 36709
rect 34609 36669 34621 36703
rect 34655 36700 34667 36703
rect 34790 36700 34796 36712
rect 34655 36672 34796 36700
rect 34655 36669 34667 36672
rect 34609 36663 34667 36669
rect 34790 36660 34796 36672
rect 34848 36700 34854 36712
rect 35434 36700 35440 36712
rect 34848 36672 35440 36700
rect 34848 36660 34854 36672
rect 35434 36660 35440 36672
rect 35492 36660 35498 36712
rect 36354 36700 36360 36712
rect 36315 36672 36360 36700
rect 36354 36660 36360 36672
rect 36412 36660 36418 36712
rect 32309 36635 32367 36641
rect 32309 36632 32321 36635
rect 25608 36604 32321 36632
rect 25409 36595 25467 36601
rect 32309 36601 32321 36604
rect 32355 36601 32367 36635
rect 33229 36635 33287 36641
rect 33229 36632 33241 36635
rect 32309 36595 32367 36601
rect 32508 36604 33241 36632
rect 15562 36524 15568 36576
rect 15620 36564 15626 36576
rect 15933 36567 15991 36573
rect 15933 36564 15945 36567
rect 15620 36536 15945 36564
rect 15620 36524 15626 36536
rect 15933 36533 15945 36536
rect 15979 36533 15991 36567
rect 15933 36527 15991 36533
rect 20901 36567 20959 36573
rect 20901 36533 20913 36567
rect 20947 36564 20959 36567
rect 20990 36564 20996 36576
rect 20947 36536 20996 36564
rect 20947 36533 20959 36536
rect 20901 36527 20959 36533
rect 20990 36524 20996 36536
rect 21048 36524 21054 36576
rect 21542 36524 21548 36576
rect 21600 36564 21606 36576
rect 23753 36567 23811 36573
rect 23753 36564 23765 36567
rect 21600 36536 23765 36564
rect 21600 36524 21606 36536
rect 23753 36533 23765 36536
rect 23799 36533 23811 36567
rect 23753 36527 23811 36533
rect 25133 36567 25191 36573
rect 25133 36533 25145 36567
rect 25179 36564 25191 36567
rect 25774 36564 25780 36576
rect 25179 36536 25780 36564
rect 25179 36533 25191 36536
rect 25133 36527 25191 36533
rect 25774 36524 25780 36536
rect 25832 36524 25838 36576
rect 26142 36524 26148 36576
rect 26200 36564 26206 36576
rect 26421 36567 26479 36573
rect 26421 36564 26433 36567
rect 26200 36536 26433 36564
rect 26200 36524 26206 36536
rect 26421 36533 26433 36536
rect 26467 36533 26479 36567
rect 26421 36527 26479 36533
rect 26786 36524 26792 36576
rect 26844 36564 26850 36576
rect 28074 36564 28080 36576
rect 26844 36536 28080 36564
rect 26844 36524 26850 36536
rect 28074 36524 28080 36536
rect 28132 36524 28138 36576
rect 28442 36564 28448 36576
rect 28403 36536 28448 36564
rect 28442 36524 28448 36536
rect 28500 36524 28506 36576
rect 29638 36564 29644 36576
rect 29599 36536 29644 36564
rect 29638 36524 29644 36536
rect 29696 36524 29702 36576
rect 30745 36567 30803 36573
rect 30745 36533 30757 36567
rect 30791 36564 30803 36567
rect 30926 36564 30932 36576
rect 30791 36536 30932 36564
rect 30791 36533 30803 36536
rect 30745 36527 30803 36533
rect 30926 36524 30932 36536
rect 30984 36564 30990 36576
rect 31110 36564 31116 36576
rect 30984 36536 31116 36564
rect 30984 36524 30990 36536
rect 31110 36524 31116 36536
rect 31168 36524 31174 36576
rect 31478 36524 31484 36576
rect 31536 36564 31542 36576
rect 32508 36564 32536 36604
rect 33229 36601 33241 36604
rect 33275 36601 33287 36635
rect 34054 36632 34060 36644
rect 34015 36604 34060 36632
rect 33229 36595 33287 36601
rect 34054 36592 34060 36604
rect 34112 36592 34118 36644
rect 31536 36536 32536 36564
rect 31536 36524 31542 36536
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 17494 36360 17500 36372
rect 17455 36332 17500 36360
rect 17494 36320 17500 36332
rect 17552 36320 17558 36372
rect 17586 36320 17592 36372
rect 17644 36360 17650 36372
rect 18417 36363 18475 36369
rect 18417 36360 18429 36363
rect 17644 36332 18429 36360
rect 17644 36320 17650 36332
rect 18417 36329 18429 36332
rect 18463 36329 18475 36363
rect 18417 36323 18475 36329
rect 18647 36363 18705 36369
rect 18647 36329 18659 36363
rect 18693 36360 18705 36363
rect 19610 36360 19616 36372
rect 18693 36332 19616 36360
rect 18693 36329 18705 36332
rect 18647 36323 18705 36329
rect 19610 36320 19616 36332
rect 19668 36360 19674 36372
rect 21177 36363 21235 36369
rect 21177 36360 21189 36363
rect 19668 36332 21189 36360
rect 19668 36320 19674 36332
rect 21177 36329 21189 36332
rect 21223 36329 21235 36363
rect 21177 36323 21235 36329
rect 24762 36320 24768 36372
rect 24820 36360 24826 36372
rect 25682 36360 25688 36372
rect 24820 36332 25688 36360
rect 24820 36320 24826 36332
rect 25682 36320 25688 36332
rect 25740 36360 25746 36372
rect 27617 36363 27675 36369
rect 25740 36332 27200 36360
rect 25740 36320 25746 36332
rect 19426 36292 19432 36304
rect 18524 36264 19432 36292
rect 17681 36227 17739 36233
rect 17681 36193 17693 36227
rect 17727 36193 17739 36227
rect 17681 36187 17739 36193
rect 17218 36156 17224 36168
rect 17179 36128 17224 36156
rect 17218 36116 17224 36128
rect 17276 36116 17282 36168
rect 17696 36156 17724 36187
rect 18524 36168 18552 36264
rect 19426 36252 19432 36264
rect 19484 36252 19490 36304
rect 20346 36292 20352 36304
rect 19536 36264 20352 36292
rect 18325 36159 18383 36165
rect 18325 36156 18337 36159
rect 17696 36128 18337 36156
rect 18325 36125 18337 36128
rect 18371 36125 18383 36159
rect 18506 36156 18512 36168
rect 18467 36128 18512 36156
rect 18325 36119 18383 36125
rect 18506 36116 18512 36128
rect 18564 36116 18570 36168
rect 18782 36156 18788 36168
rect 18743 36128 18788 36156
rect 18782 36116 18788 36128
rect 18840 36116 18846 36168
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 19392 36128 19441 36156
rect 19392 36116 19398 36128
rect 19429 36125 19441 36128
rect 19475 36156 19487 36159
rect 19536 36156 19564 36264
rect 20346 36252 20352 36264
rect 20404 36292 20410 36304
rect 20714 36292 20720 36304
rect 20404 36264 20720 36292
rect 20404 36252 20410 36264
rect 20714 36252 20720 36264
rect 20772 36252 20778 36304
rect 23198 36292 23204 36304
rect 22296 36264 23204 36292
rect 20622 36224 20628 36236
rect 20583 36196 20628 36224
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 21542 36224 21548 36236
rect 21503 36196 21548 36224
rect 21542 36184 21548 36196
rect 21600 36184 21606 36236
rect 19475 36128 19564 36156
rect 19613 36159 19671 36165
rect 19475 36125 19487 36128
rect 19429 36119 19487 36125
rect 19613 36125 19625 36159
rect 19659 36125 19671 36159
rect 19613 36119 19671 36125
rect 19628 36088 19656 36119
rect 20162 36116 20168 36168
rect 20220 36156 20226 36168
rect 20257 36159 20315 36165
rect 20257 36156 20269 36159
rect 20220 36128 20269 36156
rect 20220 36116 20226 36128
rect 20257 36125 20269 36128
rect 20303 36125 20315 36159
rect 20530 36156 20536 36168
rect 20491 36128 20536 36156
rect 20257 36119 20315 36125
rect 20530 36116 20536 36128
rect 20588 36116 20594 36168
rect 21358 36156 21364 36168
rect 21319 36128 21364 36156
rect 21358 36116 21364 36128
rect 21416 36116 21422 36168
rect 22296 36156 22324 36264
rect 23198 36252 23204 36264
rect 23256 36292 23262 36304
rect 26510 36292 26516 36304
rect 23256 36264 26516 36292
rect 23256 36252 23262 36264
rect 22370 36184 22376 36236
rect 22428 36224 22434 36236
rect 22649 36227 22707 36233
rect 22649 36224 22661 36227
rect 22428 36196 22661 36224
rect 22428 36184 22434 36196
rect 22649 36193 22661 36196
rect 22695 36193 22707 36227
rect 22649 36187 22707 36193
rect 22741 36227 22799 36233
rect 22741 36193 22753 36227
rect 22787 36224 22799 36227
rect 22922 36224 22928 36236
rect 22787 36196 22928 36224
rect 22787 36193 22799 36196
rect 22741 36187 22799 36193
rect 22922 36184 22928 36196
rect 22980 36224 22986 36236
rect 24578 36224 24584 36236
rect 22980 36196 24584 36224
rect 22980 36184 22986 36196
rect 24578 36184 24584 36196
rect 24636 36184 24642 36236
rect 22557 36159 22615 36165
rect 22557 36156 22569 36159
rect 22296 36128 22569 36156
rect 22557 36125 22569 36128
rect 22603 36125 22615 36159
rect 22557 36119 22615 36125
rect 22833 36159 22891 36165
rect 22833 36125 22845 36159
rect 22879 36156 22891 36159
rect 24486 36156 24492 36168
rect 22879 36128 24492 36156
rect 22879 36125 22891 36128
rect 22833 36119 22891 36125
rect 24486 36116 24492 36128
rect 24544 36116 24550 36168
rect 24688 36156 24716 36264
rect 26510 36252 26516 36264
rect 26568 36252 26574 36304
rect 27062 36292 27068 36304
rect 27023 36264 27068 36292
rect 27062 36252 27068 36264
rect 27120 36252 27126 36304
rect 27172 36292 27200 36332
rect 27617 36329 27629 36363
rect 27663 36360 27675 36363
rect 28902 36360 28908 36372
rect 27663 36332 28908 36360
rect 27663 36329 27675 36332
rect 27617 36323 27675 36329
rect 28902 36320 28908 36332
rect 28960 36320 28966 36372
rect 28994 36320 29000 36372
rect 29052 36360 29058 36372
rect 30098 36360 30104 36372
rect 29052 36332 30104 36360
rect 29052 36320 29058 36332
rect 30098 36320 30104 36332
rect 30156 36360 30162 36372
rect 30834 36360 30840 36372
rect 30156 36332 30840 36360
rect 30156 36320 30162 36332
rect 30834 36320 30840 36332
rect 30892 36360 30898 36372
rect 31113 36363 31171 36369
rect 31113 36360 31125 36363
rect 30892 36332 31125 36360
rect 30892 36320 30898 36332
rect 31113 36329 31125 36332
rect 31159 36329 31171 36363
rect 31113 36323 31171 36329
rect 31294 36320 31300 36372
rect 31352 36360 31358 36372
rect 31757 36363 31815 36369
rect 31757 36360 31769 36363
rect 31352 36332 31769 36360
rect 31352 36320 31358 36332
rect 31757 36329 31769 36332
rect 31803 36360 31815 36363
rect 33134 36360 33140 36372
rect 31803 36332 33140 36360
rect 31803 36329 31815 36332
rect 31757 36323 31815 36329
rect 33134 36320 33140 36332
rect 33192 36320 33198 36372
rect 27172 36264 27660 36292
rect 27632 36236 27660 36264
rect 28626 36252 28632 36304
rect 28684 36292 28690 36304
rect 33410 36292 33416 36304
rect 28684 36264 33416 36292
rect 28684 36252 28690 36264
rect 33410 36252 33416 36264
rect 33468 36292 33474 36304
rect 33597 36295 33655 36301
rect 33597 36292 33609 36295
rect 33468 36264 33609 36292
rect 33468 36252 33474 36264
rect 33597 36261 33609 36264
rect 33643 36292 33655 36295
rect 33870 36292 33876 36304
rect 33643 36264 33876 36292
rect 33643 36261 33655 36264
rect 33597 36255 33655 36261
rect 33870 36252 33876 36264
rect 33928 36252 33934 36304
rect 24765 36227 24823 36233
rect 24765 36193 24777 36227
rect 24811 36224 24823 36227
rect 25593 36227 25651 36233
rect 25593 36224 25605 36227
rect 24811 36196 25605 36224
rect 24811 36193 24823 36196
rect 24765 36187 24823 36193
rect 25593 36193 25605 36196
rect 25639 36193 25651 36227
rect 25593 36187 25651 36193
rect 26436 36196 27568 36224
rect 26436 36168 26464 36196
rect 24857 36159 24915 36165
rect 24857 36156 24869 36159
rect 24688 36128 24869 36156
rect 24857 36125 24869 36128
rect 24903 36125 24915 36159
rect 24857 36119 24915 36125
rect 24949 36159 25007 36165
rect 24949 36125 24961 36159
rect 24995 36125 25007 36159
rect 24949 36119 25007 36125
rect 20548 36088 20576 36116
rect 19628 36060 20576 36088
rect 21910 36048 21916 36100
rect 21968 36088 21974 36100
rect 23477 36091 23535 36097
rect 23477 36088 23489 36091
rect 21968 36060 23489 36088
rect 21968 36048 21974 36060
rect 23477 36057 23489 36060
rect 23523 36057 23535 36091
rect 23842 36088 23848 36100
rect 23803 36060 23848 36088
rect 23477 36051 23535 36057
rect 23842 36048 23848 36060
rect 23900 36048 23906 36100
rect 24210 36048 24216 36100
rect 24268 36088 24274 36100
rect 24964 36088 24992 36119
rect 25038 36116 25044 36168
rect 25096 36156 25102 36168
rect 25961 36159 26019 36165
rect 25096 36128 25141 36156
rect 25096 36116 25102 36128
rect 25961 36125 25973 36159
rect 26007 36156 26019 36159
rect 26418 36156 26424 36168
rect 26007 36128 26424 36156
rect 26007 36125 26019 36128
rect 25961 36119 26019 36125
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 26786 36156 26792 36168
rect 26747 36128 26792 36156
rect 26786 36116 26792 36128
rect 26844 36116 26850 36168
rect 26878 36116 26884 36168
rect 26936 36156 26942 36168
rect 27540 36165 27568 36196
rect 27614 36184 27620 36236
rect 27672 36224 27678 36236
rect 27801 36227 27859 36233
rect 27801 36224 27813 36227
rect 27672 36196 27813 36224
rect 27672 36184 27678 36196
rect 27801 36193 27813 36196
rect 27847 36193 27859 36227
rect 30009 36227 30067 36233
rect 30009 36224 30021 36227
rect 27801 36187 27859 36193
rect 27908 36196 30021 36224
rect 27525 36159 27583 36165
rect 26936 36128 26981 36156
rect 26936 36116 26942 36128
rect 27525 36125 27537 36159
rect 27571 36125 27583 36159
rect 27908 36156 27936 36196
rect 30009 36193 30021 36196
rect 30055 36224 30067 36227
rect 30650 36224 30656 36236
rect 30055 36196 30656 36224
rect 30055 36193 30067 36196
rect 30009 36187 30067 36193
rect 30650 36184 30656 36196
rect 30708 36184 30714 36236
rect 31297 36227 31355 36233
rect 31297 36224 31309 36227
rect 30760 36196 31309 36224
rect 27525 36119 27583 36125
rect 27632 36128 27936 36156
rect 24268 36060 24992 36088
rect 24268 36048 24274 36060
rect 25590 36048 25596 36100
rect 25648 36088 25654 36100
rect 25777 36091 25835 36097
rect 25777 36088 25789 36091
rect 25648 36060 25789 36088
rect 25648 36048 25654 36060
rect 25777 36057 25789 36060
rect 25823 36057 25835 36091
rect 25777 36051 25835 36057
rect 26970 36048 26976 36100
rect 27028 36088 27034 36100
rect 27065 36091 27123 36097
rect 27065 36088 27077 36091
rect 27028 36060 27077 36088
rect 27028 36048 27034 36060
rect 27065 36057 27077 36060
rect 27111 36057 27123 36091
rect 27065 36051 27123 36057
rect 19426 35980 19432 36032
rect 19484 36020 19490 36032
rect 19521 36023 19579 36029
rect 19521 36020 19533 36023
rect 19484 35992 19533 36020
rect 19484 35980 19490 35992
rect 19521 35989 19533 35992
rect 19567 35989 19579 36023
rect 20714 36020 20720 36032
rect 20675 35992 20720 36020
rect 19521 35983 19579 35989
rect 20714 35980 20720 35992
rect 20772 35980 20778 36032
rect 22094 35980 22100 36032
rect 22152 36020 22158 36032
rect 22373 36023 22431 36029
rect 22373 36020 22385 36023
rect 22152 35992 22385 36020
rect 22152 35980 22158 35992
rect 22373 35989 22385 35992
rect 22419 35989 22431 36023
rect 22373 35983 22431 35989
rect 24581 36023 24639 36029
rect 24581 35989 24593 36023
rect 24627 36020 24639 36023
rect 24762 36020 24768 36032
rect 24627 35992 24768 36020
rect 24627 35989 24639 35992
rect 24581 35983 24639 35989
rect 24762 35980 24768 35992
rect 24820 35980 24826 36032
rect 24854 35980 24860 36032
rect 24912 36020 24918 36032
rect 27632 36020 27660 36128
rect 28258 36116 28264 36168
rect 28316 36156 28322 36168
rect 29089 36159 29147 36165
rect 28316 36128 28856 36156
rect 28316 36116 28322 36128
rect 28718 36088 28724 36100
rect 28679 36060 28724 36088
rect 28718 36048 28724 36060
rect 28776 36048 28782 36100
rect 28828 36088 28856 36128
rect 29089 36125 29101 36159
rect 29135 36156 29147 36159
rect 29178 36156 29184 36168
rect 29135 36128 29184 36156
rect 29135 36125 29147 36128
rect 29089 36119 29147 36125
rect 29178 36116 29184 36128
rect 29236 36116 29242 36168
rect 29917 36159 29975 36165
rect 29917 36125 29929 36159
rect 29963 36156 29975 36159
rect 30374 36156 30380 36168
rect 29963 36128 30380 36156
rect 29963 36125 29975 36128
rect 29917 36119 29975 36125
rect 30374 36116 30380 36128
rect 30432 36116 30438 36168
rect 30558 36116 30564 36168
rect 30616 36156 30622 36168
rect 30760 36156 30788 36196
rect 31297 36193 31309 36196
rect 31343 36193 31355 36227
rect 32674 36224 32680 36236
rect 32635 36196 32680 36224
rect 31297 36187 31355 36193
rect 32674 36184 32680 36196
rect 32732 36184 32738 36236
rect 34698 36184 34704 36236
rect 34756 36224 34762 36236
rect 34756 36196 35204 36224
rect 34756 36184 34762 36196
rect 31018 36156 31024 36168
rect 30616 36128 30788 36156
rect 30979 36128 31024 36156
rect 30616 36116 30622 36128
rect 31018 36116 31024 36128
rect 31076 36116 31082 36168
rect 31478 36156 31484 36168
rect 31128 36128 31484 36156
rect 31128 36088 31156 36128
rect 31478 36116 31484 36128
rect 31536 36116 31542 36168
rect 32766 36156 32772 36168
rect 32727 36128 32772 36156
rect 32766 36116 32772 36128
rect 32824 36116 32830 36168
rect 33134 36116 33140 36168
rect 33192 36156 33198 36168
rect 33413 36159 33471 36165
rect 33413 36156 33425 36159
rect 33192 36128 33425 36156
rect 33192 36116 33198 36128
rect 33413 36125 33425 36128
rect 33459 36125 33471 36159
rect 33413 36119 33471 36125
rect 33502 36116 33508 36168
rect 33560 36156 33566 36168
rect 34149 36159 34207 36165
rect 34149 36156 34161 36159
rect 33560 36128 34161 36156
rect 33560 36116 33566 36128
rect 34149 36125 34161 36128
rect 34195 36125 34207 36159
rect 34330 36156 34336 36168
rect 34291 36128 34336 36156
rect 34149 36119 34207 36125
rect 34330 36116 34336 36128
rect 34388 36116 34394 36168
rect 34882 36156 34888 36168
rect 34843 36128 34888 36156
rect 34882 36116 34888 36128
rect 34940 36116 34946 36168
rect 35176 36165 35204 36196
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36125 35127 36159
rect 35069 36119 35127 36125
rect 35161 36159 35219 36165
rect 35161 36125 35173 36159
rect 35207 36125 35219 36159
rect 35161 36119 35219 36125
rect 28828 36060 31156 36088
rect 31297 36091 31355 36097
rect 31297 36057 31309 36091
rect 31343 36088 31355 36091
rect 32122 36088 32128 36100
rect 31343 36060 32128 36088
rect 31343 36057 31355 36060
rect 31297 36051 31355 36057
rect 32122 36048 32128 36060
rect 32180 36048 32186 36100
rect 35084 36088 35112 36119
rect 35250 36116 35256 36168
rect 35308 36156 35314 36168
rect 36541 36159 36599 36165
rect 36541 36156 36553 36159
rect 35308 36128 36553 36156
rect 35308 36116 35314 36128
rect 36541 36125 36553 36128
rect 36587 36125 36599 36159
rect 36541 36119 36599 36125
rect 34164 36060 35112 36088
rect 24912 35992 27660 36020
rect 27801 36023 27859 36029
rect 24912 35980 24918 35992
rect 27801 35989 27813 36023
rect 27847 36020 27859 36023
rect 27890 36020 27896 36032
rect 27847 35992 27896 36020
rect 27847 35989 27859 35992
rect 27801 35983 27859 35989
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 30282 36020 30288 36032
rect 30243 35992 30288 36020
rect 30282 35980 30288 35992
rect 30340 35980 30346 36032
rect 31938 35980 31944 36032
rect 31996 36020 32002 36032
rect 32401 36023 32459 36029
rect 32401 36020 32413 36023
rect 31996 35992 32413 36020
rect 31996 35980 32002 35992
rect 32401 35989 32413 35992
rect 32447 35989 32459 36023
rect 32401 35983 32459 35989
rect 33962 35980 33968 36032
rect 34020 36020 34026 36032
rect 34164 36029 34192 36060
rect 34149 36023 34207 36029
rect 34149 36020 34161 36023
rect 34020 35992 34161 36020
rect 34020 35980 34026 35992
rect 34149 35989 34161 35992
rect 34195 35989 34207 36023
rect 34149 35983 34207 35989
rect 35158 35980 35164 36032
rect 35216 36020 35222 36032
rect 35529 36023 35587 36029
rect 35529 36020 35541 36023
rect 35216 35992 35541 36020
rect 35216 35980 35222 35992
rect 35529 35989 35541 35992
rect 35575 35989 35587 36023
rect 35529 35983 35587 35989
rect 36081 36023 36139 36029
rect 36081 35989 36093 36023
rect 36127 36020 36139 36023
rect 36170 36020 36176 36032
rect 36127 35992 36176 36020
rect 36127 35989 36139 35992
rect 36081 35983 36139 35989
rect 36170 35980 36176 35992
rect 36228 35980 36234 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 14185 35819 14243 35825
rect 14185 35785 14197 35819
rect 14231 35816 14243 35819
rect 14274 35816 14280 35828
rect 14231 35788 14280 35816
rect 14231 35785 14243 35788
rect 14185 35779 14243 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 15562 35776 15568 35828
rect 15620 35776 15626 35828
rect 16114 35776 16120 35828
rect 16172 35816 16178 35828
rect 16853 35819 16911 35825
rect 16853 35816 16865 35819
rect 16172 35788 16865 35816
rect 16172 35776 16178 35788
rect 16853 35785 16865 35788
rect 16899 35785 16911 35819
rect 16853 35779 16911 35785
rect 20625 35819 20683 35825
rect 20625 35785 20637 35819
rect 20671 35816 20683 35819
rect 23750 35816 23756 35828
rect 20671 35788 23756 35816
rect 20671 35785 20683 35788
rect 20625 35779 20683 35785
rect 23750 35776 23756 35788
rect 23808 35776 23814 35828
rect 24486 35776 24492 35828
rect 24544 35816 24550 35828
rect 25041 35819 25099 35825
rect 25041 35816 25053 35819
rect 24544 35788 25053 35816
rect 24544 35776 24550 35788
rect 25041 35785 25053 35788
rect 25087 35785 25099 35819
rect 28074 35816 28080 35828
rect 25041 35779 25099 35785
rect 25424 35788 28080 35816
rect 14737 35751 14795 35757
rect 14737 35717 14749 35751
rect 14783 35748 14795 35751
rect 15194 35748 15200 35760
rect 14783 35720 15200 35748
rect 14783 35717 14795 35720
rect 14737 35711 14795 35717
rect 15194 35708 15200 35720
rect 15252 35748 15258 35760
rect 15378 35748 15384 35760
rect 15252 35720 15384 35748
rect 15252 35708 15258 35720
rect 15378 35708 15384 35720
rect 15436 35708 15442 35760
rect 15580 35748 15608 35776
rect 21450 35748 21456 35760
rect 15580 35720 15884 35748
rect 21411 35720 21456 35748
rect 14090 35680 14096 35692
rect 14051 35652 14096 35680
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 14277 35683 14335 35689
rect 14277 35649 14289 35683
rect 14323 35649 14335 35683
rect 14918 35680 14924 35692
rect 14879 35652 14924 35680
rect 14277 35643 14335 35649
rect 14292 35612 14320 35643
rect 14918 35640 14924 35652
rect 14976 35640 14982 35692
rect 15010 35640 15016 35692
rect 15068 35680 15074 35692
rect 15565 35683 15623 35689
rect 15565 35680 15577 35683
rect 15068 35652 15577 35680
rect 15068 35640 15074 35652
rect 15565 35649 15577 35652
rect 15611 35649 15623 35683
rect 15746 35680 15752 35692
rect 15707 35652 15752 35680
rect 15565 35643 15623 35649
rect 15746 35640 15752 35652
rect 15804 35640 15810 35692
rect 15856 35689 15884 35720
rect 21450 35708 21456 35720
rect 21508 35708 21514 35760
rect 22830 35748 22836 35760
rect 22791 35720 22836 35748
rect 22830 35708 22836 35720
rect 22888 35708 22894 35760
rect 22925 35751 22983 35757
rect 22925 35717 22937 35751
rect 22971 35748 22983 35751
rect 23106 35748 23112 35760
rect 22971 35720 23112 35748
rect 22971 35717 22983 35720
rect 22925 35711 22983 35717
rect 23106 35708 23112 35720
rect 23164 35748 23170 35760
rect 24210 35748 24216 35760
rect 23164 35720 23888 35748
rect 24171 35720 24216 35748
rect 23164 35708 23170 35720
rect 23860 35692 23888 35720
rect 24210 35708 24216 35720
rect 24268 35708 24274 35760
rect 25424 35757 25452 35788
rect 28074 35776 28080 35788
rect 28132 35776 28138 35828
rect 28994 35776 29000 35828
rect 29052 35776 29058 35828
rect 29288 35788 31340 35816
rect 25409 35751 25467 35757
rect 25409 35717 25421 35751
rect 25455 35717 25467 35751
rect 26142 35748 26148 35760
rect 25409 35711 25467 35717
rect 25516 35720 26148 35748
rect 15841 35683 15899 35689
rect 15841 35649 15853 35683
rect 15887 35649 15899 35683
rect 15841 35643 15899 35649
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 15988 35652 16033 35680
rect 15988 35640 15994 35652
rect 17034 35640 17040 35692
rect 17092 35680 17098 35692
rect 17221 35683 17279 35689
rect 17221 35680 17233 35683
rect 17092 35652 17233 35680
rect 17092 35640 17098 35652
rect 17221 35649 17233 35652
rect 17267 35680 17279 35683
rect 17267 35652 19104 35680
rect 17267 35649 17279 35652
rect 17221 35643 17279 35649
rect 17126 35612 17132 35624
rect 14292 35584 14780 35612
rect 17087 35584 17132 35612
rect 14752 35553 14780 35584
rect 17126 35572 17132 35584
rect 17184 35572 17190 35624
rect 19076 35553 19104 35652
rect 19518 35640 19524 35692
rect 19576 35680 19582 35692
rect 19613 35683 19671 35689
rect 19613 35680 19625 35683
rect 19576 35652 19625 35680
rect 19576 35640 19582 35652
rect 19613 35649 19625 35652
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 19702 35640 19708 35692
rect 19760 35680 19766 35692
rect 20070 35680 20076 35692
rect 19760 35652 20076 35680
rect 19760 35640 19766 35652
rect 20070 35640 20076 35652
rect 20128 35640 20134 35692
rect 20257 35683 20315 35689
rect 20257 35649 20269 35683
rect 20303 35680 20315 35683
rect 20346 35680 20352 35692
rect 20303 35652 20352 35680
rect 20303 35649 20315 35652
rect 20257 35643 20315 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20441 35683 20499 35689
rect 20441 35649 20453 35683
rect 20487 35680 20499 35683
rect 20530 35680 20536 35692
rect 20487 35652 20536 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 20530 35640 20536 35652
rect 20588 35640 20594 35692
rect 22278 35640 22284 35692
rect 22336 35680 22342 35692
rect 22738 35689 22744 35692
rect 22557 35683 22615 35689
rect 22557 35680 22569 35683
rect 22336 35652 22569 35680
rect 22336 35640 22342 35652
rect 22557 35649 22569 35652
rect 22603 35649 22615 35683
rect 22557 35643 22615 35649
rect 22705 35683 22744 35689
rect 22705 35649 22717 35683
rect 22705 35643 22744 35649
rect 19337 35615 19395 35621
rect 19337 35581 19349 35615
rect 19383 35581 19395 35615
rect 20162 35612 20168 35624
rect 20075 35584 20168 35612
rect 19337 35575 19395 35581
rect 14737 35547 14795 35553
rect 14737 35513 14749 35547
rect 14783 35513 14795 35547
rect 14737 35507 14795 35513
rect 19061 35547 19119 35553
rect 19061 35513 19073 35547
rect 19107 35513 19119 35547
rect 19352 35544 19380 35575
rect 20162 35572 20168 35584
rect 20220 35612 20226 35624
rect 20898 35612 20904 35624
rect 20220 35584 20904 35612
rect 20220 35572 20226 35584
rect 20898 35572 20904 35584
rect 20956 35572 20962 35624
rect 22572 35612 22600 35643
rect 22738 35640 22744 35643
rect 22796 35640 22802 35692
rect 23014 35640 23020 35692
rect 23072 35689 23078 35692
rect 23072 35680 23080 35689
rect 23072 35652 23117 35680
rect 23072 35643 23080 35652
rect 23072 35640 23078 35643
rect 23842 35640 23848 35692
rect 23900 35680 23906 35692
rect 24397 35683 24455 35689
rect 24397 35680 24409 35683
rect 23900 35652 24409 35680
rect 23900 35640 23906 35652
rect 24397 35649 24409 35652
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 24581 35683 24639 35689
rect 24581 35649 24593 35683
rect 24627 35680 24639 35683
rect 25225 35683 25283 35689
rect 25225 35680 25237 35683
rect 24627 35652 25237 35680
rect 24627 35649 24639 35652
rect 24581 35643 24639 35649
rect 25225 35649 25237 35652
rect 25271 35649 25283 35683
rect 25225 35643 25283 35649
rect 25317 35683 25375 35689
rect 25317 35649 25329 35683
rect 25363 35680 25375 35683
rect 25516 35680 25544 35720
rect 26142 35708 26148 35720
rect 26200 35708 26206 35760
rect 27062 35708 27068 35760
rect 27120 35748 27126 35760
rect 27157 35751 27215 35757
rect 27157 35748 27169 35751
rect 27120 35720 27169 35748
rect 27120 35708 27126 35720
rect 27157 35717 27169 35720
rect 27203 35717 27215 35751
rect 27338 35748 27344 35760
rect 27299 35720 27344 35748
rect 27157 35711 27215 35717
rect 27338 35708 27344 35720
rect 27396 35708 27402 35760
rect 29012 35748 29040 35776
rect 28184 35720 29040 35748
rect 25363 35652 25544 35680
rect 25593 35683 25651 35689
rect 25363 35649 25375 35652
rect 25317 35643 25375 35649
rect 25593 35649 25605 35683
rect 25639 35680 25651 35683
rect 25682 35680 25688 35692
rect 25639 35652 25688 35680
rect 25639 35649 25651 35652
rect 25593 35643 25651 35649
rect 23934 35612 23940 35624
rect 22572 35584 23940 35612
rect 23934 35572 23940 35584
rect 23992 35572 23998 35624
rect 24412 35612 24440 35643
rect 25682 35640 25688 35652
rect 25740 35640 25746 35692
rect 25866 35640 25872 35692
rect 25924 35680 25930 35692
rect 26421 35683 26479 35689
rect 26421 35680 26433 35683
rect 25924 35652 26433 35680
rect 25924 35640 25930 35652
rect 26421 35649 26433 35652
rect 26467 35649 26479 35683
rect 26421 35643 26479 35649
rect 26605 35683 26663 35689
rect 26605 35649 26617 35683
rect 26651 35680 26663 35683
rect 26878 35680 26884 35692
rect 26651 35652 26884 35680
rect 26651 35649 26663 35652
rect 26605 35643 26663 35649
rect 26878 35640 26884 35652
rect 26936 35640 26942 35692
rect 28184 35689 28212 35720
rect 27985 35683 28043 35689
rect 27985 35649 27997 35683
rect 28031 35649 28043 35683
rect 27985 35643 28043 35649
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35649 28227 35683
rect 28169 35643 28227 35649
rect 25406 35612 25412 35624
rect 24412 35584 25412 35612
rect 25406 35572 25412 35584
rect 25464 35612 25470 35624
rect 26326 35612 26332 35624
rect 25464 35584 26332 35612
rect 25464 35572 25470 35584
rect 26326 35572 26332 35584
rect 26384 35572 26390 35624
rect 26513 35615 26571 35621
rect 26513 35581 26525 35615
rect 26559 35612 26571 35615
rect 28000 35612 28028 35643
rect 28442 35640 28448 35692
rect 28500 35680 28506 35692
rect 28902 35680 28908 35692
rect 28500 35652 28908 35680
rect 28500 35640 28506 35652
rect 28902 35640 28908 35652
rect 28960 35680 28966 35692
rect 28997 35683 29055 35689
rect 28997 35680 29009 35683
rect 28960 35652 29009 35680
rect 28960 35640 28966 35652
rect 28997 35649 29009 35652
rect 29043 35649 29055 35683
rect 29178 35680 29184 35692
rect 29139 35652 29184 35680
rect 28997 35643 29055 35649
rect 29178 35640 29184 35652
rect 29236 35640 29242 35692
rect 26559 35584 28028 35612
rect 28721 35615 28779 35621
rect 26559 35581 26571 35584
rect 26513 35575 26571 35581
rect 26620 35556 26648 35584
rect 28721 35581 28733 35615
rect 28767 35612 28779 35615
rect 29086 35612 29092 35624
rect 28767 35584 29092 35612
rect 28767 35581 28779 35584
rect 28721 35575 28779 35581
rect 29086 35572 29092 35584
rect 29144 35572 29150 35624
rect 20070 35544 20076 35556
rect 19061 35507 19119 35513
rect 19260 35516 20076 35544
rect 18506 35436 18512 35488
rect 18564 35476 18570 35488
rect 18601 35479 18659 35485
rect 18601 35476 18613 35479
rect 18564 35448 18613 35476
rect 18564 35436 18570 35448
rect 18601 35445 18613 35448
rect 18647 35476 18659 35479
rect 19260 35476 19288 35516
rect 20070 35504 20076 35516
rect 20128 35504 20134 35556
rect 23753 35547 23811 35553
rect 23753 35513 23765 35547
rect 23799 35544 23811 35547
rect 25590 35544 25596 35556
rect 23799 35516 25596 35544
rect 23799 35513 23811 35516
rect 23753 35507 23811 35513
rect 25590 35504 25596 35516
rect 25648 35504 25654 35556
rect 26602 35504 26608 35556
rect 26660 35504 26666 35556
rect 29288 35544 29316 35788
rect 29822 35708 29828 35760
rect 29880 35748 29886 35760
rect 30101 35751 30159 35757
rect 30101 35748 30113 35751
rect 29880 35720 30113 35748
rect 29880 35708 29886 35720
rect 30101 35717 30113 35720
rect 30147 35717 30159 35751
rect 31312 35748 31340 35788
rect 31386 35776 31392 35828
rect 31444 35816 31450 35828
rect 31757 35819 31815 35825
rect 31757 35816 31769 35819
rect 31444 35788 31769 35816
rect 31444 35776 31450 35788
rect 31757 35785 31769 35788
rect 31803 35816 31815 35819
rect 32509 35819 32567 35825
rect 32509 35816 32521 35819
rect 31803 35788 32521 35816
rect 31803 35785 31815 35788
rect 31757 35779 31815 35785
rect 32509 35785 32521 35788
rect 32555 35785 32567 35819
rect 32674 35816 32680 35828
rect 32635 35788 32680 35816
rect 32509 35779 32567 35785
rect 32674 35776 32680 35788
rect 32732 35776 32738 35828
rect 33321 35819 33379 35825
rect 33321 35785 33333 35819
rect 33367 35816 33379 35819
rect 33502 35816 33508 35828
rect 33367 35788 33508 35816
rect 33367 35785 33379 35788
rect 33321 35779 33379 35785
rect 33502 35776 33508 35788
rect 33560 35776 33566 35828
rect 34333 35819 34391 35825
rect 34333 35785 34345 35819
rect 34379 35816 34391 35819
rect 34882 35816 34888 35828
rect 34379 35788 34888 35816
rect 34379 35785 34391 35788
rect 34333 35779 34391 35785
rect 34882 35776 34888 35788
rect 34940 35776 34946 35828
rect 32309 35751 32367 35757
rect 32309 35748 32321 35751
rect 30101 35711 30159 35717
rect 30852 35720 31248 35748
rect 31312 35720 32321 35748
rect 29914 35680 29920 35692
rect 29875 35652 29920 35680
rect 29914 35640 29920 35652
rect 29972 35640 29978 35692
rect 30282 35640 30288 35692
rect 30340 35680 30346 35692
rect 30745 35683 30803 35689
rect 30745 35680 30757 35683
rect 30340 35652 30757 35680
rect 30340 35640 30346 35652
rect 30745 35649 30757 35652
rect 30791 35649 30803 35683
rect 30745 35643 30803 35649
rect 29546 35612 29552 35624
rect 29507 35584 29552 35612
rect 29546 35572 29552 35584
rect 29604 35612 29610 35624
rect 30852 35612 30880 35720
rect 31110 35680 31116 35692
rect 31071 35652 31116 35680
rect 31110 35640 31116 35652
rect 31168 35640 31174 35692
rect 31220 35680 31248 35720
rect 32309 35717 32321 35720
rect 32355 35748 32367 35751
rect 32398 35748 32404 35760
rect 32355 35720 32404 35748
rect 32355 35717 32367 35720
rect 32309 35711 32367 35717
rect 32398 35708 32404 35720
rect 32456 35748 32462 35760
rect 32456 35720 33180 35748
rect 32456 35708 32462 35720
rect 33152 35689 33180 35720
rect 33137 35683 33195 35689
rect 31220 35652 33088 35680
rect 32950 35612 32956 35624
rect 29604 35584 30880 35612
rect 31036 35584 32956 35612
rect 29604 35572 29610 35584
rect 26712 35516 29316 35544
rect 19426 35476 19432 35488
rect 18647 35448 19288 35476
rect 19387 35448 19432 35476
rect 18647 35445 18659 35448
rect 18601 35439 18659 35445
rect 19426 35436 19432 35448
rect 19484 35436 19490 35488
rect 23198 35476 23204 35488
rect 23159 35448 23204 35476
rect 23198 35436 23204 35448
rect 23256 35436 23262 35488
rect 26142 35436 26148 35488
rect 26200 35476 26206 35488
rect 26712 35476 26740 35516
rect 26200 35448 26740 35476
rect 26200 35436 26206 35448
rect 27154 35436 27160 35488
rect 27212 35476 27218 35488
rect 27525 35479 27583 35485
rect 27525 35476 27537 35479
rect 27212 35448 27537 35476
rect 27212 35436 27218 35448
rect 27525 35445 27537 35448
rect 27571 35445 27583 35479
rect 27525 35439 27583 35445
rect 29086 35436 29092 35488
rect 29144 35476 29150 35488
rect 30561 35479 30619 35485
rect 30561 35476 30573 35479
rect 29144 35448 30573 35476
rect 29144 35436 29150 35448
rect 30561 35445 30573 35448
rect 30607 35445 30619 35479
rect 30561 35439 30619 35445
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 31036 35485 31064 35584
rect 32950 35572 32956 35584
rect 33008 35572 33014 35624
rect 33060 35612 33088 35652
rect 33137 35649 33149 35683
rect 33183 35649 33195 35683
rect 33520 35680 33548 35776
rect 36176 35760 36228 35766
rect 33965 35751 34023 35757
rect 33965 35717 33977 35751
rect 34011 35748 34023 35751
rect 34238 35748 34244 35760
rect 34011 35720 34244 35748
rect 34011 35717 34023 35720
rect 33965 35711 34023 35717
rect 34238 35708 34244 35720
rect 34296 35708 34302 35760
rect 36176 35702 36228 35708
rect 34149 35683 34207 35689
rect 34149 35680 34161 35683
rect 33520 35652 34161 35680
rect 33137 35643 33195 35649
rect 34149 35649 34161 35652
rect 34195 35649 34207 35683
rect 34790 35680 34796 35692
rect 34751 35652 34796 35680
rect 34149 35643 34207 35649
rect 34790 35640 34796 35652
rect 34848 35640 34854 35692
rect 35158 35680 35164 35692
rect 35119 35652 35164 35680
rect 35158 35640 35164 35652
rect 35216 35640 35222 35692
rect 35250 35640 35256 35692
rect 35308 35640 35314 35692
rect 34514 35612 34520 35624
rect 33060 35584 34520 35612
rect 34514 35572 34520 35584
rect 34572 35612 34578 35624
rect 35268 35612 35296 35640
rect 34572 35584 35296 35612
rect 34572 35572 34578 35584
rect 35986 35572 35992 35624
rect 36044 35612 36050 35624
rect 36541 35615 36599 35621
rect 36541 35612 36553 35615
rect 36044 35584 36553 35612
rect 36044 35572 36050 35584
rect 36541 35581 36553 35584
rect 36587 35581 36599 35615
rect 36541 35575 36599 35581
rect 31021 35479 31079 35485
rect 31021 35476 31033 35479
rect 30892 35448 31033 35476
rect 30892 35436 30898 35448
rect 31021 35445 31033 35448
rect 31067 35445 31079 35479
rect 32490 35476 32496 35488
rect 32451 35448 32496 35476
rect 31021 35439 31079 35445
rect 32490 35436 32496 35448
rect 32548 35436 32554 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 14090 35232 14096 35284
rect 14148 35272 14154 35284
rect 14553 35275 14611 35281
rect 14553 35272 14565 35275
rect 14148 35244 14565 35272
rect 14148 35232 14154 35244
rect 14553 35241 14565 35244
rect 14599 35241 14611 35275
rect 14553 35235 14611 35241
rect 14737 35275 14795 35281
rect 14737 35241 14749 35275
rect 14783 35272 14795 35275
rect 15010 35272 15016 35284
rect 14783 35244 15016 35272
rect 14783 35241 14795 35244
rect 14737 35235 14795 35241
rect 15010 35232 15016 35244
rect 15068 35232 15074 35284
rect 19518 35272 19524 35284
rect 19479 35244 19524 35272
rect 19518 35232 19524 35244
rect 19576 35232 19582 35284
rect 22738 35232 22744 35284
rect 22796 35272 22802 35284
rect 25593 35275 25651 35281
rect 22796 35244 23065 35272
rect 22796 35232 22802 35244
rect 17681 35207 17739 35213
rect 17681 35204 17693 35207
rect 17236 35176 17693 35204
rect 15657 35139 15715 35145
rect 15657 35105 15669 35139
rect 15703 35136 15715 35139
rect 15746 35136 15752 35148
rect 15703 35108 15752 35136
rect 15703 35105 15715 35108
rect 15657 35099 15715 35105
rect 15746 35096 15752 35108
rect 15804 35136 15810 35148
rect 16853 35139 16911 35145
rect 16853 35136 16865 35139
rect 15804 35108 16865 35136
rect 15804 35096 15810 35108
rect 16853 35105 16865 35108
rect 16899 35105 16911 35139
rect 16853 35099 16911 35105
rect 1857 35071 1915 35077
rect 1857 35037 1869 35071
rect 1903 35068 1915 35071
rect 15562 35068 15568 35080
rect 1903 35040 2084 35068
rect 15523 35040 15568 35068
rect 1903 35037 1915 35040
rect 1857 35031 1915 35037
rect 2056 34944 2084 35040
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 17034 35068 17040 35080
rect 16995 35040 17040 35068
rect 17034 35028 17040 35040
rect 17092 35028 17098 35080
rect 17126 35028 17132 35080
rect 17184 35068 17190 35080
rect 17236 35077 17264 35176
rect 17681 35173 17693 35176
rect 17727 35173 17739 35207
rect 17681 35167 17739 35173
rect 19426 35164 19432 35216
rect 19484 35164 19490 35216
rect 18141 35139 18199 35145
rect 18141 35105 18153 35139
rect 18187 35136 18199 35139
rect 18230 35136 18236 35148
rect 18187 35108 18236 35136
rect 18187 35105 18199 35108
rect 18141 35099 18199 35105
rect 18230 35096 18236 35108
rect 18288 35096 18294 35148
rect 19444 35136 19472 35164
rect 19702 35136 19708 35148
rect 18616 35108 19708 35136
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 17184 35040 17233 35068
rect 17184 35028 17190 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17221 35031 17279 35037
rect 18049 35071 18107 35077
rect 18049 35037 18061 35071
rect 18095 35068 18107 35071
rect 18616 35068 18644 35108
rect 19702 35096 19708 35108
rect 19760 35096 19766 35148
rect 20346 35096 20352 35148
rect 20404 35136 20410 35148
rect 22922 35136 22928 35148
rect 20404 35108 20852 35136
rect 20404 35096 20410 35108
rect 18095 35040 18644 35068
rect 18095 35037 18107 35040
rect 18049 35031 18107 35037
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 19392 35040 19441 35068
rect 19392 35028 19398 35040
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35068 19671 35071
rect 20530 35068 20536 35080
rect 19659 35040 20536 35068
rect 19659 35037 19671 35040
rect 19613 35031 19671 35037
rect 20530 35028 20536 35040
rect 20588 35028 20594 35080
rect 20824 35077 20852 35108
rect 22664 35108 22928 35136
rect 20717 35071 20775 35077
rect 20717 35037 20729 35071
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 20809 35071 20867 35077
rect 20809 35037 20821 35071
rect 20855 35037 20867 35071
rect 20809 35031 20867 35037
rect 14918 35000 14924 35012
rect 14879 34972 14924 35000
rect 14918 34960 14924 34972
rect 14976 35000 14982 35012
rect 15381 35003 15439 35009
rect 15381 35000 15393 35003
rect 14976 34972 15393 35000
rect 14976 34960 14982 34972
rect 15381 34969 15393 34972
rect 15427 34969 15439 35003
rect 20732 35000 20760 35031
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 22664 35077 22692 35108
rect 22922 35096 22928 35108
rect 22980 35096 22986 35148
rect 23037 35136 23065 35244
rect 25593 35241 25605 35275
rect 25639 35272 25651 35275
rect 25866 35272 25872 35284
rect 25639 35244 25872 35272
rect 25639 35241 25651 35244
rect 25593 35235 25651 35241
rect 25866 35232 25872 35244
rect 25924 35232 25930 35284
rect 30834 35272 30840 35284
rect 30795 35244 30840 35272
rect 30834 35232 30840 35244
rect 30892 35232 30898 35284
rect 29362 35164 29368 35216
rect 29420 35204 29426 35216
rect 29420 35176 30052 35204
rect 29420 35164 29426 35176
rect 24946 35136 24952 35148
rect 23032 35108 24952 35136
rect 22649 35071 22707 35077
rect 20956 35040 21001 35068
rect 20956 35028 20962 35040
rect 22649 35037 22661 35071
rect 22695 35037 22707 35071
rect 22830 35068 22836 35080
rect 22791 35040 22836 35068
rect 22649 35031 22707 35037
rect 22830 35028 22836 35040
rect 22888 35028 22894 35080
rect 23032 35077 23060 35108
rect 24946 35096 24952 35108
rect 25004 35096 25010 35148
rect 28810 35136 28816 35148
rect 26252 35108 28816 35136
rect 23017 35071 23075 35077
rect 23017 35037 23029 35071
rect 23063 35037 23075 35071
rect 24762 35068 24768 35080
rect 24723 35040 24768 35068
rect 23017 35031 23075 35037
rect 24762 35028 24768 35040
rect 24820 35028 24826 35080
rect 25038 35068 25044 35080
rect 24999 35040 25044 35068
rect 25038 35028 25044 35040
rect 25096 35028 25102 35080
rect 26252 35077 26280 35108
rect 28810 35096 28816 35108
rect 28868 35136 28874 35148
rect 29454 35136 29460 35148
rect 28868 35108 29460 35136
rect 28868 35096 28874 35108
rect 29454 35096 29460 35108
rect 29512 35096 29518 35148
rect 29822 35136 29828 35148
rect 29783 35108 29828 35136
rect 29822 35096 29828 35108
rect 29880 35096 29886 35148
rect 30024 35145 30052 35176
rect 31772 35176 32076 35204
rect 30009 35139 30067 35145
rect 30009 35105 30021 35139
rect 30055 35105 30067 35139
rect 30009 35099 30067 35105
rect 30098 35096 30104 35148
rect 30156 35136 30162 35148
rect 30156 35108 30201 35136
rect 30156 35096 30162 35108
rect 31018 35096 31024 35148
rect 31076 35136 31082 35148
rect 31478 35136 31484 35148
rect 31076 35108 31484 35136
rect 31076 35096 31082 35108
rect 31478 35096 31484 35108
rect 31536 35136 31542 35148
rect 31772 35136 31800 35176
rect 31536 35108 31800 35136
rect 31536 35096 31542 35108
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35037 26295 35071
rect 26602 35068 26608 35080
rect 26563 35040 26608 35068
rect 26237 35031 26295 35037
rect 26602 35028 26608 35040
rect 26660 35028 26666 35080
rect 27062 35028 27068 35080
rect 27120 35070 27126 35080
rect 28353 35071 28411 35077
rect 27120 35068 27200 35070
rect 27120 35040 28212 35068
rect 27120 35028 27126 35040
rect 22741 35003 22799 35009
rect 20732 34972 22600 35000
rect 15381 34963 15439 34969
rect 1670 34932 1676 34944
rect 1631 34904 1676 34932
rect 1670 34892 1676 34904
rect 1728 34892 1734 34944
rect 2038 34892 2044 34944
rect 2096 34932 2102 34944
rect 2317 34935 2375 34941
rect 2317 34932 2329 34935
rect 2096 34904 2329 34932
rect 2096 34892 2102 34904
rect 2317 34901 2329 34904
rect 2363 34901 2375 34935
rect 2317 34895 2375 34901
rect 14721 34935 14779 34941
rect 14721 34901 14733 34935
rect 14767 34932 14779 34935
rect 15194 34932 15200 34944
rect 14767 34904 15200 34932
rect 14767 34901 14779 34904
rect 14721 34895 14779 34901
rect 15194 34892 15200 34904
rect 15252 34892 15258 34944
rect 15654 34892 15660 34944
rect 15712 34932 15718 34944
rect 15930 34932 15936 34944
rect 15712 34904 15936 34932
rect 15712 34892 15718 34904
rect 15930 34892 15936 34904
rect 15988 34932 15994 34944
rect 16025 34935 16083 34941
rect 16025 34932 16037 34935
rect 15988 34904 16037 34932
rect 15988 34892 15994 34904
rect 16025 34901 16037 34904
rect 16071 34901 16083 34935
rect 16025 34895 16083 34901
rect 21082 34892 21088 34944
rect 21140 34932 21146 34944
rect 21177 34935 21235 34941
rect 21177 34932 21189 34935
rect 21140 34904 21189 34932
rect 21140 34892 21146 34904
rect 21177 34901 21189 34904
rect 21223 34901 21235 34935
rect 21634 34932 21640 34944
rect 21595 34904 21640 34932
rect 21177 34895 21235 34901
rect 21634 34892 21640 34904
rect 21692 34892 21698 34944
rect 21726 34892 21732 34944
rect 21784 34932 21790 34944
rect 22465 34935 22523 34941
rect 22465 34932 22477 34935
rect 21784 34904 22477 34932
rect 21784 34892 21790 34904
rect 22465 34901 22477 34904
rect 22511 34901 22523 34935
rect 22572 34932 22600 34972
rect 22741 34969 22753 35003
rect 22787 35000 22799 35003
rect 23382 35000 23388 35012
rect 22787 34972 23388 35000
rect 22787 34969 22799 34972
rect 22741 34963 22799 34969
rect 23382 34960 23388 34972
rect 23440 35000 23446 35012
rect 24949 35003 25007 35009
rect 24949 35000 24961 35003
rect 23440 34972 24961 35000
rect 23440 34960 23446 34972
rect 24949 34969 24961 34972
rect 24995 35000 25007 35003
rect 25682 35000 25688 35012
rect 24995 34972 25688 35000
rect 24995 34969 25007 34972
rect 24949 34963 25007 34969
rect 25682 34960 25688 34972
rect 25740 34960 25746 35012
rect 26326 35000 26332 35012
rect 26287 34972 26332 35000
rect 26326 34960 26332 34972
rect 26384 34960 26390 35012
rect 26421 35003 26479 35009
rect 26421 34969 26433 35003
rect 26467 35000 26479 35003
rect 26510 35000 26516 35012
rect 26467 34972 26516 35000
rect 26467 34969 26479 34972
rect 26421 34963 26479 34969
rect 26510 34960 26516 34972
rect 26568 35000 26574 35012
rect 27798 35000 27804 35012
rect 26568 34972 27804 35000
rect 26568 34960 26574 34972
rect 27798 34960 27804 34972
rect 27856 35000 27862 35012
rect 28077 35003 28135 35009
rect 28077 35000 28089 35003
rect 27856 34972 28089 35000
rect 27856 34960 27862 34972
rect 28077 34969 28089 34972
rect 28123 34969 28135 35003
rect 28077 34963 28135 34969
rect 23658 34932 23664 34944
rect 22572 34904 23664 34932
rect 22465 34895 22523 34901
rect 23658 34892 23664 34904
rect 23716 34892 23722 34944
rect 24578 34932 24584 34944
rect 24539 34904 24584 34932
rect 24578 34892 24584 34904
rect 24636 34892 24642 34944
rect 26050 34932 26056 34944
rect 26011 34904 26056 34932
rect 26050 34892 26056 34904
rect 26108 34892 26114 34944
rect 27246 34932 27252 34944
rect 27207 34904 27252 34932
rect 27246 34892 27252 34904
rect 27304 34892 27310 34944
rect 28184 34932 28212 35040
rect 28353 35037 28365 35071
rect 28399 35037 28411 35071
rect 28534 35068 28540 35080
rect 28495 35040 28540 35068
rect 28353 35031 28411 35037
rect 28368 35000 28396 35031
rect 28534 35028 28540 35040
rect 28592 35028 28598 35080
rect 28902 35028 28908 35080
rect 28960 35068 28966 35080
rect 29730 35068 29736 35080
rect 28960 35040 29736 35068
rect 28960 35028 28966 35040
rect 29730 35028 29736 35040
rect 29788 35028 29794 35080
rect 29914 35028 29920 35080
rect 29972 35068 29978 35080
rect 30834 35068 30840 35080
rect 29972 35040 30840 35068
rect 29972 35028 29978 35040
rect 30834 35028 30840 35040
rect 30892 35028 30898 35080
rect 31588 35077 31616 35108
rect 31846 35096 31852 35148
rect 31904 35136 31910 35148
rect 32048 35136 32076 35176
rect 33042 35164 33048 35216
rect 33100 35204 33106 35216
rect 33100 35176 34008 35204
rect 33100 35164 33106 35176
rect 33229 35139 33287 35145
rect 33229 35136 33241 35139
rect 31904 35108 31949 35136
rect 32048 35108 33241 35136
rect 31904 35096 31910 35108
rect 33229 35105 33241 35108
rect 33275 35136 33287 35139
rect 33502 35136 33508 35148
rect 33275 35108 33508 35136
rect 33275 35105 33287 35108
rect 33229 35099 33287 35105
rect 33502 35096 33508 35108
rect 33560 35096 33566 35148
rect 31573 35071 31631 35077
rect 31573 35037 31585 35071
rect 31619 35037 31631 35071
rect 31573 35031 31631 35037
rect 31757 35071 31815 35077
rect 31757 35037 31769 35071
rect 31803 35037 31815 35071
rect 31757 35031 31815 35037
rect 28718 35000 28724 35012
rect 28368 34972 28724 35000
rect 28718 34960 28724 34972
rect 28776 35000 28782 35012
rect 29178 35000 29184 35012
rect 28776 34972 29184 35000
rect 28776 34960 28782 34972
rect 29178 34960 29184 34972
rect 29236 34960 29242 35012
rect 30558 35000 30564 35012
rect 30024 34972 30564 35000
rect 28994 34932 29000 34944
rect 28184 34904 29000 34932
rect 28994 34892 29000 34904
rect 29052 34932 29058 34944
rect 30024 34932 30052 34972
rect 30558 34960 30564 34972
rect 30616 34960 30622 35012
rect 30926 34960 30932 35012
rect 30984 35000 30990 35012
rect 31772 35000 31800 35031
rect 31938 35028 31944 35080
rect 31996 35068 32002 35080
rect 31996 35040 32041 35068
rect 31996 35028 32002 35040
rect 32122 35028 32128 35080
rect 32180 35068 32186 35080
rect 32180 35040 32225 35068
rect 32180 35028 32186 35040
rect 32490 35028 32496 35080
rect 32548 35068 32554 35080
rect 33042 35068 33048 35080
rect 32548 35040 33048 35068
rect 32548 35028 32554 35040
rect 33042 35028 33048 35040
rect 33100 35068 33106 35080
rect 33137 35071 33195 35077
rect 33137 35068 33149 35071
rect 33100 35040 33149 35068
rect 33100 35028 33106 35040
rect 33137 35037 33149 35040
rect 33183 35037 33195 35071
rect 33318 35068 33324 35080
rect 33279 35040 33324 35068
rect 33137 35031 33195 35037
rect 33318 35028 33324 35040
rect 33376 35028 33382 35080
rect 33413 35071 33471 35077
rect 33413 35037 33425 35071
rect 33459 35068 33471 35071
rect 33594 35068 33600 35080
rect 33459 35040 33600 35068
rect 33459 35037 33471 35040
rect 33413 35031 33471 35037
rect 30984 34972 31800 35000
rect 30984 34960 30990 34972
rect 31846 34960 31852 35012
rect 31904 35000 31910 35012
rect 33428 35000 33456 35031
rect 33594 35028 33600 35040
rect 33652 35028 33658 35080
rect 33980 35077 34008 35176
rect 34790 35096 34796 35148
rect 34848 35136 34854 35148
rect 35805 35139 35863 35145
rect 35805 35136 35817 35139
rect 34848 35108 35817 35136
rect 34848 35096 34854 35108
rect 35805 35105 35817 35108
rect 35851 35105 35863 35139
rect 35805 35099 35863 35105
rect 33965 35071 34023 35077
rect 33965 35037 33977 35071
rect 34011 35037 34023 35071
rect 33965 35031 34023 35037
rect 34054 35028 34060 35080
rect 34112 35068 34118 35080
rect 34149 35071 34207 35077
rect 34149 35068 34161 35071
rect 34112 35040 34161 35068
rect 34112 35028 34118 35040
rect 34149 35037 34161 35040
rect 34195 35037 34207 35071
rect 34149 35031 34207 35037
rect 36081 35071 36139 35077
rect 36081 35037 36093 35071
rect 36127 35068 36139 35071
rect 36127 35040 36676 35068
rect 36127 35037 36139 35040
rect 36081 35031 36139 35037
rect 31904 34972 33456 35000
rect 31904 34960 31910 34972
rect 29052 34904 30052 34932
rect 30285 34935 30343 34941
rect 29052 34892 29058 34904
rect 30285 34901 30297 34935
rect 30331 34932 30343 34935
rect 31110 34932 31116 34944
rect 30331 34904 31116 34932
rect 30331 34901 30343 34904
rect 30285 34895 30343 34901
rect 31110 34892 31116 34904
rect 31168 34892 31174 34944
rect 31389 34935 31447 34941
rect 31389 34901 31401 34935
rect 31435 34932 31447 34935
rect 31570 34932 31576 34944
rect 31435 34904 31576 34932
rect 31435 34901 31447 34904
rect 31389 34895 31447 34901
rect 31570 34892 31576 34904
rect 31628 34892 31634 34944
rect 32674 34892 32680 34944
rect 32732 34932 32738 34944
rect 32953 34935 33011 34941
rect 32953 34932 32965 34935
rect 32732 34904 32965 34932
rect 32732 34892 32738 34904
rect 32953 34901 32965 34904
rect 32999 34901 33011 34935
rect 32953 34895 33011 34901
rect 33134 34892 33140 34944
rect 33192 34932 33198 34944
rect 33318 34932 33324 34944
rect 33192 34904 33324 34932
rect 33192 34892 33198 34904
rect 33318 34892 33324 34904
rect 33376 34892 33382 34944
rect 33410 34892 33416 34944
rect 33468 34932 33474 34944
rect 36648 34941 36676 35040
rect 34057 34935 34115 34941
rect 34057 34932 34069 34935
rect 33468 34904 34069 34932
rect 33468 34892 33474 34904
rect 34057 34901 34069 34904
rect 34103 34901 34115 34935
rect 34057 34895 34115 34901
rect 36633 34935 36691 34941
rect 36633 34901 36645 34935
rect 36679 34932 36691 34935
rect 36906 34932 36912 34944
rect 36679 34904 36912 34932
rect 36679 34901 36691 34904
rect 36633 34895 36691 34901
rect 36906 34892 36912 34904
rect 36964 34892 36970 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 14918 34688 14924 34740
rect 14976 34728 14982 34740
rect 15473 34731 15531 34737
rect 15473 34728 15485 34731
rect 14976 34700 15485 34728
rect 14976 34688 14982 34700
rect 15473 34697 15485 34700
rect 15519 34697 15531 34731
rect 18230 34728 18236 34740
rect 18191 34700 18236 34728
rect 15473 34691 15531 34697
rect 18230 34688 18236 34700
rect 18288 34688 18294 34740
rect 20898 34688 20904 34740
rect 20956 34728 20962 34740
rect 20956 34700 22508 34728
rect 20956 34688 20962 34700
rect 15194 34660 15200 34672
rect 15028 34632 15200 34660
rect 15028 34533 15056 34632
rect 15194 34620 15200 34632
rect 15252 34620 15258 34672
rect 18506 34620 18512 34672
rect 18564 34660 18570 34672
rect 18601 34663 18659 34669
rect 18601 34660 18613 34663
rect 18564 34632 18613 34660
rect 18564 34620 18570 34632
rect 18601 34629 18613 34632
rect 18647 34660 18659 34663
rect 18782 34660 18788 34672
rect 18647 34632 18788 34660
rect 18647 34629 18659 34632
rect 18601 34623 18659 34629
rect 18782 34620 18788 34632
rect 18840 34620 18846 34672
rect 19797 34663 19855 34669
rect 19797 34629 19809 34663
rect 19843 34660 19855 34663
rect 20070 34660 20076 34672
rect 19843 34632 20076 34660
rect 19843 34629 19855 34632
rect 19797 34623 19855 34629
rect 20070 34620 20076 34632
rect 20128 34660 20134 34672
rect 22370 34660 22376 34672
rect 20128 34632 22376 34660
rect 20128 34620 20134 34632
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 22480 34660 22508 34700
rect 22554 34688 22560 34740
rect 22612 34728 22618 34740
rect 22925 34731 22983 34737
rect 22925 34728 22937 34731
rect 22612 34700 22937 34728
rect 22612 34688 22618 34700
rect 22925 34697 22937 34700
rect 22971 34728 22983 34731
rect 23014 34728 23020 34740
rect 22971 34700 23020 34728
rect 22971 34697 22983 34700
rect 22925 34691 22983 34697
rect 23014 34688 23020 34700
rect 23072 34688 23078 34740
rect 24857 34731 24915 34737
rect 23124 34700 24808 34728
rect 23124 34660 23152 34700
rect 22480 34632 23152 34660
rect 23198 34620 23204 34672
rect 23256 34660 23262 34672
rect 23256 34632 23612 34660
rect 23256 34620 23262 34632
rect 18417 34595 18475 34601
rect 18417 34561 18429 34595
rect 18463 34561 18475 34595
rect 18417 34555 18475 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34592 21051 34595
rect 21726 34592 21732 34604
rect 21039 34564 21732 34592
rect 21039 34561 21051 34564
rect 20993 34555 21051 34561
rect 15013 34527 15071 34533
rect 15013 34493 15025 34527
rect 15059 34493 15071 34527
rect 15013 34487 15071 34493
rect 15102 34484 15108 34536
rect 15160 34524 15166 34536
rect 18432 34524 18460 34555
rect 21726 34552 21732 34564
rect 21784 34552 21790 34604
rect 22465 34595 22523 34601
rect 22465 34561 22477 34595
rect 22511 34592 22523 34595
rect 23385 34595 23443 34601
rect 23385 34592 23397 34595
rect 22511 34564 23397 34592
rect 22511 34561 22523 34564
rect 22465 34555 22523 34561
rect 23385 34561 23397 34564
rect 23431 34592 23443 34595
rect 23474 34592 23480 34604
rect 23431 34564 23480 34592
rect 23431 34561 23443 34564
rect 23385 34555 23443 34561
rect 23474 34552 23480 34564
rect 23532 34552 23538 34604
rect 23584 34601 23612 34632
rect 23569 34595 23627 34601
rect 23569 34561 23581 34595
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 23658 34552 23664 34604
rect 23716 34592 23722 34604
rect 24780 34601 24808 34700
rect 24857 34697 24869 34731
rect 24903 34728 24915 34731
rect 24946 34728 24952 34740
rect 24903 34700 24952 34728
rect 24903 34697 24915 34700
rect 24857 34691 24915 34697
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 25038 34688 25044 34740
rect 25096 34728 25102 34740
rect 25096 34700 28028 34728
rect 25096 34688 25102 34700
rect 25222 34660 25228 34672
rect 24964 34632 25228 34660
rect 24964 34601 24992 34632
rect 25222 34620 25228 34632
rect 25280 34660 25286 34672
rect 26050 34660 26056 34672
rect 25280 34632 26056 34660
rect 25280 34620 25286 34632
rect 26050 34620 26056 34632
rect 26108 34620 26114 34672
rect 26605 34663 26663 34669
rect 26605 34629 26617 34663
rect 26651 34660 26663 34663
rect 26786 34660 26792 34672
rect 26651 34632 26792 34660
rect 26651 34629 26663 34632
rect 26605 34623 26663 34629
rect 26786 34620 26792 34632
rect 26844 34620 26850 34672
rect 27157 34663 27215 34669
rect 27157 34629 27169 34663
rect 27203 34660 27215 34663
rect 27614 34660 27620 34672
rect 27203 34632 27620 34660
rect 27203 34629 27215 34632
rect 27157 34623 27215 34629
rect 27614 34620 27620 34632
rect 27672 34620 27678 34672
rect 27890 34660 27896 34672
rect 27851 34632 27896 34660
rect 27890 34620 27896 34632
rect 27948 34620 27954 34672
rect 28000 34660 28028 34700
rect 28994 34688 29000 34740
rect 29052 34728 29058 34740
rect 29089 34731 29147 34737
rect 29089 34728 29101 34731
rect 29052 34700 29101 34728
rect 29052 34688 29058 34700
rect 29089 34697 29101 34700
rect 29135 34697 29147 34731
rect 29089 34691 29147 34697
rect 29472 34700 31754 34728
rect 29472 34660 29500 34700
rect 28000 34632 29500 34660
rect 29822 34620 29828 34672
rect 29880 34660 29886 34672
rect 29880 34632 30052 34660
rect 29880 34620 29886 34632
rect 24765 34595 24823 34601
rect 23716 34564 23761 34592
rect 23716 34552 23722 34564
rect 24765 34561 24777 34595
rect 24811 34561 24823 34595
rect 24765 34555 24823 34561
rect 24949 34595 25007 34601
rect 24949 34561 24961 34595
rect 24995 34561 25007 34595
rect 25590 34592 25596 34604
rect 25551 34564 25596 34592
rect 24949 34555 25007 34561
rect 19153 34527 19211 34533
rect 19153 34524 19165 34527
rect 15160 34496 15205 34524
rect 18432 34496 19165 34524
rect 15160 34484 15166 34496
rect 19153 34493 19165 34496
rect 19199 34524 19211 34527
rect 19242 34524 19248 34536
rect 19199 34496 19248 34524
rect 19199 34493 19211 34496
rect 19153 34487 19211 34493
rect 19242 34484 19248 34496
rect 19300 34484 19306 34536
rect 21082 34524 21088 34536
rect 21043 34496 21088 34524
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 22002 34484 22008 34536
rect 22060 34524 22066 34536
rect 22281 34527 22339 34533
rect 22281 34524 22293 34527
rect 22060 34496 22293 34524
rect 22060 34484 22066 34496
rect 22281 34493 22293 34496
rect 22327 34493 22339 34527
rect 22281 34487 22339 34493
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34524 22615 34527
rect 22646 34524 22652 34536
rect 22603 34496 22652 34524
rect 22603 34493 22615 34496
rect 22557 34487 22615 34493
rect 22646 34484 22652 34496
rect 22704 34484 22710 34536
rect 24780 34524 24808 34555
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 27246 34552 27252 34604
rect 27304 34592 27310 34604
rect 27709 34595 27767 34601
rect 27709 34592 27721 34595
rect 27304 34564 27721 34592
rect 27304 34552 27310 34564
rect 27709 34561 27721 34564
rect 27755 34561 27767 34595
rect 27709 34555 27767 34561
rect 25498 34524 25504 34536
rect 24780 34496 25504 34524
rect 25498 34484 25504 34496
rect 25556 34484 25562 34536
rect 25777 34527 25835 34533
rect 25777 34493 25789 34527
rect 25823 34524 25835 34527
rect 26418 34524 26424 34536
rect 25823 34496 26424 34524
rect 25823 34493 25835 34496
rect 25777 34487 25835 34493
rect 26418 34484 26424 34496
rect 26476 34484 26482 34536
rect 27724 34524 27752 34555
rect 27798 34552 27804 34604
rect 27856 34592 27862 34604
rect 27985 34595 28043 34601
rect 27985 34592 27997 34595
rect 27856 34564 27997 34592
rect 27856 34552 27862 34564
rect 27985 34561 27997 34564
rect 28031 34561 28043 34595
rect 27985 34555 28043 34561
rect 28074 34552 28080 34604
rect 28132 34592 28138 34604
rect 28810 34592 28816 34604
rect 28132 34564 28177 34592
rect 28771 34564 28816 34592
rect 28132 34552 28138 34564
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 29270 34552 29276 34604
rect 29328 34592 29334 34604
rect 29641 34595 29699 34601
rect 29641 34592 29653 34595
rect 29328 34564 29653 34592
rect 29328 34552 29334 34564
rect 29641 34561 29653 34564
rect 29687 34561 29699 34595
rect 29641 34555 29699 34561
rect 29730 34552 29736 34604
rect 29788 34592 29794 34604
rect 30024 34601 30052 34632
rect 30852 34632 31248 34660
rect 30009 34595 30067 34601
rect 29788 34564 29833 34592
rect 29788 34552 29794 34564
rect 30009 34561 30021 34595
rect 30055 34561 30067 34595
rect 30009 34555 30067 34561
rect 30190 34552 30196 34604
rect 30248 34592 30254 34604
rect 30852 34601 30880 34632
rect 30837 34595 30895 34601
rect 30837 34592 30849 34595
rect 30248 34564 30849 34592
rect 30248 34552 30254 34564
rect 30837 34561 30849 34564
rect 30883 34561 30895 34595
rect 31110 34592 31116 34604
rect 31071 34564 31116 34592
rect 30837 34555 30895 34561
rect 31110 34552 31116 34564
rect 31168 34552 31174 34604
rect 29825 34527 29883 34533
rect 29825 34524 29837 34527
rect 27724 34496 29837 34524
rect 29825 34493 29837 34496
rect 29871 34524 29883 34527
rect 29914 34524 29920 34536
rect 29871 34496 29920 34524
rect 29871 34493 29883 34496
rect 29825 34487 29883 34493
rect 29914 34484 29920 34496
rect 29972 34484 29978 34536
rect 30650 34524 30656 34536
rect 30611 34496 30656 34524
rect 30650 34484 30656 34496
rect 30708 34484 30714 34536
rect 30926 34524 30932 34536
rect 30887 34496 30932 34524
rect 30926 34484 30932 34496
rect 30984 34484 30990 34536
rect 31018 34484 31024 34536
rect 31076 34524 31082 34536
rect 31220 34524 31248 34632
rect 31726 34592 31754 34700
rect 57882 34688 57888 34740
rect 57940 34728 57946 34740
rect 58253 34731 58311 34737
rect 58253 34728 58265 34731
rect 57940 34700 58265 34728
rect 57940 34688 57946 34700
rect 58253 34697 58265 34700
rect 58299 34697 58311 34731
rect 58253 34691 58311 34697
rect 33045 34663 33103 34669
rect 33045 34629 33057 34663
rect 33091 34660 33103 34663
rect 33134 34660 33140 34672
rect 33091 34632 33140 34660
rect 33091 34629 33103 34632
rect 33045 34623 33103 34629
rect 33134 34620 33140 34632
rect 33192 34660 33198 34672
rect 34054 34660 34060 34672
rect 33192 34632 34060 34660
rect 33192 34620 33198 34632
rect 34054 34620 34060 34632
rect 34112 34660 34118 34672
rect 34517 34663 34575 34669
rect 34517 34660 34529 34663
rect 34112 34632 34529 34660
rect 34112 34620 34118 34632
rect 34517 34629 34529 34632
rect 34563 34629 34575 34663
rect 34517 34623 34575 34629
rect 32309 34595 32367 34601
rect 32309 34592 32321 34595
rect 31726 34564 32321 34592
rect 32309 34561 32321 34564
rect 32355 34561 32367 34595
rect 32309 34555 32367 34561
rect 33318 34552 33324 34604
rect 33376 34592 33382 34604
rect 33686 34592 33692 34604
rect 33376 34564 33692 34592
rect 33376 34552 33382 34564
rect 33686 34552 33692 34564
rect 33744 34592 33750 34604
rect 33870 34592 33876 34604
rect 33744 34564 33876 34592
rect 33744 34552 33750 34564
rect 33870 34552 33876 34564
rect 33928 34552 33934 34604
rect 35526 34592 35532 34604
rect 35487 34564 35532 34592
rect 35526 34552 35532 34564
rect 35584 34552 35590 34604
rect 35710 34592 35716 34604
rect 35671 34564 35716 34592
rect 35710 34552 35716 34564
rect 35768 34552 35774 34604
rect 36541 34595 36599 34601
rect 36541 34561 36553 34595
rect 36587 34561 36599 34595
rect 36541 34555 36599 34561
rect 31386 34524 31392 34536
rect 31076 34496 31121 34524
rect 31220 34496 31392 34524
rect 31076 34484 31082 34496
rect 31386 34484 31392 34496
rect 31444 34524 31450 34536
rect 31665 34527 31723 34533
rect 31665 34524 31677 34527
rect 31444 34496 31677 34524
rect 31444 34484 31450 34496
rect 31665 34493 31677 34496
rect 31711 34493 31723 34527
rect 31665 34487 31723 34493
rect 31938 34484 31944 34536
rect 31996 34524 32002 34536
rect 32401 34527 32459 34533
rect 32401 34524 32413 34527
rect 31996 34496 32413 34524
rect 31996 34484 32002 34496
rect 32401 34493 32413 34496
rect 32447 34493 32459 34527
rect 33962 34524 33968 34536
rect 33923 34496 33968 34524
rect 32401 34487 32459 34493
rect 33962 34484 33968 34496
rect 34020 34484 34026 34536
rect 35544 34524 35572 34552
rect 36556 34524 36584 34555
rect 37458 34552 37464 34604
rect 37516 34592 37522 34604
rect 37645 34595 37703 34601
rect 37645 34592 37657 34595
rect 37516 34564 37657 34592
rect 37516 34552 37522 34564
rect 37645 34561 37657 34564
rect 37691 34561 37703 34595
rect 58069 34595 58127 34601
rect 58069 34592 58081 34595
rect 37645 34555 37703 34561
rect 57440 34564 58081 34592
rect 57440 34536 57468 34564
rect 58069 34561 58081 34564
rect 58115 34561 58127 34595
rect 58069 34555 58127 34561
rect 35544 34496 36584 34524
rect 36633 34527 36691 34533
rect 36633 34493 36645 34527
rect 36679 34524 36691 34527
rect 36722 34524 36728 34536
rect 36679 34496 36728 34524
rect 36679 34493 36691 34496
rect 36633 34487 36691 34493
rect 36722 34484 36728 34496
rect 36780 34484 36786 34536
rect 36909 34527 36967 34533
rect 36909 34493 36921 34527
rect 36955 34524 36967 34527
rect 37553 34527 37611 34533
rect 37553 34524 37565 34527
rect 36955 34496 37565 34524
rect 36955 34493 36967 34496
rect 36909 34487 36967 34493
rect 37553 34493 37565 34496
rect 37599 34493 37611 34527
rect 57422 34524 57428 34536
rect 57383 34496 57428 34524
rect 37553 34487 37611 34493
rect 57422 34484 57428 34496
rect 57480 34484 57486 34536
rect 21361 34459 21419 34465
rect 21361 34425 21373 34459
rect 21407 34456 21419 34459
rect 21726 34456 21732 34468
rect 21407 34428 21732 34456
rect 21407 34425 21419 34428
rect 21361 34419 21419 34425
rect 21726 34416 21732 34428
rect 21784 34416 21790 34468
rect 22738 34416 22744 34468
rect 22796 34456 22802 34468
rect 26786 34456 26792 34468
rect 22796 34428 26792 34456
rect 22796 34416 22802 34428
rect 26786 34416 26792 34428
rect 26844 34416 26850 34468
rect 33042 34416 33048 34468
rect 33100 34456 33106 34468
rect 33505 34459 33563 34465
rect 33505 34456 33517 34459
rect 33100 34428 33517 34456
rect 33100 34416 33106 34428
rect 33505 34425 33517 34428
rect 33551 34425 33563 34459
rect 33505 34419 33563 34425
rect 38013 34459 38071 34465
rect 38013 34425 38025 34459
rect 38059 34456 38071 34459
rect 38930 34456 38936 34468
rect 38059 34428 38936 34456
rect 38059 34425 38071 34428
rect 38013 34419 38071 34425
rect 38930 34416 38936 34428
rect 38988 34416 38994 34468
rect 14829 34391 14887 34397
rect 14829 34357 14841 34391
rect 14875 34388 14887 34391
rect 15378 34388 15384 34400
rect 14875 34360 15384 34388
rect 14875 34357 14887 34360
rect 14829 34351 14887 34357
rect 15378 34348 15384 34360
rect 15436 34348 15442 34400
rect 20346 34388 20352 34400
rect 20307 34360 20352 34388
rect 20346 34348 20352 34360
rect 20404 34348 20410 34400
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 27982 34388 27988 34400
rect 21140 34360 27988 34388
rect 21140 34348 21146 34360
rect 27982 34348 27988 34360
rect 28040 34348 28046 34400
rect 28258 34388 28264 34400
rect 28219 34360 28264 34388
rect 28258 34348 28264 34360
rect 28316 34348 28322 34400
rect 28994 34348 29000 34400
rect 29052 34388 29058 34400
rect 30009 34391 30067 34397
rect 30009 34388 30021 34391
rect 29052 34360 30021 34388
rect 29052 34348 29058 34360
rect 30009 34357 30021 34360
rect 30055 34357 30067 34391
rect 35618 34388 35624 34400
rect 35579 34360 35624 34388
rect 30009 34351 30067 34357
rect 35618 34348 35624 34360
rect 35676 34348 35682 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 15654 34184 15660 34196
rect 15615 34156 15660 34184
rect 15654 34144 15660 34156
rect 15712 34144 15718 34196
rect 20346 34144 20352 34196
rect 20404 34184 20410 34196
rect 20901 34187 20959 34193
rect 20901 34184 20913 34187
rect 20404 34156 20913 34184
rect 20404 34144 20410 34156
rect 20901 34153 20913 34156
rect 20947 34184 20959 34187
rect 21450 34184 21456 34196
rect 20947 34156 21456 34184
rect 20947 34153 20959 34156
rect 20901 34147 20959 34153
rect 21450 34144 21456 34156
rect 21508 34144 21514 34196
rect 23566 34184 23572 34196
rect 23527 34156 23572 34184
rect 23566 34144 23572 34156
rect 23624 34144 23630 34196
rect 30653 34187 30711 34193
rect 24688 34156 28994 34184
rect 17402 34116 17408 34128
rect 17363 34088 17408 34116
rect 17402 34076 17408 34088
rect 17460 34076 17466 34128
rect 18506 34116 18512 34128
rect 17604 34088 18512 34116
rect 15381 34051 15439 34057
rect 15381 34017 15393 34051
rect 15427 34048 15439 34051
rect 16206 34048 16212 34060
rect 15427 34020 16212 34048
rect 15427 34017 15439 34020
rect 15381 34011 15439 34017
rect 16206 34008 16212 34020
rect 16264 34008 16270 34060
rect 15286 33980 15292 33992
rect 15247 33952 15292 33980
rect 15286 33940 15292 33952
rect 15344 33940 15350 33992
rect 17604 33989 17632 34088
rect 18506 34076 18512 34088
rect 18564 34076 18570 34128
rect 20364 34116 20392 34144
rect 20088 34088 20392 34116
rect 23385 34119 23443 34125
rect 18417 34051 18475 34057
rect 18417 34048 18429 34051
rect 17696 34020 18429 34048
rect 17696 33989 17724 34020
rect 18417 34017 18429 34020
rect 18463 34048 18475 34051
rect 19426 34048 19432 34060
rect 18463 34020 19432 34048
rect 18463 34017 18475 34020
rect 18417 34011 18475 34017
rect 19426 34008 19432 34020
rect 19484 34008 19490 34060
rect 20088 34057 20116 34088
rect 23385 34085 23397 34119
rect 23431 34116 23443 34119
rect 23474 34116 23480 34128
rect 23431 34088 23480 34116
rect 23431 34085 23443 34088
rect 23385 34079 23443 34085
rect 23474 34076 23480 34088
rect 23532 34076 23538 34128
rect 20073 34051 20131 34057
rect 20073 34017 20085 34051
rect 20119 34017 20131 34051
rect 20073 34011 20131 34017
rect 20349 34051 20407 34057
rect 20349 34017 20361 34051
rect 20395 34048 20407 34051
rect 20530 34048 20536 34060
rect 20395 34020 20536 34048
rect 20395 34017 20407 34020
rect 20349 34011 20407 34017
rect 20530 34008 20536 34020
rect 20588 34008 20594 34060
rect 20809 34051 20867 34057
rect 20809 34017 20821 34051
rect 20855 34048 20867 34051
rect 22281 34051 22339 34057
rect 20855 34020 21680 34048
rect 20855 34017 20867 34020
rect 20809 34011 20867 34017
rect 21652 33992 21680 34020
rect 22281 34017 22293 34051
rect 22327 34048 22339 34051
rect 24688 34048 24716 34156
rect 28966 34116 28994 34156
rect 30653 34153 30665 34187
rect 30699 34184 30711 34187
rect 33781 34187 33839 34193
rect 30699 34156 33732 34184
rect 30699 34153 30711 34156
rect 30653 34147 30711 34153
rect 29181 34119 29239 34125
rect 28966 34088 29132 34116
rect 22327 34020 24716 34048
rect 24765 34051 24823 34057
rect 22327 34017 22339 34020
rect 22281 34011 22339 34017
rect 24765 34017 24777 34051
rect 24811 34048 24823 34051
rect 24946 34048 24952 34060
rect 24811 34020 24952 34048
rect 24811 34017 24823 34020
rect 24765 34011 24823 34017
rect 24946 34008 24952 34020
rect 25004 34008 25010 34060
rect 25222 34048 25228 34060
rect 25183 34020 25228 34048
rect 25222 34008 25228 34020
rect 25280 34008 25286 34060
rect 25777 34051 25835 34057
rect 25777 34017 25789 34051
rect 25823 34048 25835 34051
rect 27154 34048 27160 34060
rect 25823 34020 27160 34048
rect 25823 34017 25835 34020
rect 25777 34011 25835 34017
rect 27154 34008 27160 34020
rect 27212 34008 27218 34060
rect 27522 34048 27528 34060
rect 27483 34020 27528 34048
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 27706 34048 27712 34060
rect 27667 34020 27712 34048
rect 27706 34008 27712 34020
rect 27764 34008 27770 34060
rect 28629 34051 28687 34057
rect 28629 34017 28641 34051
rect 28675 34048 28687 34051
rect 28994 34048 29000 34060
rect 28675 34020 29000 34048
rect 28675 34017 28687 34020
rect 28629 34011 28687 34017
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 29104 34048 29132 34088
rect 29181 34085 29193 34119
rect 29227 34116 29239 34119
rect 31018 34116 31024 34128
rect 29227 34088 31024 34116
rect 29227 34085 29239 34088
rect 29181 34079 29239 34085
rect 31018 34076 31024 34088
rect 31076 34076 31082 34128
rect 31110 34076 31116 34128
rect 31168 34116 31174 34128
rect 32122 34116 32128 34128
rect 31168 34088 32128 34116
rect 31168 34076 31174 34088
rect 32122 34076 32128 34088
rect 32180 34116 32186 34128
rect 32585 34119 32643 34125
rect 32180 34088 32444 34116
rect 32180 34076 32186 34088
rect 29104 34020 29776 34048
rect 17589 33983 17647 33989
rect 17589 33949 17601 33983
rect 17635 33949 17647 33983
rect 17589 33943 17647 33949
rect 17681 33983 17739 33989
rect 17681 33949 17693 33983
rect 17727 33949 17739 33983
rect 18322 33980 18328 33992
rect 18283 33952 18328 33980
rect 17681 33943 17739 33949
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 18506 33980 18512 33992
rect 18467 33952 18512 33980
rect 18506 33940 18512 33952
rect 18564 33940 18570 33992
rect 18598 33940 18604 33992
rect 18656 33980 18662 33992
rect 19978 33980 19984 33992
rect 18656 33952 18701 33980
rect 19939 33952 19984 33980
rect 18656 33940 18662 33952
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 21085 33983 21143 33989
rect 21085 33949 21097 33983
rect 21131 33949 21143 33983
rect 21085 33943 21143 33949
rect 17405 33915 17463 33921
rect 17405 33881 17417 33915
rect 17451 33912 17463 33915
rect 18616 33912 18644 33940
rect 17451 33884 18644 33912
rect 19996 33912 20024 33940
rect 21100 33912 21128 33943
rect 21634 33940 21640 33992
rect 21692 33980 21698 33992
rect 21729 33983 21787 33989
rect 21729 33980 21741 33983
rect 21692 33952 21741 33980
rect 21692 33940 21698 33952
rect 21729 33949 21741 33952
rect 21775 33980 21787 33983
rect 22738 33980 22744 33992
rect 21775 33952 22744 33980
rect 21775 33949 21787 33952
rect 21729 33943 21787 33949
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 23014 33940 23020 33992
rect 23072 33980 23078 33992
rect 24857 33983 24915 33989
rect 24857 33980 24869 33983
rect 23072 33952 24869 33980
rect 23072 33940 23078 33952
rect 24780 33924 24808 33952
rect 24857 33949 24869 33952
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 25958 33940 25964 33992
rect 26016 33980 26022 33992
rect 26145 33983 26203 33989
rect 26145 33980 26157 33983
rect 26016 33952 26157 33980
rect 26016 33940 26022 33952
rect 26145 33949 26157 33952
rect 26191 33949 26203 33983
rect 26145 33943 26203 33949
rect 26237 33983 26295 33989
rect 26237 33949 26249 33983
rect 26283 33980 26295 33983
rect 26602 33980 26608 33992
rect 26283 33952 26608 33980
rect 26283 33949 26295 33952
rect 26237 33943 26295 33949
rect 26602 33940 26608 33952
rect 26660 33940 26666 33992
rect 26970 33940 26976 33992
rect 27028 33980 27034 33992
rect 27433 33983 27491 33989
rect 27433 33980 27445 33983
rect 27028 33952 27445 33980
rect 27028 33940 27034 33952
rect 27433 33949 27445 33952
rect 27479 33949 27491 33983
rect 27433 33943 27491 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33980 27675 33983
rect 29086 33980 29092 33992
rect 27663 33952 29092 33980
rect 27663 33949 27675 33952
rect 27617 33943 27675 33949
rect 29086 33940 29092 33952
rect 29144 33940 29150 33992
rect 29748 33980 29776 34020
rect 29822 34008 29828 34060
rect 29880 34048 29886 34060
rect 30009 34051 30067 34057
rect 30009 34048 30021 34051
rect 29880 34020 30021 34048
rect 29880 34008 29886 34020
rect 30009 34017 30021 34020
rect 30055 34017 30067 34051
rect 30009 34011 30067 34017
rect 30926 34008 30932 34060
rect 30984 34048 30990 34060
rect 31389 34051 31447 34057
rect 31389 34048 31401 34051
rect 30984 34020 31401 34048
rect 30984 34008 30990 34020
rect 31110 33980 31116 33992
rect 29748 33952 31116 33980
rect 31110 33940 31116 33952
rect 31168 33940 31174 33992
rect 19996 33884 21404 33912
rect 17451 33881 17463 33884
rect 17405 33875 17463 33881
rect 17954 33804 17960 33856
rect 18012 33844 18018 33856
rect 18141 33847 18199 33853
rect 18141 33844 18153 33847
rect 18012 33816 18153 33844
rect 18012 33804 18018 33816
rect 18141 33813 18153 33816
rect 18187 33813 18199 33847
rect 18141 33807 18199 33813
rect 18322 33804 18328 33856
rect 18380 33844 18386 33856
rect 20254 33844 20260 33856
rect 18380 33816 20260 33844
rect 18380 33804 18386 33816
rect 20254 33804 20260 33816
rect 20312 33804 20318 33856
rect 21266 33844 21272 33856
rect 21227 33816 21272 33844
rect 21266 33804 21272 33816
rect 21324 33804 21330 33856
rect 21376 33844 21404 33884
rect 21450 33872 21456 33924
rect 21508 33912 21514 33924
rect 21508 33884 22048 33912
rect 21508 33872 21514 33884
rect 22020 33853 22048 33884
rect 22094 33872 22100 33924
rect 22152 33912 22158 33924
rect 23750 33912 23756 33924
rect 22152 33884 22197 33912
rect 23711 33884 23756 33912
rect 22152 33872 22158 33884
rect 23750 33872 23756 33884
rect 23808 33872 23814 33924
rect 24762 33872 24768 33924
rect 24820 33872 24826 33924
rect 25682 33872 25688 33924
rect 25740 33912 25746 33924
rect 26421 33915 26479 33921
rect 25740 33884 26096 33912
rect 25740 33872 25746 33884
rect 21913 33847 21971 33853
rect 21913 33844 21925 33847
rect 21376 33816 21925 33844
rect 21913 33813 21925 33816
rect 21959 33813 21971 33847
rect 21913 33807 21971 33813
rect 22005 33847 22063 33853
rect 22005 33813 22017 33847
rect 22051 33844 22063 33847
rect 22186 33844 22192 33856
rect 22051 33816 22192 33844
rect 22051 33813 22063 33816
rect 22005 33807 22063 33813
rect 22186 33804 22192 33816
rect 22244 33804 22250 33856
rect 23553 33847 23611 33853
rect 23553 33813 23565 33847
rect 23599 33844 23611 33847
rect 24026 33844 24032 33856
rect 23599 33816 24032 33844
rect 23599 33813 23611 33816
rect 23553 33807 23611 33813
rect 24026 33804 24032 33816
rect 24084 33804 24090 33856
rect 24581 33847 24639 33853
rect 24581 33813 24593 33847
rect 24627 33844 24639 33847
rect 24670 33844 24676 33856
rect 24627 33816 24676 33844
rect 24627 33813 24639 33816
rect 24581 33807 24639 33813
rect 24670 33804 24676 33816
rect 24728 33804 24734 33856
rect 24946 33844 24952 33856
rect 24907 33816 24952 33844
rect 24946 33804 24952 33816
rect 25004 33804 25010 33856
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 25133 33847 25191 33853
rect 25133 33844 25145 33847
rect 25096 33816 25145 33844
rect 25096 33804 25102 33816
rect 25133 33813 25145 33816
rect 25179 33813 25191 33847
rect 25133 33807 25191 33813
rect 25774 33804 25780 33856
rect 25832 33844 25838 33856
rect 26068 33853 26096 33884
rect 26421 33881 26433 33915
rect 26467 33912 26479 33915
rect 28813 33915 28871 33921
rect 28813 33912 28825 33915
rect 26467 33884 28825 33912
rect 26467 33881 26479 33884
rect 26421 33875 26479 33881
rect 28813 33881 28825 33884
rect 28859 33881 28871 33915
rect 28813 33875 28871 33881
rect 30285 33915 30343 33921
rect 30285 33881 30297 33915
rect 30331 33912 30343 33915
rect 30331 33884 31156 33912
rect 30331 33881 30343 33884
rect 30285 33875 30343 33881
rect 25869 33847 25927 33853
rect 25869 33844 25881 33847
rect 25832 33816 25881 33844
rect 25832 33804 25838 33816
rect 25869 33813 25881 33816
rect 25915 33813 25927 33847
rect 25869 33807 25927 33813
rect 26053 33847 26111 33853
rect 26053 33813 26065 33847
rect 26099 33844 26111 33847
rect 27430 33844 27436 33856
rect 26099 33816 27436 33844
rect 26099 33813 26111 33816
rect 26053 33807 26111 33813
rect 27430 33804 27436 33816
rect 27488 33804 27494 33856
rect 27893 33847 27951 33853
rect 27893 33813 27905 33847
rect 27939 33844 27951 33847
rect 28442 33844 28448 33856
rect 27939 33816 28448 33844
rect 27939 33813 27951 33816
rect 27893 33807 27951 33813
rect 28442 33804 28448 33816
rect 28500 33804 28506 33856
rect 28718 33844 28724 33856
rect 28679 33816 28724 33844
rect 28718 33804 28724 33816
rect 28776 33804 28782 33856
rect 30193 33847 30251 33853
rect 30193 33813 30205 33847
rect 30239 33844 30251 33847
rect 30558 33844 30564 33856
rect 30239 33816 30564 33844
rect 30239 33813 30251 33816
rect 30193 33807 30251 33813
rect 30558 33804 30564 33816
rect 30616 33804 30622 33856
rect 31128 33853 31156 33884
rect 31113 33847 31171 33853
rect 31113 33813 31125 33847
rect 31159 33813 31171 33847
rect 31220 33844 31248 34020
rect 31389 34017 31401 34020
rect 31435 34017 31447 34051
rect 31389 34011 31447 34017
rect 31573 34051 31631 34057
rect 31573 34017 31585 34051
rect 31619 34048 31631 34051
rect 31754 34048 31760 34060
rect 31619 34020 31760 34048
rect 31619 34017 31631 34020
rect 31573 34011 31631 34017
rect 31754 34008 31760 34020
rect 31812 34008 31818 34060
rect 32416 34057 32444 34088
rect 32585 34085 32597 34119
rect 32631 34116 32643 34119
rect 33410 34116 33416 34128
rect 32631 34088 33416 34116
rect 32631 34085 32643 34088
rect 32585 34079 32643 34085
rect 33410 34076 33416 34088
rect 33468 34076 33474 34128
rect 32401 34051 32459 34057
rect 32401 34017 32413 34051
rect 32447 34017 32459 34051
rect 33505 34051 33563 34057
rect 33505 34048 33517 34051
rect 32401 34011 32459 34017
rect 32692 34020 33517 34048
rect 32692 33992 32720 34020
rect 33505 34017 33517 34020
rect 33551 34017 33563 34051
rect 33704 34048 33732 34156
rect 33781 34153 33793 34187
rect 33827 34184 33839 34187
rect 35526 34184 35532 34196
rect 33827 34156 35532 34184
rect 33827 34153 33839 34156
rect 33781 34147 33839 34153
rect 35526 34144 35532 34156
rect 35584 34144 35590 34196
rect 35544 34116 35572 34144
rect 38933 34119 38991 34125
rect 35544 34088 36308 34116
rect 34974 34048 34980 34060
rect 33704 34020 34980 34048
rect 33505 34011 33563 34017
rect 34974 34008 34980 34020
rect 35032 34008 35038 34060
rect 35437 34051 35495 34057
rect 35437 34017 35449 34051
rect 35483 34017 35495 34051
rect 35437 34011 35495 34017
rect 31297 33983 31355 33989
rect 31297 33949 31309 33983
rect 31343 33980 31355 33983
rect 31343 33952 31432 33980
rect 31343 33949 31355 33952
rect 31297 33943 31355 33949
rect 31404 33924 31432 33952
rect 31478 33940 31484 33992
rect 31536 33980 31542 33992
rect 32674 33980 32680 33992
rect 31536 33952 31581 33980
rect 32635 33952 32680 33980
rect 31536 33940 31542 33952
rect 32674 33940 32680 33952
rect 32732 33940 32738 33992
rect 33134 33980 33140 33992
rect 33095 33952 33140 33980
rect 33134 33940 33140 33952
rect 33192 33940 33198 33992
rect 33321 33983 33379 33989
rect 33321 33949 33333 33983
rect 33367 33949 33379 33983
rect 33321 33943 33379 33949
rect 33597 33983 33655 33989
rect 33597 33949 33609 33983
rect 33643 33949 33655 33983
rect 33597 33943 33655 33949
rect 31386 33872 31392 33924
rect 31444 33872 31450 33924
rect 32401 33915 32459 33921
rect 32401 33881 32413 33915
rect 32447 33912 32459 33915
rect 33336 33912 33364 33943
rect 32447 33884 33364 33912
rect 32447 33881 32459 33884
rect 32401 33875 32459 33881
rect 31294 33844 31300 33856
rect 31220 33816 31300 33844
rect 31113 33807 31171 33813
rect 31294 33804 31300 33816
rect 31352 33844 31358 33856
rect 31846 33844 31852 33856
rect 31352 33816 31852 33844
rect 31352 33804 31358 33816
rect 31846 33804 31852 33816
rect 31904 33804 31910 33856
rect 32766 33804 32772 33856
rect 32824 33844 32830 33856
rect 33612 33844 33640 33943
rect 34422 33940 34428 33992
rect 34480 33980 34486 33992
rect 35069 33983 35127 33989
rect 35069 33980 35081 33983
rect 34480 33952 35081 33980
rect 34480 33940 34486 33952
rect 35069 33949 35081 33952
rect 35115 33949 35127 33983
rect 35452 33980 35480 34011
rect 35710 33980 35716 33992
rect 35452 33952 35716 33980
rect 35069 33943 35127 33949
rect 35710 33940 35716 33952
rect 35768 33980 35774 33992
rect 36280 33989 36308 34088
rect 38933 34085 38945 34119
rect 38979 34116 38991 34119
rect 40218 34116 40224 34128
rect 38979 34088 40224 34116
rect 38979 34085 38991 34088
rect 38933 34079 38991 34085
rect 40218 34076 40224 34088
rect 40276 34076 40282 34128
rect 36081 33983 36139 33989
rect 36081 33980 36093 33983
rect 35768 33952 36093 33980
rect 35768 33940 35774 33952
rect 36081 33949 36093 33952
rect 36127 33949 36139 33983
rect 36081 33943 36139 33949
rect 36265 33983 36323 33989
rect 36265 33949 36277 33983
rect 36311 33980 36323 33983
rect 36630 33980 36636 33992
rect 36311 33952 36636 33980
rect 36311 33949 36323 33952
rect 36265 33943 36323 33949
rect 36630 33940 36636 33952
rect 36688 33940 36694 33992
rect 38657 33983 38715 33989
rect 38657 33949 38669 33983
rect 38703 33949 38715 33983
rect 38930 33980 38936 33992
rect 38891 33952 38936 33980
rect 38657 33943 38715 33949
rect 38672 33912 38700 33943
rect 38930 33940 38936 33952
rect 38988 33940 38994 33992
rect 38838 33912 38844 33924
rect 38672 33884 38844 33912
rect 38838 33872 38844 33884
rect 38896 33872 38902 33924
rect 34241 33847 34299 33853
rect 34241 33844 34253 33847
rect 32824 33816 34253 33844
rect 32824 33804 32830 33816
rect 34241 33813 34253 33816
rect 34287 33813 34299 33847
rect 34241 33807 34299 33813
rect 35802 33804 35808 33856
rect 35860 33844 35866 33856
rect 35897 33847 35955 33853
rect 35897 33844 35909 33847
rect 35860 33816 35909 33844
rect 35860 33804 35866 33816
rect 35897 33813 35909 33816
rect 35943 33813 35955 33847
rect 38746 33844 38752 33856
rect 38707 33816 38752 33844
rect 35897 33807 35955 33813
rect 38746 33804 38752 33816
rect 38804 33804 38810 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 19521 33643 19579 33649
rect 19521 33640 19533 33643
rect 19484 33612 19533 33640
rect 19484 33600 19490 33612
rect 19521 33609 19533 33612
rect 19567 33609 19579 33643
rect 19521 33603 19579 33609
rect 19705 33643 19763 33649
rect 19705 33609 19717 33643
rect 19751 33640 19763 33643
rect 21082 33640 21088 33652
rect 19751 33612 21088 33640
rect 19751 33609 19763 33612
rect 19705 33603 19763 33609
rect 19720 33572 19748 33603
rect 21082 33600 21088 33612
rect 21140 33600 21146 33652
rect 22186 33640 22192 33652
rect 22147 33612 22192 33640
rect 22186 33600 22192 33612
rect 22244 33600 22250 33652
rect 23014 33640 23020 33652
rect 22975 33612 23020 33640
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 25133 33643 25191 33649
rect 23308 33612 25008 33640
rect 17788 33544 19748 33572
rect 15013 33507 15071 33513
rect 15013 33473 15025 33507
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33473 15899 33507
rect 15841 33467 15899 33473
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 16206 33504 16212 33516
rect 16071 33476 16212 33504
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 15028 33368 15056 33467
rect 15105 33439 15163 33445
rect 15105 33405 15117 33439
rect 15151 33436 15163 33439
rect 15194 33436 15200 33448
rect 15151 33408 15200 33436
rect 15151 33405 15163 33408
rect 15105 33399 15163 33405
rect 15194 33396 15200 33408
rect 15252 33396 15258 33448
rect 15286 33396 15292 33448
rect 15344 33436 15350 33448
rect 15381 33439 15439 33445
rect 15381 33436 15393 33439
rect 15344 33408 15393 33436
rect 15344 33396 15350 33408
rect 15381 33405 15393 33408
rect 15427 33436 15439 33439
rect 15856 33436 15884 33467
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 15427 33408 15884 33436
rect 17788 33436 17816 33544
rect 23198 33532 23204 33584
rect 23256 33572 23262 33584
rect 23308 33572 23336 33612
rect 24026 33572 24032 33584
rect 23256 33544 23336 33572
rect 23939 33544 24032 33572
rect 23256 33532 23262 33544
rect 17954 33504 17960 33516
rect 17915 33476 17960 33504
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 18506 33464 18512 33516
rect 18564 33504 18570 33516
rect 19337 33507 19395 33513
rect 19337 33504 19349 33507
rect 18564 33476 19349 33504
rect 18564 33464 18570 33476
rect 19337 33473 19349 33476
rect 19383 33473 19395 33507
rect 19337 33467 19395 33473
rect 19613 33507 19671 33513
rect 19613 33473 19625 33507
rect 19659 33504 19671 33507
rect 20254 33504 20260 33516
rect 19659 33476 20260 33504
rect 19659 33473 19671 33476
rect 19613 33467 19671 33473
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 20714 33464 20720 33516
rect 20772 33504 20778 33516
rect 20809 33507 20867 33513
rect 20809 33504 20821 33507
rect 20772 33476 20821 33504
rect 20772 33464 20778 33476
rect 20809 33473 20821 33476
rect 20855 33473 20867 33507
rect 20990 33504 20996 33516
rect 20951 33476 20996 33504
rect 20809 33467 20867 33473
rect 20990 33464 20996 33476
rect 21048 33464 21054 33516
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22833 33507 22891 33513
rect 22833 33504 22845 33507
rect 22428 33476 22845 33504
rect 22428 33464 22434 33476
rect 22833 33473 22845 33476
rect 22879 33504 22891 33507
rect 23106 33504 23112 33516
rect 22879 33476 23112 33504
rect 22879 33473 22891 33476
rect 22833 33467 22891 33473
rect 23106 33464 23112 33476
rect 23164 33464 23170 33516
rect 23308 33513 23336 33544
rect 24026 33532 24032 33544
rect 24084 33572 24090 33584
rect 24578 33572 24584 33584
rect 24084 33544 24584 33572
rect 24084 33532 24090 33544
rect 24578 33532 24584 33544
rect 24636 33532 24642 33584
rect 24762 33572 24768 33584
rect 24723 33544 24768 33572
rect 24762 33532 24768 33544
rect 24820 33532 24826 33584
rect 24980 33572 25008 33612
rect 25133 33609 25145 33643
rect 25179 33640 25191 33643
rect 25590 33640 25596 33652
rect 25179 33612 25596 33640
rect 25179 33609 25191 33612
rect 25133 33603 25191 33609
rect 25590 33600 25596 33612
rect 25648 33600 25654 33652
rect 26602 33600 26608 33652
rect 26660 33600 26666 33652
rect 27246 33640 27252 33652
rect 27207 33612 27252 33640
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 28166 33640 28172 33652
rect 28127 33612 28172 33640
rect 28166 33600 28172 33612
rect 28224 33600 28230 33652
rect 28718 33600 28724 33652
rect 28776 33640 28782 33652
rect 30377 33643 30435 33649
rect 30377 33640 30389 33643
rect 28776 33612 30389 33640
rect 28776 33600 28782 33612
rect 30377 33609 30389 33612
rect 30423 33640 30435 33643
rect 31754 33640 31760 33652
rect 30423 33612 31760 33640
rect 30423 33609 30435 33612
rect 30377 33603 30435 33609
rect 31754 33600 31760 33612
rect 31812 33600 31818 33652
rect 33870 33600 33876 33652
rect 33928 33640 33934 33652
rect 34793 33643 34851 33649
rect 34793 33640 34805 33643
rect 33928 33612 34805 33640
rect 33928 33600 33934 33612
rect 34793 33609 34805 33612
rect 34839 33609 34851 33643
rect 34793 33603 34851 33609
rect 34974 33600 34980 33652
rect 35032 33640 35038 33652
rect 36265 33643 36323 33649
rect 36265 33640 36277 33643
rect 35032 33612 36277 33640
rect 35032 33600 35038 33612
rect 36265 33609 36277 33612
rect 36311 33640 36323 33643
rect 37458 33640 37464 33652
rect 36311 33612 37464 33640
rect 36311 33609 36323 33612
rect 36265 33603 36323 33609
rect 37458 33600 37464 33612
rect 37516 33600 37522 33652
rect 37829 33643 37887 33649
rect 37829 33609 37841 33643
rect 37875 33640 37887 33643
rect 38381 33643 38439 33649
rect 38381 33640 38393 33643
rect 37875 33612 38393 33640
rect 37875 33609 37887 33612
rect 37829 33603 37887 33609
rect 38381 33609 38393 33612
rect 38427 33640 38439 33643
rect 38746 33640 38752 33652
rect 38427 33612 38752 33640
rect 38427 33609 38439 33612
rect 38381 33603 38439 33609
rect 38746 33600 38752 33612
rect 38804 33600 38810 33652
rect 25038 33572 25044 33584
rect 24980 33541 25044 33572
rect 23293 33507 23351 33513
rect 23293 33473 23305 33507
rect 23339 33473 23351 33507
rect 23293 33467 23351 33473
rect 23566 33464 23572 33516
rect 23624 33504 23630 33516
rect 23753 33507 23811 33513
rect 23753 33504 23765 33507
rect 23624 33476 23765 33504
rect 23624 33464 23630 33476
rect 23753 33473 23765 33476
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 24980 33510 25007 33541
rect 24995 33507 25007 33510
rect 25041 33532 25044 33541
rect 25096 33532 25102 33584
rect 26418 33572 26424 33584
rect 26379 33544 26424 33572
rect 26418 33532 26424 33544
rect 26476 33532 26482 33584
rect 26620 33572 26648 33600
rect 27433 33575 27491 33581
rect 26620 33544 27292 33572
rect 25041 33507 25053 33532
rect 23900 33476 23945 33504
rect 24995 33501 25053 33507
rect 25590 33504 25596 33516
rect 25551 33476 25596 33504
rect 23900 33464 23906 33476
rect 25590 33464 25596 33476
rect 25648 33464 25654 33516
rect 25777 33507 25835 33513
rect 25777 33473 25789 33507
rect 25823 33473 25835 33507
rect 25777 33467 25835 33473
rect 26605 33507 26663 33513
rect 26605 33473 26617 33507
rect 26651 33473 26663 33507
rect 27154 33504 27160 33516
rect 27115 33476 27160 33504
rect 26605 33467 26663 33473
rect 17865 33439 17923 33445
rect 17865 33436 17877 33439
rect 17788 33408 17877 33436
rect 15427 33405 15439 33408
rect 15381 33399 15439 33405
rect 17865 33405 17877 33408
rect 17911 33405 17923 33439
rect 20625 33439 20683 33445
rect 20625 33436 20637 33439
rect 17865 33399 17923 33405
rect 17972 33408 20637 33436
rect 15654 33368 15660 33380
rect 15028 33340 15660 33368
rect 15654 33328 15660 33340
rect 15712 33368 15718 33380
rect 17972 33368 18000 33408
rect 20625 33405 20637 33408
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 20901 33439 20959 33445
rect 20901 33405 20913 33439
rect 20947 33405 20959 33439
rect 20901 33399 20959 33405
rect 21085 33439 21143 33445
rect 21085 33405 21097 33439
rect 21131 33436 21143 33439
rect 22649 33439 22707 33445
rect 22649 33436 22661 33439
rect 21131 33408 22661 33436
rect 21131 33405 21143 33408
rect 21085 33399 21143 33405
rect 22649 33405 22661 33408
rect 22695 33405 22707 33439
rect 22649 33399 22707 33405
rect 15712 33340 18000 33368
rect 20916 33368 20944 33399
rect 22922 33396 22928 33448
rect 22980 33436 22986 33448
rect 23201 33439 23259 33445
rect 22980 33408 23025 33436
rect 22980 33396 22986 33408
rect 23201 33405 23213 33439
rect 23247 33436 23259 33439
rect 23658 33436 23664 33448
rect 23247 33408 23664 33436
rect 23247 33405 23259 33408
rect 23201 33399 23259 33405
rect 23658 33396 23664 33408
rect 23716 33436 23722 33448
rect 24946 33436 24952 33448
rect 23716 33408 24952 33436
rect 23716 33396 23722 33408
rect 24946 33396 24952 33408
rect 25004 33396 25010 33448
rect 25792 33436 25820 33467
rect 26620 33436 26648 33467
rect 27154 33464 27160 33476
rect 27212 33464 27218 33516
rect 27264 33504 27292 33544
rect 27433 33541 27445 33575
rect 27479 33572 27491 33575
rect 30466 33572 30472 33584
rect 27479 33544 30472 33572
rect 27479 33541 27491 33544
rect 27433 33535 27491 33541
rect 30466 33532 30472 33544
rect 30524 33532 30530 33584
rect 31294 33572 31300 33584
rect 31036 33544 31300 33572
rect 30282 33504 30288 33516
rect 27264 33476 30288 33504
rect 30282 33464 30288 33476
rect 30340 33464 30346 33516
rect 31036 33513 31064 33544
rect 31294 33532 31300 33544
rect 31352 33532 31358 33584
rect 33134 33572 33140 33584
rect 32324 33544 33140 33572
rect 31021 33507 31079 33513
rect 31021 33473 31033 33507
rect 31067 33473 31079 33507
rect 31202 33504 31208 33516
rect 31163 33476 31208 33504
rect 31021 33467 31079 33473
rect 31202 33464 31208 33476
rect 31260 33464 31266 33516
rect 31386 33464 31392 33516
rect 31444 33504 31450 33516
rect 32324 33513 32352 33544
rect 33134 33532 33140 33544
rect 33192 33532 33198 33584
rect 33594 33572 33600 33584
rect 33555 33544 33600 33572
rect 33594 33532 33600 33544
rect 33652 33532 33658 33584
rect 33781 33575 33839 33581
rect 33781 33541 33793 33575
rect 33827 33572 33839 33575
rect 34146 33572 34152 33584
rect 33827 33544 34152 33572
rect 33827 33541 33839 33544
rect 33781 33535 33839 33541
rect 34146 33532 34152 33544
rect 34204 33532 34210 33584
rect 38838 33572 38844 33584
rect 35636 33544 38844 33572
rect 35636 33516 35664 33544
rect 31665 33507 31723 33513
rect 31665 33504 31677 33507
rect 31444 33476 31677 33504
rect 31444 33464 31450 33476
rect 31665 33473 31677 33476
rect 31711 33473 31723 33507
rect 31665 33467 31723 33473
rect 32309 33507 32367 33513
rect 32309 33473 32321 33507
rect 32355 33473 32367 33507
rect 32490 33504 32496 33516
rect 32451 33476 32496 33504
rect 32309 33467 32367 33473
rect 32490 33464 32496 33476
rect 32548 33464 32554 33516
rect 32585 33507 32643 33513
rect 32585 33473 32597 33507
rect 32631 33473 32643 33507
rect 32585 33467 32643 33473
rect 32677 33507 32735 33513
rect 32677 33473 32689 33507
rect 32723 33504 32735 33507
rect 32766 33504 32772 33516
rect 32723 33476 32772 33504
rect 32723 33473 32735 33476
rect 32677 33467 32735 33473
rect 25792 33408 27476 33436
rect 21634 33368 21640 33380
rect 20916 33340 21640 33368
rect 15712 33328 15718 33340
rect 21634 33328 21640 33340
rect 21692 33328 21698 33380
rect 15930 33260 15936 33312
rect 15988 33300 15994 33312
rect 16025 33303 16083 33309
rect 16025 33300 16037 33303
rect 15988 33272 16037 33300
rect 15988 33260 15994 33272
rect 16025 33269 16037 33272
rect 16071 33269 16083 33303
rect 16025 33263 16083 33269
rect 17589 33303 17647 33309
rect 17589 33269 17601 33303
rect 17635 33300 17647 33303
rect 18414 33300 18420 33312
rect 17635 33272 18420 33300
rect 17635 33269 17647 33272
rect 17589 33263 17647 33269
rect 18414 33260 18420 33272
rect 18472 33260 18478 33312
rect 19889 33303 19947 33309
rect 19889 33269 19901 33303
rect 19935 33300 19947 33303
rect 20438 33300 20444 33312
rect 19935 33272 20444 33300
rect 19935 33269 19947 33272
rect 19889 33263 19947 33269
rect 20438 33260 20444 33272
rect 20496 33260 20502 33312
rect 23566 33260 23572 33312
rect 23624 33300 23630 33312
rect 24980 33309 25008 33396
rect 25685 33371 25743 33377
rect 25685 33337 25697 33371
rect 25731 33368 25743 33371
rect 26694 33368 26700 33380
rect 25731 33340 26700 33368
rect 25731 33337 25743 33340
rect 25685 33331 25743 33337
rect 26694 33328 26700 33340
rect 26752 33328 26758 33380
rect 27448 33377 27476 33408
rect 32214 33396 32220 33448
rect 32272 33436 32278 33448
rect 32600 33436 32628 33467
rect 32766 33464 32772 33476
rect 32824 33504 32830 33516
rect 34241 33507 34299 33513
rect 34241 33504 34253 33507
rect 32824 33476 34253 33504
rect 32824 33464 32830 33476
rect 34241 33473 34253 33476
rect 34287 33473 34299 33507
rect 35618 33504 35624 33516
rect 35579 33476 35624 33504
rect 34241 33467 34299 33473
rect 35618 33464 35624 33476
rect 35676 33464 35682 33516
rect 35802 33504 35808 33516
rect 35763 33476 35808 33504
rect 35802 33464 35808 33476
rect 35860 33464 35866 33516
rect 36630 33504 36636 33516
rect 36591 33476 36636 33504
rect 36630 33464 36636 33476
rect 36688 33464 36694 33516
rect 37458 33504 37464 33516
rect 37419 33476 37464 33504
rect 37458 33464 37464 33476
rect 37516 33464 37522 33516
rect 38304 33513 38332 33544
rect 38838 33532 38844 33544
rect 38896 33532 38902 33584
rect 37645 33507 37703 33513
rect 37645 33473 37657 33507
rect 37691 33473 37703 33507
rect 37645 33467 37703 33473
rect 38289 33507 38347 33513
rect 38289 33473 38301 33507
rect 38335 33473 38347 33507
rect 38289 33467 38347 33473
rect 38565 33507 38623 33513
rect 38565 33473 38577 33507
rect 38611 33504 38623 33507
rect 38930 33504 38936 33516
rect 38611 33476 38936 33504
rect 38611 33473 38623 33476
rect 38565 33467 38623 33473
rect 33413 33439 33471 33445
rect 33413 33436 33425 33439
rect 32272 33408 33425 33436
rect 32272 33396 32278 33408
rect 33413 33405 33425 33408
rect 33459 33405 33471 33439
rect 35526 33436 35532 33448
rect 33413 33399 33471 33405
rect 33612 33408 35532 33436
rect 27433 33371 27491 33377
rect 27433 33337 27445 33371
rect 27479 33337 27491 33371
rect 29178 33368 29184 33380
rect 29091 33340 29184 33368
rect 27433 33331 27491 33337
rect 29178 33328 29184 33340
rect 29236 33368 29242 33380
rect 33612 33368 33640 33408
rect 35526 33396 35532 33408
rect 35584 33396 35590 33448
rect 36722 33436 36728 33448
rect 36683 33408 36728 33436
rect 36722 33396 36728 33408
rect 36780 33396 36786 33448
rect 29236 33340 33640 33368
rect 29236 33328 29242 33340
rect 34422 33328 34428 33380
rect 34480 33368 34486 33380
rect 37660 33368 37688 33467
rect 38930 33464 38936 33476
rect 38988 33464 38994 33516
rect 39666 33504 39672 33516
rect 39627 33476 39672 33504
rect 39666 33464 39672 33476
rect 39724 33464 39730 33516
rect 40034 33504 40040 33516
rect 39995 33476 40040 33504
rect 40034 33464 40040 33476
rect 40092 33464 40098 33516
rect 40681 33439 40739 33445
rect 40681 33405 40693 33439
rect 40727 33436 40739 33439
rect 52270 33436 52276 33448
rect 40727 33408 52276 33436
rect 40727 33405 40739 33408
rect 40681 33399 40739 33405
rect 52270 33396 52276 33408
rect 52328 33396 52334 33448
rect 34480 33340 37688 33368
rect 34480 33328 34486 33340
rect 24029 33303 24087 33309
rect 24029 33300 24041 33303
rect 23624 33272 24041 33300
rect 23624 33260 23630 33272
rect 24029 33269 24041 33272
rect 24075 33269 24087 33303
rect 24029 33263 24087 33269
rect 24971 33303 25029 33309
rect 24971 33269 24983 33303
rect 25017 33269 25029 33303
rect 24971 33263 25029 33269
rect 26237 33303 26295 33309
rect 26237 33269 26249 33303
rect 26283 33300 26295 33303
rect 26326 33300 26332 33312
rect 26283 33272 26332 33300
rect 26283 33269 26295 33272
rect 26237 33263 26295 33269
rect 26326 33260 26332 33272
rect 26384 33260 26390 33312
rect 30834 33260 30840 33312
rect 30892 33300 30898 33312
rect 31205 33303 31263 33309
rect 31205 33300 31217 33303
rect 30892 33272 31217 33300
rect 30892 33260 30898 33272
rect 31205 33269 31217 33272
rect 31251 33269 31263 33303
rect 32950 33300 32956 33312
rect 32911 33272 32956 33300
rect 31205 33263 31263 33269
rect 32950 33260 32956 33272
rect 33008 33260 33014 33312
rect 35710 33300 35716 33312
rect 35671 33272 35716 33300
rect 35710 33260 35716 33272
rect 35768 33260 35774 33312
rect 36814 33260 36820 33312
rect 36872 33300 36878 33312
rect 36909 33303 36967 33309
rect 36909 33300 36921 33303
rect 36872 33272 36921 33300
rect 36872 33260 36878 33272
rect 36909 33269 36921 33272
rect 36955 33269 36967 33303
rect 38746 33300 38752 33312
rect 38707 33272 38752 33300
rect 36909 33263 36967 33269
rect 38746 33260 38752 33272
rect 38804 33260 38810 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 21266 33056 21272 33108
rect 21324 33096 21330 33108
rect 22097 33099 22155 33105
rect 22097 33096 22109 33099
rect 21324 33068 22109 33096
rect 21324 33056 21330 33068
rect 22097 33065 22109 33068
rect 22143 33065 22155 33099
rect 22097 33059 22155 33065
rect 22830 33056 22836 33108
rect 22888 33096 22894 33108
rect 26602 33096 26608 33108
rect 22888 33068 26608 33096
rect 22888 33056 22894 33068
rect 26602 33056 26608 33068
rect 26660 33056 26666 33108
rect 26786 33056 26792 33108
rect 26844 33096 26850 33108
rect 31294 33096 31300 33108
rect 26844 33068 31300 33096
rect 26844 33056 26850 33068
rect 31294 33056 31300 33068
rect 31352 33056 31358 33108
rect 31938 33096 31944 33108
rect 31899 33068 31944 33096
rect 31938 33056 31944 33068
rect 31996 33056 32002 33108
rect 32309 33099 32367 33105
rect 32309 33065 32321 33099
rect 32355 33096 32367 33099
rect 32490 33096 32496 33108
rect 32355 33068 32496 33096
rect 32355 33065 32367 33068
rect 32309 33059 32367 33065
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 33226 33096 33232 33108
rect 33187 33068 33232 33096
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 34054 33096 34060 33108
rect 34015 33068 34060 33096
rect 34054 33056 34060 33068
rect 34112 33056 34118 33108
rect 38838 33096 38844 33108
rect 38799 33068 38844 33096
rect 38838 33056 38844 33068
rect 38896 33056 38902 33108
rect 40034 33056 40040 33108
rect 40092 33096 40098 33108
rect 40405 33099 40463 33105
rect 40405 33096 40417 33099
rect 40092 33068 40417 33096
rect 40092 33056 40098 33068
rect 40405 33065 40417 33068
rect 40451 33065 40463 33099
rect 40405 33059 40463 33065
rect 15194 32988 15200 33040
rect 15252 33028 15258 33040
rect 15933 33031 15991 33037
rect 15933 33028 15945 33031
rect 15252 33000 15945 33028
rect 15252 32988 15258 33000
rect 15933 32997 15945 33000
rect 15979 33028 15991 33031
rect 16761 33031 16819 33037
rect 16761 33028 16773 33031
rect 15979 33000 16773 33028
rect 15979 32997 15991 33000
rect 15933 32991 15991 32997
rect 16761 32997 16773 33000
rect 16807 32997 16819 33031
rect 16761 32991 16819 32997
rect 20438 32988 20444 33040
rect 20496 33028 20502 33040
rect 20496 33000 23244 33028
rect 20496 32988 20502 33000
rect 15654 32960 15660 32972
rect 15615 32932 15660 32960
rect 15654 32920 15660 32932
rect 15712 32920 15718 32972
rect 17221 32963 17279 32969
rect 17221 32929 17233 32963
rect 17267 32960 17279 32963
rect 18322 32960 18328 32972
rect 17267 32932 18328 32960
rect 17267 32929 17279 32932
rect 17221 32923 17279 32929
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 20993 32963 21051 32969
rect 20993 32929 21005 32963
rect 21039 32960 21051 32963
rect 22094 32960 22100 32972
rect 21039 32932 21956 32960
rect 21039 32929 21051 32932
rect 20993 32923 21051 32929
rect 17129 32895 17187 32901
rect 17129 32861 17141 32895
rect 17175 32892 17187 32895
rect 17402 32892 17408 32904
rect 17175 32864 17408 32892
rect 17175 32861 17187 32864
rect 17129 32855 17187 32861
rect 17402 32852 17408 32864
rect 17460 32852 17466 32904
rect 17770 32852 17776 32904
rect 17828 32892 17834 32904
rect 20809 32895 20867 32901
rect 20809 32892 20821 32895
rect 17828 32864 20821 32892
rect 17828 32852 17834 32864
rect 20809 32861 20821 32864
rect 20855 32861 20867 32895
rect 21266 32892 21272 32904
rect 21227 32864 21272 32892
rect 20809 32855 20867 32861
rect 18877 32827 18935 32833
rect 18877 32793 18889 32827
rect 18923 32824 18935 32827
rect 19242 32824 19248 32836
rect 18923 32796 19248 32824
rect 18923 32793 18935 32796
rect 18877 32787 18935 32793
rect 19242 32784 19248 32796
rect 19300 32824 19306 32836
rect 19521 32827 19579 32833
rect 19521 32824 19533 32827
rect 19300 32796 19533 32824
rect 19300 32784 19306 32796
rect 19521 32793 19533 32796
rect 19567 32793 19579 32827
rect 19521 32787 19579 32793
rect 16114 32756 16120 32768
rect 16075 32728 16120 32756
rect 16114 32716 16120 32728
rect 16172 32716 16178 32768
rect 18598 32716 18604 32768
rect 18656 32756 18662 32768
rect 19797 32759 19855 32765
rect 19797 32756 19809 32759
rect 18656 32728 19809 32756
rect 18656 32716 18662 32728
rect 19797 32725 19809 32728
rect 19843 32756 19855 32759
rect 20622 32756 20628 32768
rect 19843 32728 20628 32756
rect 19843 32725 19855 32728
rect 19797 32719 19855 32725
rect 20622 32716 20628 32728
rect 20680 32716 20686 32768
rect 20824 32756 20852 32855
rect 21266 32852 21272 32864
rect 21324 32852 21330 32904
rect 21928 32901 21956 32932
rect 22066 32920 22100 32960
rect 22152 32960 22158 32972
rect 22189 32963 22247 32969
rect 22189 32960 22201 32963
rect 22152 32932 22201 32960
rect 22152 32920 22158 32932
rect 22189 32929 22201 32932
rect 22235 32929 22247 32963
rect 22189 32923 22247 32929
rect 21913 32895 21971 32901
rect 21913 32861 21925 32895
rect 21959 32861 21971 32895
rect 21913 32855 21971 32861
rect 21177 32827 21235 32833
rect 21177 32793 21189 32827
rect 21223 32824 21235 32827
rect 22066 32824 22094 32920
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 23017 32895 23075 32901
rect 23017 32892 23029 32895
rect 22888 32864 23029 32892
rect 22888 32852 22894 32864
rect 23017 32861 23029 32864
rect 23063 32861 23075 32895
rect 23017 32855 23075 32861
rect 23216 32833 23244 33000
rect 23382 32988 23388 33040
rect 23440 33028 23446 33040
rect 26050 33028 26056 33040
rect 23440 33000 26056 33028
rect 23440 32988 23446 33000
rect 26050 32988 26056 33000
rect 26108 32988 26114 33040
rect 26510 32988 26516 33040
rect 26568 33028 26574 33040
rect 27801 33031 27859 33037
rect 26568 33000 27384 33028
rect 26568 32988 26574 33000
rect 25682 32960 25688 32972
rect 23308 32932 25688 32960
rect 23308 32904 23336 32932
rect 25682 32920 25688 32932
rect 25740 32920 25746 32972
rect 25866 32920 25872 32972
rect 25924 32960 25930 32972
rect 26236 32963 26294 32969
rect 26236 32960 26248 32963
rect 25924 32932 26248 32960
rect 25924 32920 25930 32932
rect 26236 32929 26248 32932
rect 26282 32929 26294 32963
rect 26236 32923 26294 32929
rect 26429 32963 26487 32969
rect 26429 32929 26441 32963
rect 26475 32960 26487 32963
rect 26694 32960 26700 32972
rect 26475 32932 26700 32960
rect 26475 32929 26487 32932
rect 26429 32923 26487 32929
rect 26694 32920 26700 32932
rect 26752 32920 26758 32972
rect 27356 32969 27384 33000
rect 27801 32997 27813 33031
rect 27847 32997 27859 33031
rect 27801 32991 27859 32997
rect 29825 33031 29883 33037
rect 29825 32997 29837 33031
rect 29871 33028 29883 33031
rect 34422 33028 34428 33040
rect 29871 33000 34428 33028
rect 29871 32997 29883 33000
rect 29825 32991 29883 32997
rect 27341 32963 27399 32969
rect 27341 32929 27353 32963
rect 27387 32929 27399 32963
rect 27341 32923 27399 32929
rect 23290 32852 23296 32904
rect 23348 32892 23354 32904
rect 24581 32895 24639 32901
rect 23348 32864 23441 32892
rect 23348 32852 23354 32864
rect 24581 32861 24593 32895
rect 24627 32892 24639 32895
rect 24670 32892 24676 32904
rect 24627 32864 24676 32892
rect 24627 32861 24639 32864
rect 24581 32855 24639 32861
rect 24670 32852 24676 32864
rect 24728 32852 24734 32904
rect 24854 32852 24860 32904
rect 24912 32892 24918 32904
rect 26145 32895 26203 32901
rect 26145 32892 26157 32895
rect 24912 32864 26157 32892
rect 24912 32852 24918 32864
rect 26145 32861 26157 32864
rect 26191 32861 26203 32895
rect 26145 32855 26203 32861
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26384 32864 26428 32892
rect 26384 32852 26390 32864
rect 27154 32852 27160 32904
rect 27212 32892 27218 32904
rect 27433 32895 27491 32901
rect 27433 32892 27445 32895
rect 27212 32864 27445 32892
rect 27212 32852 27218 32864
rect 27433 32861 27445 32864
rect 27479 32861 27491 32895
rect 27816 32892 27844 32991
rect 34422 32988 34428 33000
rect 34480 32988 34486 33040
rect 36630 33028 36636 33040
rect 36556 33000 36636 33028
rect 28258 32920 28264 32972
rect 28316 32960 28322 32972
rect 28537 32963 28595 32969
rect 28537 32960 28549 32963
rect 28316 32932 28549 32960
rect 28316 32920 28322 32932
rect 28537 32929 28549 32932
rect 28583 32929 28595 32963
rect 28537 32923 28595 32929
rect 28997 32963 29055 32969
rect 28997 32929 29009 32963
rect 29043 32929 29055 32963
rect 28997 32923 29055 32929
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 27816 32864 28641 32892
rect 27433 32855 27491 32861
rect 28629 32861 28641 32864
rect 28675 32892 28687 32895
rect 28810 32892 28816 32904
rect 28675 32864 28816 32892
rect 28675 32861 28687 32864
rect 28629 32855 28687 32861
rect 28810 32852 28816 32864
rect 28868 32852 28874 32904
rect 29012 32892 29040 32923
rect 29086 32920 29092 32972
rect 29144 32960 29150 32972
rect 32214 32960 32220 32972
rect 29144 32932 29960 32960
rect 32175 32932 32220 32960
rect 29144 32920 29150 32932
rect 29932 32901 29960 32932
rect 32214 32920 32220 32932
rect 32272 32920 32278 32972
rect 32766 32920 32772 32972
rect 32824 32960 32830 32972
rect 36556 32969 36584 33000
rect 36630 32988 36636 33000
rect 36688 32988 36694 33040
rect 36541 32963 36599 32969
rect 32824 32932 33364 32960
rect 32824 32920 32830 32932
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 29012 32864 29745 32892
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29917 32895 29975 32901
rect 29917 32861 29929 32895
rect 29963 32861 29975 32895
rect 29917 32855 29975 32861
rect 31754 32852 31760 32904
rect 31812 32892 31818 32904
rect 31849 32895 31907 32901
rect 31849 32892 31861 32895
rect 31812 32864 31861 32892
rect 31812 32852 31818 32864
rect 31849 32861 31861 32864
rect 31895 32861 31907 32895
rect 32122 32892 32128 32904
rect 32083 32864 32128 32892
rect 31849 32855 31907 32861
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 32674 32852 32680 32904
rect 32732 32892 32738 32904
rect 33336 32901 33364 32932
rect 36541 32929 36553 32963
rect 36587 32929 36599 32963
rect 36541 32923 36599 32929
rect 37001 32963 37059 32969
rect 37001 32929 37013 32963
rect 37047 32960 37059 32963
rect 37274 32960 37280 32972
rect 37047 32932 37280 32960
rect 37047 32929 37059 32932
rect 37001 32923 37059 32929
rect 37274 32920 37280 32932
rect 37332 32960 37338 32972
rect 37332 32932 37688 32960
rect 37332 32920 37338 32932
rect 33229 32895 33287 32901
rect 33229 32892 33241 32895
rect 32732 32864 33241 32892
rect 32732 32852 32738 32864
rect 33229 32861 33241 32864
rect 33275 32861 33287 32895
rect 33229 32855 33287 32861
rect 33321 32895 33379 32901
rect 33321 32861 33333 32895
rect 33367 32892 33379 32895
rect 34885 32895 34943 32901
rect 34885 32892 34897 32895
rect 33367 32864 34897 32892
rect 33367 32861 33379 32864
rect 33321 32855 33379 32861
rect 34885 32861 34897 32864
rect 34931 32861 34943 32895
rect 35802 32892 35808 32904
rect 35763 32864 35808 32892
rect 34885 32855 34943 32861
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 35986 32892 35992 32904
rect 35947 32864 35992 32892
rect 35986 32852 35992 32864
rect 36044 32852 36050 32904
rect 36633 32895 36691 32901
rect 36633 32861 36645 32895
rect 36679 32861 36691 32895
rect 36814 32892 36820 32904
rect 36775 32864 36820 32892
rect 36633 32855 36691 32861
rect 21223 32796 22094 32824
rect 23201 32827 23259 32833
rect 21223 32793 21235 32796
rect 21177 32787 21235 32793
rect 23201 32793 23213 32827
rect 23247 32824 23259 32827
rect 25041 32827 25099 32833
rect 23247 32796 24808 32824
rect 23247 32793 23259 32796
rect 23201 32787 23259 32793
rect 21358 32756 21364 32768
rect 20824 32728 21364 32756
rect 21358 32716 21364 32728
rect 21416 32716 21422 32768
rect 21729 32759 21787 32765
rect 21729 32725 21741 32759
rect 21775 32756 21787 32759
rect 21818 32756 21824 32768
rect 21775 32728 21824 32756
rect 21775 32725 21787 32728
rect 21729 32719 21787 32725
rect 21818 32716 21824 32728
rect 21876 32716 21882 32768
rect 22833 32759 22891 32765
rect 22833 32725 22845 32759
rect 22879 32756 22891 32759
rect 23014 32756 23020 32768
rect 22879 32728 23020 32756
rect 22879 32725 22891 32728
rect 22833 32719 22891 32725
rect 23014 32716 23020 32728
rect 23072 32716 23078 32768
rect 23106 32716 23112 32768
rect 23164 32756 23170 32768
rect 23382 32756 23388 32768
rect 23164 32728 23388 32756
rect 23164 32716 23170 32728
rect 23382 32716 23388 32728
rect 23440 32756 23446 32768
rect 23753 32759 23811 32765
rect 23753 32756 23765 32759
rect 23440 32728 23765 32756
rect 23440 32716 23446 32728
rect 23753 32725 23765 32728
rect 23799 32725 23811 32759
rect 23753 32719 23811 32725
rect 24486 32716 24492 32768
rect 24544 32756 24550 32768
rect 24673 32759 24731 32765
rect 24673 32756 24685 32759
rect 24544 32728 24685 32756
rect 24544 32716 24550 32728
rect 24673 32725 24685 32728
rect 24719 32725 24731 32759
rect 24780 32756 24808 32796
rect 25041 32793 25053 32827
rect 25087 32824 25099 32827
rect 36648 32824 36676 32855
rect 36814 32852 36820 32864
rect 36872 32852 36878 32904
rect 37550 32892 37556 32904
rect 37511 32864 37556 32892
rect 37550 32852 37556 32864
rect 37608 32852 37614 32904
rect 37660 32901 37688 32932
rect 37645 32895 37703 32901
rect 37645 32861 37657 32895
rect 37691 32861 37703 32895
rect 40218 32892 40224 32904
rect 40179 32864 40224 32892
rect 37645 32855 37703 32861
rect 40218 32852 40224 32864
rect 40276 32852 40282 32904
rect 36722 32824 36728 32836
rect 25087 32796 36728 32824
rect 25087 32793 25099 32796
rect 25041 32787 25099 32793
rect 36722 32784 36728 32796
rect 36780 32784 36786 32836
rect 38654 32824 38660 32836
rect 38615 32796 38660 32824
rect 38654 32784 38660 32796
rect 38712 32784 38718 32836
rect 38930 32833 38936 32836
rect 38873 32827 38936 32833
rect 38873 32793 38885 32827
rect 38919 32793 38936 32827
rect 38873 32787 38936 32793
rect 38930 32784 38936 32787
rect 38988 32784 38994 32836
rect 40037 32827 40095 32833
rect 40037 32824 40049 32827
rect 39040 32796 40049 32824
rect 39040 32768 39068 32796
rect 40037 32793 40049 32796
rect 40083 32793 40095 32827
rect 40037 32787 40095 32793
rect 25958 32756 25964 32768
rect 24780 32728 25964 32756
rect 24673 32719 24731 32725
rect 25958 32716 25964 32728
rect 26016 32716 26022 32768
rect 26605 32759 26663 32765
rect 26605 32725 26617 32759
rect 26651 32756 26663 32759
rect 31110 32756 31116 32768
rect 26651 32728 31116 32756
rect 26651 32725 26663 32728
rect 26605 32719 26663 32725
rect 31110 32716 31116 32728
rect 31168 32716 31174 32768
rect 31294 32716 31300 32768
rect 31352 32756 31358 32768
rect 31754 32756 31760 32768
rect 31352 32728 31760 32756
rect 31352 32716 31358 32728
rect 31754 32716 31760 32728
rect 31812 32756 31818 32768
rect 32766 32756 32772 32768
rect 31812 32728 32772 32756
rect 31812 32716 31818 32728
rect 32766 32716 32772 32728
rect 32824 32716 32830 32768
rect 33594 32756 33600 32768
rect 33555 32728 33600 32756
rect 33594 32716 33600 32728
rect 33652 32716 33658 32768
rect 35618 32716 35624 32768
rect 35676 32756 35682 32768
rect 35805 32759 35863 32765
rect 35805 32756 35817 32759
rect 35676 32728 35817 32756
rect 35676 32716 35682 32728
rect 35805 32725 35817 32728
rect 35851 32725 35863 32759
rect 35805 32719 35863 32725
rect 37829 32759 37887 32765
rect 37829 32725 37841 32759
rect 37875 32756 37887 32759
rect 37918 32756 37924 32768
rect 37875 32728 37924 32756
rect 37875 32725 37887 32728
rect 37829 32719 37887 32725
rect 37918 32716 37924 32728
rect 37976 32716 37982 32768
rect 39022 32716 39028 32768
rect 39080 32756 39086 32768
rect 39080 32728 39173 32756
rect 39080 32716 39086 32728
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 19242 32512 19248 32564
rect 19300 32552 19306 32564
rect 25498 32552 25504 32564
rect 19300 32524 25504 32552
rect 19300 32512 19306 32524
rect 25498 32512 25504 32524
rect 25556 32512 25562 32564
rect 25958 32552 25964 32564
rect 25919 32524 25964 32552
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 26326 32512 26332 32564
rect 26384 32552 26390 32564
rect 26384 32524 28948 32552
rect 26384 32512 26390 32524
rect 20533 32487 20591 32493
rect 20533 32484 20545 32487
rect 19628 32456 20545 32484
rect 18414 32416 18420 32428
rect 18375 32388 18420 32416
rect 18414 32376 18420 32388
rect 18472 32376 18478 32428
rect 19628 32425 19656 32456
rect 20533 32453 20545 32456
rect 20579 32453 20591 32487
rect 24854 32484 24860 32496
rect 24815 32456 24860 32484
rect 20533 32447 20591 32453
rect 24854 32444 24860 32456
rect 24912 32444 24918 32496
rect 25682 32444 25688 32496
rect 25740 32484 25746 32496
rect 25879 32487 25937 32493
rect 25879 32484 25891 32487
rect 25740 32456 25891 32484
rect 25740 32444 25746 32456
rect 25879 32453 25891 32456
rect 25925 32453 25937 32487
rect 27246 32484 27252 32496
rect 27207 32456 27252 32484
rect 25879 32447 25937 32453
rect 27246 32444 27252 32456
rect 27304 32484 27310 32496
rect 27985 32487 28043 32493
rect 27985 32484 27997 32487
rect 27304 32456 27997 32484
rect 27304 32444 27310 32456
rect 27985 32453 27997 32456
rect 28031 32484 28043 32487
rect 28350 32484 28356 32496
rect 28031 32456 28356 32484
rect 28031 32453 28043 32456
rect 27985 32447 28043 32453
rect 28350 32444 28356 32456
rect 28408 32444 28414 32496
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 20438 32416 20444 32428
rect 20399 32388 20444 32416
rect 19613 32379 19671 32385
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 20622 32376 20628 32428
rect 20680 32416 20686 32428
rect 22830 32416 22836 32428
rect 20680 32388 22836 32416
rect 20680 32376 20686 32388
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 22922 32376 22928 32428
rect 22980 32416 22986 32428
rect 23385 32419 23443 32425
rect 23385 32416 23397 32419
rect 22980 32388 23397 32416
rect 22980 32376 22986 32388
rect 23385 32385 23397 32388
rect 23431 32385 23443 32419
rect 23385 32379 23443 32385
rect 15838 32348 15844 32360
rect 15799 32320 15844 32348
rect 15838 32308 15844 32320
rect 15896 32308 15902 32360
rect 18230 32348 18236 32360
rect 18191 32320 18236 32348
rect 18230 32308 18236 32320
rect 18288 32308 18294 32360
rect 19705 32351 19763 32357
rect 19705 32317 19717 32351
rect 19751 32348 19763 32351
rect 23290 32348 23296 32360
rect 19751 32320 23296 32348
rect 19751 32317 19763 32320
rect 19705 32311 19763 32317
rect 23290 32308 23296 32320
rect 23348 32308 23354 32360
rect 15194 32240 15200 32292
rect 15252 32280 15258 32292
rect 15473 32283 15531 32289
rect 15473 32280 15485 32283
rect 15252 32252 15485 32280
rect 15252 32240 15258 32252
rect 15473 32249 15485 32252
rect 15519 32249 15531 32283
rect 15473 32243 15531 32249
rect 15378 32212 15384 32224
rect 15339 32184 15384 32212
rect 15378 32172 15384 32184
rect 15436 32172 15442 32224
rect 18598 32212 18604 32224
rect 18559 32184 18604 32212
rect 18598 32172 18604 32184
rect 18656 32172 18662 32224
rect 19889 32215 19947 32221
rect 19889 32181 19901 32215
rect 19935 32212 19947 32215
rect 19978 32212 19984 32224
rect 19935 32184 19984 32212
rect 19935 32181 19947 32184
rect 19889 32175 19947 32181
rect 19978 32172 19984 32184
rect 20036 32172 20042 32224
rect 21358 32212 21364 32224
rect 21319 32184 21364 32212
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 21450 32172 21456 32224
rect 21508 32212 21514 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 21508 32184 23213 32212
rect 21508 32172 21514 32184
rect 23201 32181 23213 32184
rect 23247 32181 23259 32215
rect 23400 32212 23428 32379
rect 23474 32376 23480 32428
rect 23532 32416 23538 32428
rect 23532 32388 23577 32416
rect 23532 32376 23538 32388
rect 23658 32376 23664 32428
rect 23716 32416 23722 32428
rect 24581 32419 24639 32425
rect 23716 32388 23761 32416
rect 23716 32376 23722 32388
rect 24581 32385 24593 32419
rect 24627 32416 24639 32419
rect 24670 32416 24676 32428
rect 24627 32388 24676 32416
rect 24627 32385 24639 32388
rect 24581 32379 24639 32385
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32385 25007 32419
rect 25774 32416 25780 32428
rect 25735 32388 25780 32416
rect 24949 32379 25007 32385
rect 23566 32348 23572 32360
rect 23527 32320 23572 32348
rect 23566 32308 23572 32320
rect 23624 32308 23630 32360
rect 24486 32348 24492 32360
rect 24447 32320 24492 32348
rect 24486 32308 24492 32320
rect 24544 32308 24550 32360
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 24964 32348 24992 32379
rect 25774 32376 25780 32388
rect 25832 32376 25838 32428
rect 26145 32419 26203 32425
rect 26145 32385 26157 32419
rect 26191 32416 26203 32419
rect 26602 32416 26608 32428
rect 26191 32388 26608 32416
rect 26191 32385 26203 32388
rect 26145 32379 26203 32385
rect 26602 32376 26608 32388
rect 26660 32376 26666 32428
rect 27430 32416 27436 32428
rect 27391 32388 27436 32416
rect 27430 32376 27436 32388
rect 27488 32376 27494 32428
rect 27522 32376 27528 32428
rect 27580 32416 27586 32428
rect 28810 32416 28816 32428
rect 27580 32388 27625 32416
rect 28771 32388 28816 32416
rect 27580 32376 27586 32388
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 28920 32416 28948 32524
rect 30282 32512 30288 32564
rect 30340 32552 30346 32564
rect 30469 32555 30527 32561
rect 30469 32552 30481 32555
rect 30340 32524 30481 32552
rect 30340 32512 30346 32524
rect 30469 32521 30481 32524
rect 30515 32521 30527 32555
rect 30469 32515 30527 32521
rect 31757 32555 31815 32561
rect 31757 32521 31769 32555
rect 31803 32552 31815 32555
rect 35253 32555 35311 32561
rect 35253 32552 35265 32555
rect 31803 32524 35265 32552
rect 31803 32521 31815 32524
rect 31757 32515 31815 32521
rect 35253 32521 35265 32524
rect 35299 32521 35311 32555
rect 35253 32515 35311 32521
rect 30650 32484 30656 32496
rect 30392 32456 30656 32484
rect 28997 32419 29055 32425
rect 28997 32416 29009 32419
rect 28920 32388 29009 32416
rect 28997 32385 29009 32388
rect 29043 32416 29055 32419
rect 29362 32416 29368 32428
rect 29043 32388 29368 32416
rect 29043 32385 29055 32388
rect 28997 32379 29055 32385
rect 29362 32376 29368 32388
rect 29420 32416 29426 32428
rect 29457 32419 29515 32425
rect 29457 32416 29469 32419
rect 29420 32388 29469 32416
rect 29420 32376 29426 32388
rect 29457 32385 29469 32388
rect 29503 32385 29515 32419
rect 30392 32416 30420 32456
rect 30650 32444 30656 32456
rect 30708 32444 30714 32496
rect 32769 32487 32827 32493
rect 32769 32453 32781 32487
rect 32815 32484 32827 32487
rect 32815 32456 33732 32484
rect 32815 32453 32827 32456
rect 32769 32447 32827 32453
rect 31202 32416 31208 32428
rect 29457 32379 29515 32385
rect 30208 32388 30420 32416
rect 30852 32388 31208 32416
rect 29086 32348 29092 32360
rect 24820 32320 29092 32348
rect 24820 32308 24826 32320
rect 29086 32308 29092 32320
rect 29144 32308 29150 32360
rect 30208 32357 30236 32388
rect 30193 32351 30251 32357
rect 30193 32317 30205 32351
rect 30239 32317 30251 32351
rect 30374 32348 30380 32360
rect 30335 32320 30380 32348
rect 30193 32311 30251 32317
rect 30374 32308 30380 32320
rect 30432 32308 30438 32360
rect 25593 32283 25651 32289
rect 25593 32249 25605 32283
rect 25639 32280 25651 32283
rect 25682 32280 25688 32292
rect 25639 32252 25688 32280
rect 25639 32249 25651 32252
rect 25593 32243 25651 32249
rect 25682 32240 25688 32252
rect 25740 32240 25746 32292
rect 28813 32283 28871 32289
rect 28813 32249 28825 32283
rect 28859 32280 28871 32283
rect 30466 32280 30472 32292
rect 28859 32252 30472 32280
rect 28859 32249 28871 32252
rect 28813 32243 28871 32249
rect 30466 32240 30472 32252
rect 30524 32240 30530 32292
rect 30852 32289 30880 32388
rect 31202 32376 31208 32388
rect 31260 32416 31266 32428
rect 31297 32419 31355 32425
rect 31297 32416 31309 32419
rect 31260 32388 31309 32416
rect 31260 32376 31266 32388
rect 31297 32385 31309 32388
rect 31343 32385 31355 32419
rect 31297 32379 31355 32385
rect 32674 32376 32680 32428
rect 32732 32416 32738 32428
rect 32953 32419 33011 32425
rect 32953 32416 32965 32419
rect 32732 32388 32965 32416
rect 32732 32376 32738 32388
rect 32953 32385 32965 32388
rect 32999 32385 33011 32419
rect 32953 32379 33011 32385
rect 33045 32419 33103 32425
rect 33045 32385 33057 32419
rect 33091 32416 33103 32419
rect 33226 32416 33232 32428
rect 33091 32388 33232 32416
rect 33091 32385 33103 32388
rect 33045 32379 33103 32385
rect 33226 32376 33232 32388
rect 33284 32376 33290 32428
rect 33594 32416 33600 32428
rect 33555 32388 33600 32416
rect 33594 32376 33600 32388
rect 33652 32376 33658 32428
rect 33704 32425 33732 32456
rect 33689 32419 33747 32425
rect 33689 32385 33701 32419
rect 33735 32416 33747 32419
rect 33778 32416 33784 32428
rect 33735 32388 33784 32416
rect 33735 32385 33747 32388
rect 33689 32379 33747 32385
rect 33778 32376 33784 32388
rect 33836 32376 33842 32428
rect 33965 32419 34023 32425
rect 33965 32385 33977 32419
rect 34011 32385 34023 32419
rect 33965 32379 34023 32385
rect 32122 32308 32128 32360
rect 32180 32348 32186 32360
rect 32769 32351 32827 32357
rect 32769 32348 32781 32351
rect 32180 32320 32781 32348
rect 32180 32308 32186 32320
rect 32769 32317 32781 32320
rect 32815 32317 32827 32351
rect 32769 32311 32827 32317
rect 33502 32308 33508 32360
rect 33560 32348 33566 32360
rect 33980 32348 34008 32379
rect 34054 32376 34060 32428
rect 34112 32416 34118 32428
rect 34333 32419 34391 32425
rect 34333 32416 34345 32419
rect 34112 32388 34345 32416
rect 34112 32376 34118 32388
rect 34333 32385 34345 32388
rect 34379 32385 34391 32419
rect 34333 32379 34391 32385
rect 35161 32419 35219 32425
rect 35161 32385 35173 32419
rect 35207 32385 35219 32419
rect 35161 32379 35219 32385
rect 33560 32320 34008 32348
rect 33560 32308 33566 32320
rect 30837 32283 30895 32289
rect 30837 32249 30849 32283
rect 30883 32249 30895 32283
rect 30837 32243 30895 32249
rect 33686 32240 33692 32292
rect 33744 32280 33750 32292
rect 34072 32280 34100 32376
rect 34149 32351 34207 32357
rect 34149 32317 34161 32351
rect 34195 32348 34207 32351
rect 34422 32348 34428 32360
rect 34195 32320 34428 32348
rect 34195 32317 34207 32320
rect 34149 32311 34207 32317
rect 34422 32308 34428 32320
rect 34480 32348 34486 32360
rect 35176 32348 35204 32379
rect 34480 32320 35204 32348
rect 35268 32348 35296 32515
rect 35986 32512 35992 32564
rect 36044 32552 36050 32564
rect 36081 32555 36139 32561
rect 36081 32552 36093 32555
rect 36044 32524 36093 32552
rect 36044 32512 36050 32524
rect 36081 32521 36093 32524
rect 36127 32521 36139 32555
rect 39577 32555 39635 32561
rect 36081 32515 36139 32521
rect 37476 32524 39160 32552
rect 36357 32487 36415 32493
rect 36357 32484 36369 32487
rect 35728 32456 36369 32484
rect 35728 32428 35756 32456
rect 36357 32453 36369 32456
rect 36403 32453 36415 32487
rect 36357 32447 36415 32453
rect 35437 32419 35495 32425
rect 35437 32385 35449 32419
rect 35483 32416 35495 32419
rect 35710 32416 35716 32428
rect 35483 32388 35716 32416
rect 35483 32385 35495 32388
rect 35437 32379 35495 32385
rect 35710 32376 35716 32388
rect 35768 32376 35774 32428
rect 36081 32419 36139 32425
rect 36081 32385 36093 32419
rect 36127 32385 36139 32419
rect 36081 32379 36139 32385
rect 36173 32419 36231 32425
rect 36173 32385 36185 32419
rect 36219 32385 36231 32419
rect 36173 32379 36231 32385
rect 36096 32348 36124 32379
rect 35268 32320 36124 32348
rect 34480 32308 34486 32320
rect 33744 32252 34100 32280
rect 35176 32280 35204 32320
rect 36188 32280 36216 32379
rect 37476 32348 37504 32524
rect 38746 32484 38752 32496
rect 38580 32456 38752 32484
rect 37642 32416 37648 32428
rect 37603 32388 37648 32416
rect 37642 32376 37648 32388
rect 37700 32376 37706 32428
rect 37918 32416 37924 32428
rect 37879 32388 37924 32416
rect 37918 32376 37924 32388
rect 37976 32376 37982 32428
rect 38580 32425 38608 32456
rect 38746 32444 38752 32456
rect 38804 32444 38810 32496
rect 39132 32484 39160 32524
rect 39577 32521 39589 32555
rect 39623 32552 39635 32555
rect 39666 32552 39672 32564
rect 39623 32524 39672 32552
rect 39623 32521 39635 32524
rect 39577 32515 39635 32521
rect 39666 32512 39672 32524
rect 39724 32512 39730 32564
rect 39132 32456 39620 32484
rect 38565 32419 38623 32425
rect 38565 32385 38577 32419
rect 38611 32385 38623 32419
rect 38565 32379 38623 32385
rect 38841 32419 38899 32425
rect 38841 32385 38853 32419
rect 38887 32416 38899 32419
rect 39022 32416 39028 32428
rect 38887 32388 39028 32416
rect 38887 32385 38899 32388
rect 38841 32379 38899 32385
rect 39022 32376 39028 32388
rect 39080 32376 39086 32428
rect 35176 32252 36216 32280
rect 36372 32320 37504 32348
rect 38657 32351 38715 32357
rect 38657 32340 38669 32351
rect 33744 32240 33750 32252
rect 26970 32212 26976 32224
rect 23400 32184 26976 32212
rect 23201 32175 23259 32181
rect 26970 32172 26976 32184
rect 27028 32172 27034 32224
rect 27246 32212 27252 32224
rect 27207 32184 27252 32212
rect 27246 32172 27252 32184
rect 27304 32172 27310 32224
rect 31110 32172 31116 32224
rect 31168 32212 31174 32224
rect 31389 32215 31447 32221
rect 31389 32212 31401 32215
rect 31168 32184 31401 32212
rect 31168 32172 31174 32184
rect 31389 32181 31401 32184
rect 31435 32181 31447 32215
rect 31389 32175 31447 32181
rect 33594 32172 33600 32224
rect 33652 32212 33658 32224
rect 33870 32212 33876 32224
rect 33652 32184 33876 32212
rect 33652 32172 33658 32184
rect 33870 32172 33876 32184
rect 33928 32172 33934 32224
rect 35621 32215 35679 32221
rect 35621 32181 35633 32215
rect 35667 32212 35679 32215
rect 35802 32212 35808 32224
rect 35667 32184 35808 32212
rect 35667 32181 35679 32184
rect 35621 32175 35679 32181
rect 35802 32172 35808 32184
rect 35860 32212 35866 32224
rect 36372 32212 36400 32320
rect 38580 32317 38669 32340
rect 38703 32317 38715 32351
rect 38580 32312 38715 32317
rect 36446 32240 36452 32292
rect 36504 32280 36510 32292
rect 38580 32280 38608 32312
rect 38657 32311 38715 32312
rect 38749 32351 38807 32357
rect 38749 32317 38761 32351
rect 38795 32348 38807 32351
rect 39132 32348 39160 32456
rect 39592 32425 39620 32456
rect 39393 32419 39451 32425
rect 39393 32385 39405 32419
rect 39439 32385 39451 32419
rect 39393 32379 39451 32385
rect 39577 32419 39635 32425
rect 39577 32385 39589 32419
rect 39623 32385 39635 32419
rect 39577 32379 39635 32385
rect 38795 32320 39160 32348
rect 38795 32317 38807 32320
rect 38749 32311 38807 32317
rect 39408 32280 39436 32379
rect 36504 32252 39436 32280
rect 36504 32240 36510 32252
rect 37458 32212 37464 32224
rect 35860 32184 36400 32212
rect 37419 32184 37464 32212
rect 35860 32172 35866 32184
rect 37458 32172 37464 32184
rect 37516 32172 37522 32224
rect 37829 32215 37887 32221
rect 37829 32181 37841 32215
rect 37875 32212 37887 32215
rect 38381 32215 38439 32221
rect 38381 32212 38393 32215
rect 37875 32184 38393 32212
rect 37875 32181 37887 32184
rect 37829 32175 37887 32181
rect 38381 32181 38393 32184
rect 38427 32181 38439 32215
rect 38381 32175 38439 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 18230 31968 18236 32020
rect 18288 32008 18294 32020
rect 22005 32011 22063 32017
rect 22005 32008 22017 32011
rect 18288 31980 22017 32008
rect 18288 31968 18294 31980
rect 22005 31977 22017 31980
rect 22051 31977 22063 32011
rect 22005 31971 22063 31977
rect 23658 31968 23664 32020
rect 23716 32008 23722 32020
rect 24581 32011 24639 32017
rect 24581 32008 24593 32011
rect 23716 31980 24593 32008
rect 23716 31968 23722 31980
rect 24581 31977 24593 31980
rect 24627 31977 24639 32011
rect 24581 31971 24639 31977
rect 24670 31968 24676 32020
rect 24728 32008 24734 32020
rect 24949 32011 25007 32017
rect 24949 32008 24961 32011
rect 24728 31980 24961 32008
rect 24728 31968 24734 31980
rect 24949 31977 24961 31980
rect 24995 31977 25007 32011
rect 26970 32008 26976 32020
rect 26931 31980 26976 32008
rect 24949 31971 25007 31977
rect 26970 31968 26976 31980
rect 27028 31968 27034 32020
rect 28350 32008 28356 32020
rect 28311 31980 28356 32008
rect 28350 31968 28356 31980
rect 28408 31968 28414 32020
rect 30374 32008 30380 32020
rect 30335 31980 30380 32008
rect 30374 31968 30380 31980
rect 30432 31968 30438 32020
rect 30466 31968 30472 32020
rect 30524 32008 30530 32020
rect 30524 31980 35388 32008
rect 30524 31968 30530 31980
rect 18046 31940 18052 31952
rect 16960 31912 18052 31940
rect 16666 31872 16672 31884
rect 16627 31844 16672 31872
rect 16666 31832 16672 31844
rect 16724 31832 16730 31884
rect 16960 31881 16988 31912
rect 18046 31900 18052 31912
rect 18104 31900 18110 31952
rect 25774 31940 25780 31952
rect 19996 31912 21128 31940
rect 19996 31884 20024 31912
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31841 17003 31875
rect 17678 31872 17684 31884
rect 16945 31835 17003 31841
rect 17052 31844 17684 31872
rect 15286 31804 15292 31816
rect 15247 31776 15292 31804
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 15378 31764 15384 31816
rect 15436 31804 15442 31816
rect 17052 31813 17080 31844
rect 17678 31832 17684 31844
rect 17736 31872 17742 31884
rect 18598 31872 18604 31884
rect 17736 31844 18276 31872
rect 18559 31844 18604 31872
rect 17736 31832 17742 31844
rect 15749 31807 15807 31813
rect 15749 31804 15761 31807
rect 15436 31776 15761 31804
rect 15436 31764 15442 31776
rect 15749 31773 15761 31776
rect 15795 31773 15807 31807
rect 15749 31767 15807 31773
rect 17037 31807 17095 31813
rect 17037 31773 17049 31807
rect 17083 31773 17095 31807
rect 18046 31804 18052 31816
rect 18007 31776 18052 31804
rect 17037 31767 17095 31773
rect 18046 31764 18052 31776
rect 18104 31764 18110 31816
rect 18248 31813 18276 31844
rect 18598 31832 18604 31844
rect 18656 31832 18662 31884
rect 19978 31872 19984 31884
rect 19939 31844 19984 31872
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 20438 31872 20444 31884
rect 20399 31844 20444 31872
rect 20438 31832 20444 31844
rect 20496 31832 20502 31884
rect 18233 31807 18291 31813
rect 18233 31773 18245 31807
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 20073 31807 20131 31813
rect 20073 31773 20085 31807
rect 20119 31804 20131 31807
rect 20898 31804 20904 31816
rect 20119 31776 20760 31804
rect 20859 31776 20904 31804
rect 20119 31773 20131 31776
rect 20073 31767 20131 31773
rect 14648 31748 14700 31754
rect 20732 31736 20760 31776
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 21100 31813 21128 31912
rect 24872 31912 25780 31940
rect 23109 31875 23167 31881
rect 23109 31841 23121 31875
rect 23155 31872 23167 31875
rect 24872 31872 24900 31912
rect 25774 31900 25780 31912
rect 25832 31900 25838 31952
rect 26878 31940 26884 31952
rect 26791 31912 26884 31940
rect 26878 31900 26884 31912
rect 26936 31940 26942 31952
rect 27246 31940 27252 31952
rect 26936 31912 27252 31940
rect 26936 31900 26942 31912
rect 27246 31900 27252 31912
rect 27304 31900 27310 31952
rect 31665 31943 31723 31949
rect 31665 31909 31677 31943
rect 31711 31940 31723 31943
rect 35360 31940 35388 31980
rect 35434 31968 35440 32020
rect 35492 32008 35498 32020
rect 36081 32011 36139 32017
rect 36081 32008 36093 32011
rect 35492 31980 36093 32008
rect 35492 31968 35498 31980
rect 36081 31977 36093 31980
rect 36127 31977 36139 32011
rect 37642 32008 37648 32020
rect 37603 31980 37648 32008
rect 36081 31971 36139 31977
rect 37642 31968 37648 31980
rect 37700 31968 37706 32020
rect 37550 31940 37556 31952
rect 31711 31912 33180 31940
rect 35360 31912 37556 31940
rect 31711 31909 31723 31912
rect 31665 31903 31723 31909
rect 23155 31844 24900 31872
rect 23155 31841 23167 31844
rect 23109 31835 23167 31841
rect 25866 31832 25872 31884
rect 25924 31872 25930 31884
rect 27154 31872 27160 31884
rect 25924 31844 27160 31872
rect 25924 31832 25930 31844
rect 27154 31832 27160 31844
rect 27212 31872 27218 31884
rect 27525 31875 27583 31881
rect 27525 31872 27537 31875
rect 27212 31844 27537 31872
rect 27212 31832 27218 31844
rect 27525 31841 27537 31844
rect 27571 31841 27583 31875
rect 30558 31872 30564 31884
rect 27525 31835 27583 31841
rect 30484 31844 30564 31872
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21269 31807 21327 31813
rect 21269 31804 21281 31807
rect 21085 31767 21143 31773
rect 21192 31776 21281 31804
rect 21192 31736 21220 31776
rect 21269 31773 21281 31776
rect 21315 31804 21327 31807
rect 21450 31804 21456 31816
rect 21315 31776 21456 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21450 31764 21456 31776
rect 21508 31764 21514 31816
rect 21726 31804 21732 31816
rect 21687 31776 21732 31804
rect 21726 31764 21732 31776
rect 21784 31764 21790 31816
rect 22005 31807 22063 31813
rect 22005 31773 22017 31807
rect 22051 31804 22063 31807
rect 22278 31804 22284 31816
rect 22051 31776 22284 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 22278 31764 22284 31776
rect 22336 31764 22342 31816
rect 23014 31804 23020 31816
rect 22975 31776 23020 31804
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 24762 31804 24768 31816
rect 24723 31776 24768 31804
rect 24762 31764 24768 31776
rect 24820 31764 24826 31816
rect 25041 31807 25099 31813
rect 25041 31773 25053 31807
rect 25087 31773 25099 31807
rect 25041 31767 25099 31773
rect 20732 31708 21220 31736
rect 21634 31696 21640 31748
rect 21692 31736 21698 31748
rect 21821 31739 21879 31745
rect 21821 31736 21833 31739
rect 21692 31708 21833 31736
rect 21692 31696 21698 31708
rect 21821 31705 21833 31708
rect 21867 31705 21879 31739
rect 21821 31699 21879 31705
rect 24486 31696 24492 31748
rect 24544 31736 24550 31748
rect 25056 31736 25084 31767
rect 25314 31764 25320 31816
rect 25372 31804 25378 31816
rect 25501 31807 25559 31813
rect 25501 31804 25513 31807
rect 25372 31776 25513 31804
rect 25372 31764 25378 31776
rect 25501 31773 25513 31776
rect 25547 31773 25559 31807
rect 25501 31767 25559 31773
rect 25590 31764 25596 31816
rect 25648 31804 25654 31816
rect 25685 31807 25743 31813
rect 25685 31804 25697 31807
rect 25648 31776 25697 31804
rect 25648 31764 25654 31776
rect 25685 31773 25697 31776
rect 25731 31804 25743 31807
rect 26326 31804 26332 31816
rect 25731 31776 26332 31804
rect 25731 31773 25743 31776
rect 25685 31767 25743 31773
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 26970 31764 26976 31816
rect 27028 31804 27034 31816
rect 30484 31813 30512 31844
rect 30558 31832 30564 31844
rect 30616 31832 30622 31884
rect 31202 31872 31208 31884
rect 31163 31844 31208 31872
rect 31202 31832 31208 31844
rect 31260 31832 31266 31884
rect 32950 31872 32956 31884
rect 32508 31844 32956 31872
rect 30469 31807 30527 31813
rect 30469 31804 30481 31807
rect 27028 31776 27073 31804
rect 30392 31776 30481 31804
rect 27028 31764 27034 31776
rect 25866 31736 25872 31748
rect 24544 31708 25872 31736
rect 24544 31696 24550 31708
rect 25866 31696 25872 31708
rect 25924 31696 25930 31748
rect 26237 31739 26295 31745
rect 26237 31705 26249 31739
rect 26283 31736 26295 31739
rect 26697 31739 26755 31745
rect 26697 31736 26709 31739
rect 26283 31708 26709 31736
rect 26283 31705 26295 31708
rect 26237 31699 26295 31705
rect 26697 31705 26709 31708
rect 26743 31736 26755 31739
rect 27062 31736 27068 31748
rect 26743 31708 27068 31736
rect 26743 31705 26755 31708
rect 26697 31699 26755 31705
rect 27062 31696 27068 31708
rect 27120 31696 27126 31748
rect 27798 31736 27804 31748
rect 27759 31708 27804 31736
rect 27798 31696 27804 31708
rect 27856 31696 27862 31748
rect 29178 31696 29184 31748
rect 29236 31736 29242 31748
rect 30392 31736 30420 31776
rect 30469 31773 30481 31776
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 31110 31764 31116 31816
rect 31168 31804 31174 31816
rect 32508 31813 32536 31844
rect 32950 31832 32956 31844
rect 33008 31832 33014 31884
rect 31297 31807 31355 31813
rect 31297 31804 31309 31807
rect 31168 31776 31309 31804
rect 31168 31764 31174 31776
rect 31297 31773 31309 31776
rect 31343 31773 31355 31807
rect 31297 31767 31355 31773
rect 32493 31807 32551 31813
rect 32493 31773 32505 31807
rect 32539 31773 32551 31807
rect 32674 31804 32680 31816
rect 32635 31776 32680 31804
rect 32493 31767 32551 31773
rect 32674 31764 32680 31776
rect 32732 31764 32738 31816
rect 33152 31804 33180 31912
rect 33778 31872 33784 31884
rect 33739 31844 33784 31872
rect 33778 31832 33784 31844
rect 33836 31832 33842 31884
rect 33870 31832 33876 31884
rect 33928 31872 33934 31884
rect 33928 31844 33973 31872
rect 33928 31832 33934 31844
rect 34054 31832 34060 31884
rect 34112 31872 34118 31884
rect 34885 31875 34943 31881
rect 34885 31872 34897 31875
rect 34112 31844 34897 31872
rect 34112 31832 34118 31844
rect 34885 31841 34897 31844
rect 34931 31841 34943 31875
rect 34885 31835 34943 31841
rect 35529 31875 35587 31881
rect 35529 31841 35541 31875
rect 35575 31872 35587 31875
rect 36446 31872 36452 31884
rect 35575 31844 36308 31872
rect 36407 31844 36452 31872
rect 35575 31841 35587 31844
rect 35529 31835 35587 31841
rect 33502 31804 33508 31816
rect 33152 31776 33508 31804
rect 33502 31764 33508 31776
rect 33560 31804 33566 31816
rect 33597 31807 33655 31813
rect 33597 31804 33609 31807
rect 33560 31776 33609 31804
rect 33560 31764 33566 31776
rect 33597 31773 33609 31776
rect 33643 31773 33655 31807
rect 33597 31767 33655 31773
rect 33689 31807 33747 31813
rect 33689 31773 33701 31807
rect 33735 31804 33747 31807
rect 34072 31804 34100 31832
rect 35434 31804 35440 31816
rect 33735 31776 34100 31804
rect 35395 31776 35440 31804
rect 33735 31773 33747 31776
rect 33689 31767 33747 31773
rect 35434 31764 35440 31776
rect 35492 31764 35498 31816
rect 35618 31804 35624 31816
rect 35579 31776 35624 31804
rect 35618 31764 35624 31776
rect 35676 31764 35682 31816
rect 36280 31813 36308 31844
rect 36446 31832 36452 31844
rect 36504 31832 36510 31884
rect 36265 31807 36323 31813
rect 36265 31773 36277 31807
rect 36311 31773 36323 31807
rect 37274 31804 37280 31816
rect 37235 31776 37280 31804
rect 36265 31767 36323 31773
rect 37274 31764 37280 31776
rect 37332 31764 37338 31816
rect 37476 31813 37504 31912
rect 37550 31900 37556 31912
rect 37608 31900 37614 31952
rect 37461 31807 37519 31813
rect 37461 31773 37473 31807
rect 37507 31773 37519 31807
rect 37461 31767 37519 31773
rect 29236 31708 30420 31736
rect 29236 31696 29242 31708
rect 14648 31690 14700 31696
rect 18506 31668 18512 31680
rect 18467 31640 18512 31668
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 22649 31671 22707 31677
rect 22649 31637 22661 31671
rect 22695 31668 22707 31671
rect 22738 31668 22744 31680
rect 22695 31640 22744 31668
rect 22695 31637 22707 31640
rect 22649 31631 22707 31637
rect 22738 31628 22744 31640
rect 22796 31628 22802 31680
rect 25685 31671 25743 31677
rect 25685 31637 25697 31671
rect 25731 31668 25743 31671
rect 26050 31668 26056 31680
rect 25731 31640 26056 31668
rect 25731 31637 25743 31640
rect 25685 31631 25743 31637
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 26510 31628 26516 31680
rect 26568 31668 26574 31680
rect 28626 31668 28632 31680
rect 26568 31640 28632 31668
rect 26568 31628 26574 31640
rect 28626 31628 28632 31640
rect 28684 31628 28690 31680
rect 32582 31668 32588 31680
rect 32543 31640 32588 31668
rect 32582 31628 32588 31640
rect 32640 31628 32646 31680
rect 34054 31668 34060 31680
rect 34015 31640 34060 31668
rect 34054 31628 34060 31640
rect 34112 31628 34118 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 15565 31467 15623 31473
rect 15565 31464 15577 31467
rect 15120 31436 15577 31464
rect 15120 31405 15148 31436
rect 15565 31433 15577 31436
rect 15611 31464 15623 31467
rect 15838 31464 15844 31476
rect 15611 31436 15844 31464
rect 15611 31433 15623 31436
rect 15565 31427 15623 31433
rect 15838 31424 15844 31436
rect 15896 31424 15902 31476
rect 21634 31424 21640 31476
rect 21692 31464 21698 31476
rect 22097 31467 22155 31473
rect 22097 31464 22109 31467
rect 21692 31436 22109 31464
rect 21692 31424 21698 31436
rect 22097 31433 22109 31436
rect 22143 31464 22155 31467
rect 24486 31464 24492 31476
rect 22143 31436 24492 31464
rect 22143 31433 22155 31436
rect 22097 31427 22155 31433
rect 24486 31424 24492 31436
rect 24544 31464 24550 31476
rect 24765 31467 24823 31473
rect 24765 31464 24777 31467
rect 24544 31436 24777 31464
rect 24544 31424 24550 31436
rect 24765 31433 24777 31436
rect 24811 31433 24823 31467
rect 24765 31427 24823 31433
rect 26970 31424 26976 31476
rect 27028 31464 27034 31476
rect 27249 31467 27307 31473
rect 27249 31464 27261 31467
rect 27028 31436 27261 31464
rect 27028 31424 27034 31436
rect 27249 31433 27261 31436
rect 27295 31433 27307 31467
rect 28077 31467 28135 31473
rect 28077 31464 28089 31467
rect 27249 31427 27307 31433
rect 27356 31436 28089 31464
rect 15105 31399 15163 31405
rect 15105 31365 15117 31399
rect 15151 31365 15163 31399
rect 16666 31396 16672 31408
rect 15105 31359 15163 31365
rect 15764 31368 16672 31396
rect 14829 31331 14887 31337
rect 14829 31297 14841 31331
rect 14875 31297 14887 31331
rect 14829 31291 14887 31297
rect 14921 31331 14979 31337
rect 14921 31297 14933 31331
rect 14967 31328 14979 31331
rect 15194 31328 15200 31340
rect 14967 31300 15200 31328
rect 14967 31297 14979 31300
rect 14921 31291 14979 31297
rect 14844 31260 14872 31291
rect 15194 31288 15200 31300
rect 15252 31288 15258 31340
rect 15764 31337 15792 31368
rect 16666 31356 16672 31368
rect 16724 31356 16730 31408
rect 27356 31396 27384 31436
rect 28077 31433 28089 31436
rect 28123 31433 28135 31467
rect 32674 31464 32680 31476
rect 32635 31436 32680 31464
rect 28077 31427 28135 31433
rect 32674 31424 32680 31436
rect 32732 31464 32738 31476
rect 32732 31436 33364 31464
rect 32732 31424 32738 31436
rect 27430 31405 27436 31408
rect 24872 31368 27384 31396
rect 27417 31399 27436 31405
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 15930 31328 15936 31340
rect 15891 31300 15936 31328
rect 15749 31291 15807 31297
rect 15930 31288 15936 31300
rect 15988 31288 15994 31340
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16114 31328 16120 31340
rect 16071 31300 16120 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16114 31288 16120 31300
rect 16172 31288 16178 31340
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31328 18107 31331
rect 18230 31328 18236 31340
rect 18095 31300 18236 31328
rect 18095 31297 18107 31300
rect 18049 31291 18107 31297
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 22002 31328 22008 31340
rect 21963 31300 22008 31328
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 22278 31328 22284 31340
rect 22239 31300 22284 31328
rect 22278 31288 22284 31300
rect 22336 31328 22342 31340
rect 24581 31331 24639 31337
rect 24581 31328 24593 31331
rect 22336 31300 24593 31328
rect 22336 31288 22342 31300
rect 24581 31297 24593 31300
rect 24627 31328 24639 31331
rect 24762 31328 24768 31340
rect 24627 31300 24768 31328
rect 24627 31297 24639 31300
rect 24581 31291 24639 31297
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 24872 31337 24900 31368
rect 27417 31365 27429 31399
rect 27417 31359 27436 31365
rect 27430 31356 27436 31359
rect 27488 31356 27494 31408
rect 27614 31396 27620 31408
rect 27575 31368 27620 31396
rect 27614 31356 27620 31368
rect 27672 31356 27678 31408
rect 30837 31399 30895 31405
rect 30837 31396 30849 31399
rect 28368 31368 30849 31396
rect 24857 31331 24915 31337
rect 24857 31297 24869 31331
rect 24903 31297 24915 31331
rect 25866 31328 25872 31340
rect 25827 31300 25872 31328
rect 24857 31291 24915 31297
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 26050 31328 26056 31340
rect 26011 31300 26056 31328
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 28368 31328 28396 31368
rect 30837 31365 30849 31368
rect 30883 31396 30895 31399
rect 31386 31396 31392 31408
rect 30883 31368 31392 31396
rect 30883 31365 30895 31368
rect 30837 31359 30895 31365
rect 31386 31356 31392 31368
rect 31444 31356 31450 31408
rect 32950 31356 32956 31408
rect 33008 31396 33014 31408
rect 33336 31405 33364 31436
rect 34054 31424 34060 31476
rect 34112 31464 34118 31476
rect 34349 31467 34407 31473
rect 34349 31464 34361 31467
rect 34112 31436 34361 31464
rect 34112 31424 34118 31436
rect 34349 31433 34361 31436
rect 34395 31433 34407 31467
rect 34349 31427 34407 31433
rect 34517 31467 34575 31473
rect 34517 31433 34529 31467
rect 34563 31464 34575 31467
rect 34563 31436 36768 31464
rect 34563 31433 34575 31436
rect 34517 31427 34575 31433
rect 33137 31399 33195 31405
rect 33137 31396 33149 31399
rect 33008 31368 33149 31396
rect 33008 31356 33014 31368
rect 33137 31365 33149 31368
rect 33183 31365 33195 31399
rect 33137 31359 33195 31365
rect 33321 31399 33379 31405
rect 33321 31365 33333 31399
rect 33367 31365 33379 31399
rect 33321 31359 33379 31365
rect 34149 31399 34207 31405
rect 34149 31365 34161 31399
rect 34195 31396 34207 31399
rect 34238 31396 34244 31408
rect 34195 31368 34244 31396
rect 34195 31365 34207 31368
rect 34149 31359 34207 31365
rect 34238 31356 34244 31368
rect 34296 31356 34302 31408
rect 36740 31405 36768 31436
rect 36725 31399 36783 31405
rect 36725 31365 36737 31399
rect 36771 31365 36783 31399
rect 36725 31359 36783 31365
rect 26252 31300 28396 31328
rect 28445 31331 28503 31337
rect 15286 31260 15292 31272
rect 14844 31232 15292 31260
rect 15286 31220 15292 31232
rect 15344 31220 15350 31272
rect 17678 31260 17684 31272
rect 17639 31232 17684 31260
rect 17678 31220 17684 31232
rect 17736 31220 17742 31272
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31260 18199 31263
rect 18414 31260 18420 31272
rect 18187 31232 18420 31260
rect 18187 31229 18199 31232
rect 18141 31223 18199 31229
rect 18414 31220 18420 31232
rect 18472 31220 18478 31272
rect 24780 31260 24808 31288
rect 25777 31263 25835 31269
rect 25777 31260 25789 31263
rect 24780 31232 25789 31260
rect 25777 31229 25789 31232
rect 25823 31229 25835 31263
rect 25958 31260 25964 31272
rect 25919 31232 25964 31260
rect 25777 31223 25835 31229
rect 25958 31220 25964 31232
rect 26016 31220 26022 31272
rect 26252 31269 26280 31300
rect 28445 31297 28457 31331
rect 28491 31328 28503 31331
rect 28626 31328 28632 31340
rect 28491 31300 28632 31328
rect 28491 31297 28503 31300
rect 28445 31291 28503 31297
rect 28626 31288 28632 31300
rect 28684 31288 28690 31340
rect 29178 31328 29184 31340
rect 29139 31300 29184 31328
rect 29178 31288 29184 31300
rect 29236 31288 29242 31340
rect 29638 31288 29644 31340
rect 29696 31288 29702 31340
rect 31018 31328 31024 31340
rect 30979 31300 31024 31328
rect 31018 31288 31024 31300
rect 31076 31288 31082 31340
rect 31478 31288 31484 31340
rect 31536 31328 31542 31340
rect 32493 31331 32551 31337
rect 32493 31328 32505 31331
rect 31536 31300 32505 31328
rect 31536 31288 31542 31300
rect 32493 31297 32505 31300
rect 32539 31297 32551 31331
rect 35342 31328 35348 31340
rect 35303 31300 35348 31328
rect 32493 31291 32551 31297
rect 35342 31288 35348 31300
rect 35400 31288 35406 31340
rect 35894 31288 35900 31340
rect 35952 31328 35958 31340
rect 36541 31331 36599 31337
rect 36541 31328 36553 31331
rect 35952 31300 36553 31328
rect 35952 31288 35958 31300
rect 36541 31297 36553 31300
rect 36587 31297 36599 31331
rect 36541 31291 36599 31297
rect 26237 31263 26295 31269
rect 26237 31229 26249 31263
rect 26283 31229 26295 31263
rect 28534 31260 28540 31272
rect 28495 31232 28540 31260
rect 26237 31223 26295 31229
rect 28534 31220 28540 31232
rect 28592 31220 28598 31272
rect 30098 31260 30104 31272
rect 30059 31232 30104 31260
rect 30098 31220 30104 31232
rect 30156 31220 30162 31272
rect 31205 31263 31263 31269
rect 31205 31229 31217 31263
rect 31251 31260 31263 31263
rect 32309 31263 32367 31269
rect 32309 31260 32321 31263
rect 31251 31232 32321 31260
rect 31251 31229 31263 31232
rect 31205 31223 31263 31229
rect 32309 31229 32321 31232
rect 32355 31260 32367 31263
rect 33962 31260 33968 31272
rect 32355 31232 33968 31260
rect 32355 31229 32367 31232
rect 32309 31223 32367 31229
rect 33962 31220 33968 31232
rect 34020 31220 34026 31272
rect 34790 31220 34796 31272
rect 34848 31260 34854 31272
rect 35161 31263 35219 31269
rect 35161 31260 35173 31263
rect 34848 31232 35173 31260
rect 34848 31220 34854 31232
rect 35161 31229 35173 31232
rect 35207 31229 35219 31263
rect 35161 31223 35219 31229
rect 15105 31195 15163 31201
rect 15105 31161 15117 31195
rect 15151 31192 15163 31195
rect 15151 31164 16574 31192
rect 15151 31161 15163 31164
rect 15105 31155 15163 31161
rect 16546 31124 16574 31164
rect 18874 31152 18880 31204
rect 18932 31192 18938 31204
rect 57422 31192 57428 31204
rect 18932 31164 57428 31192
rect 18932 31152 18938 31164
rect 57422 31152 57428 31164
rect 57480 31152 57486 31204
rect 16942 31124 16948 31136
rect 16546 31096 16948 31124
rect 16942 31084 16948 31096
rect 17000 31084 17006 31136
rect 22465 31127 22523 31133
rect 22465 31093 22477 31127
rect 22511 31124 22523 31127
rect 22554 31124 22560 31136
rect 22511 31096 22560 31124
rect 22511 31093 22523 31096
rect 22465 31087 22523 31093
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 24578 31124 24584 31136
rect 24539 31096 24584 31124
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 27154 31084 27160 31136
rect 27212 31124 27218 31136
rect 27433 31127 27491 31133
rect 27433 31124 27445 31127
rect 27212 31096 27445 31124
rect 27212 31084 27218 31096
rect 27433 31093 27445 31096
rect 27479 31124 27491 31127
rect 28350 31124 28356 31136
rect 27479 31096 28356 31124
rect 27479 31093 27491 31096
rect 27433 31087 27491 31093
rect 28350 31084 28356 31096
rect 28408 31084 28414 31136
rect 32950 31084 32956 31136
rect 33008 31124 33014 31136
rect 33505 31127 33563 31133
rect 33505 31124 33517 31127
rect 33008 31096 33517 31124
rect 33008 31084 33014 31096
rect 33505 31093 33517 31096
rect 33551 31093 33563 31127
rect 34330 31124 34336 31136
rect 34291 31096 34336 31124
rect 33505 31087 33563 31093
rect 34330 31084 34336 31096
rect 34388 31084 34394 31136
rect 35529 31127 35587 31133
rect 35529 31093 35541 31127
rect 35575 31124 35587 31127
rect 35986 31124 35992 31136
rect 35575 31096 35992 31124
rect 35575 31093 35587 31096
rect 35529 31087 35587 31093
rect 35986 31084 35992 31096
rect 36044 31084 36050 31136
rect 36909 31127 36967 31133
rect 36909 31093 36921 31127
rect 36955 31124 36967 31127
rect 37182 31124 37188 31136
rect 36955 31096 37188 31124
rect 36955 31093 36967 31096
rect 36909 31087 36967 31093
rect 37182 31084 37188 31096
rect 37240 31084 37246 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 15194 30880 15200 30932
rect 15252 30920 15258 30932
rect 15841 30923 15899 30929
rect 15841 30920 15853 30923
rect 15252 30892 15853 30920
rect 15252 30880 15258 30892
rect 15841 30889 15853 30892
rect 15887 30889 15899 30923
rect 15841 30883 15899 30889
rect 15930 30880 15936 30932
rect 15988 30920 15994 30932
rect 16025 30923 16083 30929
rect 16025 30920 16037 30923
rect 15988 30892 16037 30920
rect 15988 30880 15994 30892
rect 16025 30889 16037 30892
rect 16071 30889 16083 30923
rect 16025 30883 16083 30889
rect 20438 30880 20444 30932
rect 20496 30920 20502 30932
rect 20533 30923 20591 30929
rect 20533 30920 20545 30923
rect 20496 30892 20545 30920
rect 20496 30880 20502 30892
rect 20533 30889 20545 30892
rect 20579 30889 20591 30923
rect 25958 30920 25964 30932
rect 25919 30892 25964 30920
rect 20533 30883 20591 30889
rect 25958 30880 25964 30892
rect 26016 30880 26022 30932
rect 26878 30880 26884 30932
rect 26936 30920 26942 30932
rect 27433 30923 27491 30929
rect 27433 30920 27445 30923
rect 26936 30892 27445 30920
rect 26936 30880 26942 30892
rect 27433 30889 27445 30892
rect 27479 30889 27491 30923
rect 29178 30920 29184 30932
rect 27433 30883 27491 30889
rect 28966 30892 29184 30920
rect 22097 30855 22155 30861
rect 22097 30821 22109 30855
rect 22143 30852 22155 30855
rect 22278 30852 22284 30864
rect 22143 30824 22284 30852
rect 22143 30821 22155 30824
rect 22097 30815 22155 30821
rect 22278 30812 22284 30824
rect 22336 30812 22342 30864
rect 24581 30855 24639 30861
rect 24581 30821 24593 30855
rect 24627 30852 24639 30855
rect 24762 30852 24768 30864
rect 24627 30824 24768 30852
rect 24627 30821 24639 30824
rect 24581 30815 24639 30821
rect 24762 30812 24768 30824
rect 24820 30812 24826 30864
rect 16114 30784 16120 30796
rect 16075 30756 16120 30784
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 17954 30784 17960 30796
rect 17915 30756 17960 30784
rect 17954 30744 17960 30756
rect 18012 30744 18018 30796
rect 20254 30784 20260 30796
rect 18248 30756 20260 30784
rect 16209 30719 16267 30725
rect 16209 30685 16221 30719
rect 16255 30716 16267 30719
rect 16666 30716 16672 30728
rect 16255 30688 16672 30716
rect 16255 30685 16267 30688
rect 16209 30679 16267 30685
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 18248 30725 18276 30756
rect 20254 30744 20260 30756
rect 20312 30744 20318 30796
rect 21269 30787 21327 30793
rect 21269 30753 21281 30787
rect 21315 30784 21327 30787
rect 24302 30784 24308 30796
rect 21315 30756 24308 30784
rect 21315 30753 21327 30756
rect 21269 30747 21327 30753
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30685 18291 30719
rect 18874 30716 18880 30728
rect 18835 30688 18880 30716
rect 18233 30679 18291 30685
rect 18874 30676 18880 30688
rect 18932 30676 18938 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 20162 30716 20168 30728
rect 19751 30688 20168 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 20162 30676 20168 30688
rect 20220 30676 20226 30728
rect 20530 30657 20536 30660
rect 19889 30651 19947 30657
rect 19889 30617 19901 30651
rect 19935 30648 19947 30651
rect 20517 30651 20536 30657
rect 19935 30620 20392 30648
rect 19935 30617 19947 30620
rect 19889 30611 19947 30617
rect 19426 30540 19432 30592
rect 19484 30580 19490 30592
rect 20364 30589 20392 30620
rect 20517 30617 20529 30651
rect 20517 30611 20536 30617
rect 20530 30608 20536 30611
rect 20588 30608 20594 30660
rect 20714 30608 20720 30660
rect 20772 30648 20778 30660
rect 21284 30648 21312 30747
rect 24302 30744 24308 30756
rect 24360 30744 24366 30796
rect 25682 30784 25688 30796
rect 24872 30756 25688 30784
rect 21818 30716 21824 30728
rect 21779 30688 21824 30716
rect 21818 30676 21824 30688
rect 21876 30676 21882 30728
rect 22554 30716 22560 30728
rect 22515 30688 22560 30716
rect 22554 30676 22560 30688
rect 22612 30676 22618 30728
rect 22738 30716 22744 30728
rect 22699 30688 22744 30716
rect 22738 30676 22744 30688
rect 22796 30676 22802 30728
rect 23845 30719 23903 30725
rect 23845 30685 23857 30719
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 24029 30719 24087 30725
rect 24029 30685 24041 30719
rect 24075 30716 24087 30719
rect 24670 30716 24676 30728
rect 24075 30688 24676 30716
rect 24075 30685 24087 30688
rect 24029 30679 24087 30685
rect 20772 30620 21312 30648
rect 20772 30608 20778 30620
rect 22094 30608 22100 30660
rect 22152 30648 22158 30660
rect 22152 30620 22197 30648
rect 22152 30608 22158 30620
rect 19521 30583 19579 30589
rect 19521 30580 19533 30583
rect 19484 30552 19533 30580
rect 19484 30540 19490 30552
rect 19521 30549 19533 30552
rect 19567 30549 19579 30583
rect 19521 30543 19579 30549
rect 20349 30583 20407 30589
rect 20349 30549 20361 30583
rect 20395 30580 20407 30583
rect 20990 30580 20996 30592
rect 20395 30552 20996 30580
rect 20395 30549 20407 30552
rect 20349 30543 20407 30549
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 21913 30583 21971 30589
rect 21913 30549 21925 30583
rect 21959 30580 21971 30583
rect 22557 30583 22615 30589
rect 22557 30580 22569 30583
rect 21959 30552 22569 30580
rect 21959 30549 21971 30552
rect 21913 30543 21971 30549
rect 22557 30549 22569 30552
rect 22603 30549 22615 30583
rect 23860 30580 23888 30679
rect 24670 30676 24676 30688
rect 24728 30716 24734 30728
rect 24872 30725 24900 30756
rect 25682 30744 25688 30756
rect 25740 30784 25746 30796
rect 28966 30784 28994 30892
rect 29178 30880 29184 30892
rect 29236 30880 29242 30932
rect 31478 30920 31484 30932
rect 31439 30892 31484 30920
rect 31478 30880 31484 30892
rect 31536 30880 31542 30932
rect 34146 30920 34152 30932
rect 34107 30892 34152 30920
rect 34146 30880 34152 30892
rect 34204 30880 34210 30932
rect 34333 30923 34391 30929
rect 34333 30889 34345 30923
rect 34379 30920 34391 30923
rect 35342 30920 35348 30932
rect 34379 30892 35348 30920
rect 34379 30889 34391 30892
rect 34333 30883 34391 30889
rect 35342 30880 35348 30892
rect 35400 30880 35406 30932
rect 36173 30923 36231 30929
rect 36173 30889 36185 30923
rect 36219 30920 36231 30923
rect 36446 30920 36452 30932
rect 36219 30892 36452 30920
rect 36219 30889 36231 30892
rect 36173 30883 36231 30889
rect 36446 30880 36452 30892
rect 36504 30880 36510 30932
rect 32122 30852 32128 30864
rect 25740 30756 28994 30784
rect 30576 30824 32128 30852
rect 25740 30744 25746 30756
rect 24765 30719 24823 30725
rect 24765 30716 24777 30719
rect 24728 30688 24777 30716
rect 24728 30676 24734 30688
rect 24765 30685 24777 30688
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 25314 30676 25320 30728
rect 25372 30716 25378 30728
rect 25593 30719 25651 30725
rect 25593 30716 25605 30719
rect 25372 30688 25605 30716
rect 25372 30676 25378 30688
rect 25593 30685 25605 30688
rect 25639 30685 25651 30719
rect 26418 30716 26424 30728
rect 26379 30688 26424 30716
rect 25593 30679 25651 30685
rect 26418 30676 26424 30688
rect 26476 30676 26482 30728
rect 26970 30676 26976 30728
rect 27028 30716 27034 30728
rect 27433 30719 27491 30725
rect 27433 30716 27445 30719
rect 27028 30688 27445 30716
rect 27028 30676 27034 30688
rect 27433 30685 27445 30688
rect 27479 30685 27491 30719
rect 27433 30679 27491 30685
rect 27525 30719 27583 30725
rect 27525 30685 27537 30719
rect 27571 30685 27583 30719
rect 28258 30716 28264 30728
rect 28219 30688 28264 30716
rect 27525 30679 27583 30685
rect 23937 30651 23995 30657
rect 23937 30617 23949 30651
rect 23983 30648 23995 30651
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 23983 30620 24593 30648
rect 23983 30617 23995 30620
rect 23937 30611 23995 30617
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 25777 30651 25835 30657
rect 25777 30617 25789 30651
rect 25823 30648 25835 30651
rect 26510 30648 26516 30660
rect 25823 30620 26516 30648
rect 25823 30617 25835 30620
rect 25777 30611 25835 30617
rect 26510 30608 26516 30620
rect 26568 30608 26574 30660
rect 27540 30648 27568 30679
rect 28258 30676 28264 30688
rect 28316 30676 28322 30728
rect 28442 30716 28448 30728
rect 28403 30688 28448 30716
rect 28442 30676 28448 30688
rect 28500 30716 28506 30728
rect 28718 30716 28724 30728
rect 28500 30688 28724 30716
rect 28500 30676 28506 30688
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 30576 30725 30604 30824
rect 32122 30812 32128 30824
rect 32180 30812 32186 30864
rect 32490 30812 32496 30864
rect 32548 30852 32554 30864
rect 32769 30855 32827 30861
rect 32769 30852 32781 30855
rect 32548 30824 32781 30852
rect 32548 30812 32554 30824
rect 32769 30821 32781 30824
rect 32815 30821 32827 30855
rect 32769 30815 32827 30821
rect 30653 30787 30711 30793
rect 30653 30753 30665 30787
rect 30699 30784 30711 30787
rect 30834 30784 30840 30796
rect 30699 30756 30840 30784
rect 30699 30753 30711 30756
rect 30653 30747 30711 30753
rect 30834 30744 30840 30756
rect 30892 30744 30898 30796
rect 31018 30744 31024 30796
rect 31076 30784 31082 30796
rect 34238 30784 34244 30796
rect 31076 30756 31616 30784
rect 31076 30744 31082 30756
rect 30561 30719 30619 30725
rect 30561 30685 30573 30719
rect 30607 30685 30619 30719
rect 31386 30716 31392 30728
rect 31347 30688 31392 30716
rect 30561 30679 30619 30685
rect 31386 30676 31392 30688
rect 31444 30676 31450 30728
rect 31588 30725 31616 30756
rect 33888 30756 34244 30784
rect 31573 30719 31631 30725
rect 31573 30685 31585 30719
rect 31619 30685 31631 30719
rect 31573 30679 31631 30685
rect 32582 30676 32588 30728
rect 32640 30716 32646 30728
rect 32677 30719 32735 30725
rect 32677 30716 32689 30719
rect 32640 30688 32689 30716
rect 32640 30676 32646 30688
rect 32677 30685 32689 30688
rect 32723 30685 32735 30719
rect 32950 30716 32956 30728
rect 32911 30688 32956 30716
rect 32677 30679 32735 30685
rect 32692 30648 32720 30679
rect 32950 30676 32956 30688
rect 33008 30676 33014 30728
rect 33888 30725 33916 30756
rect 34238 30744 34244 30756
rect 34296 30784 34302 30796
rect 34977 30787 35035 30793
rect 34977 30784 34989 30787
rect 34296 30756 34989 30784
rect 34296 30744 34302 30756
rect 34977 30753 34989 30756
rect 35023 30753 35035 30787
rect 36078 30784 36084 30796
rect 34977 30747 35035 30753
rect 35912 30756 36084 30784
rect 33873 30719 33931 30725
rect 33873 30685 33885 30719
rect 33919 30685 33931 30719
rect 33873 30679 33931 30685
rect 33962 30676 33968 30728
rect 34020 30716 34026 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 34020 30688 34897 30716
rect 34020 30676 34026 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 35621 30719 35679 30725
rect 35621 30685 35633 30719
rect 35667 30685 35679 30719
rect 35621 30679 35679 30685
rect 33594 30648 33600 30660
rect 27540 30620 29040 30648
rect 32692 30620 33600 30648
rect 26326 30580 26332 30592
rect 23860 30552 26332 30580
rect 22557 30543 22615 30549
rect 26326 30540 26332 30552
rect 26384 30540 26390 30592
rect 26605 30583 26663 30589
rect 26605 30549 26617 30583
rect 26651 30580 26663 30583
rect 26878 30580 26884 30592
rect 26651 30552 26884 30580
rect 26651 30549 26663 30552
rect 26605 30543 26663 30549
rect 26878 30540 26884 30552
rect 26936 30540 26942 30592
rect 27062 30540 27068 30592
rect 27120 30580 27126 30592
rect 27430 30580 27436 30592
rect 27120 30552 27436 30580
rect 27120 30540 27126 30552
rect 27430 30540 27436 30552
rect 27488 30580 27494 30592
rect 27540 30580 27568 30620
rect 27798 30580 27804 30592
rect 27488 30552 27568 30580
rect 27759 30552 27804 30580
rect 27488 30540 27494 30552
rect 27798 30540 27804 30552
rect 27856 30540 27862 30592
rect 28353 30583 28411 30589
rect 28353 30549 28365 30583
rect 28399 30580 28411 30583
rect 28442 30580 28448 30592
rect 28399 30552 28448 30580
rect 28399 30549 28411 30552
rect 28353 30543 28411 30549
rect 28442 30540 28448 30552
rect 28500 30540 28506 30592
rect 29012 30589 29040 30620
rect 33594 30608 33600 30620
rect 33652 30648 33658 30660
rect 35084 30648 35112 30679
rect 33652 30620 35112 30648
rect 35636 30648 35664 30679
rect 35710 30676 35716 30728
rect 35768 30716 35774 30728
rect 35912 30725 35940 30756
rect 36078 30744 36084 30756
rect 36136 30744 36142 30796
rect 37274 30784 37280 30796
rect 37235 30756 37280 30784
rect 37274 30744 37280 30756
rect 37332 30744 37338 30796
rect 38013 30787 38071 30793
rect 38013 30753 38025 30787
rect 38059 30784 38071 30787
rect 41322 30784 41328 30796
rect 38059 30756 41328 30784
rect 38059 30753 38071 30756
rect 38013 30747 38071 30753
rect 41322 30744 41328 30756
rect 41380 30744 41386 30796
rect 35897 30719 35955 30725
rect 35768 30688 35813 30716
rect 35768 30676 35774 30688
rect 35897 30685 35909 30719
rect 35943 30685 35955 30719
rect 35897 30679 35955 30685
rect 35986 30676 35992 30728
rect 36044 30716 36050 30728
rect 37182 30716 37188 30728
rect 36044 30688 36089 30716
rect 37143 30688 37188 30716
rect 36044 30676 36050 30688
rect 37182 30676 37188 30688
rect 37240 30676 37246 30728
rect 35636 30620 35940 30648
rect 33652 30608 33658 30620
rect 35912 30592 35940 30620
rect 28997 30583 29055 30589
rect 28997 30549 29009 30583
rect 29043 30580 29055 30583
rect 29270 30580 29276 30592
rect 29043 30552 29276 30580
rect 29043 30549 29055 30552
rect 28997 30543 29055 30549
rect 29270 30540 29276 30552
rect 29328 30580 29334 30592
rect 29546 30580 29552 30592
rect 29328 30552 29552 30580
rect 29328 30540 29334 30552
rect 29546 30540 29552 30552
rect 29604 30540 29610 30592
rect 30926 30580 30932 30592
rect 30887 30552 30932 30580
rect 30926 30540 30932 30552
rect 30984 30540 30990 30592
rect 35894 30540 35900 30592
rect 35952 30540 35958 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 17954 30376 17960 30388
rect 17915 30348 17960 30376
rect 17954 30336 17960 30348
rect 18012 30336 18018 30388
rect 20438 30376 20444 30388
rect 20180 30348 20444 30376
rect 20180 30317 20208 30348
rect 20438 30336 20444 30348
rect 20496 30336 20502 30388
rect 23845 30379 23903 30385
rect 23845 30345 23857 30379
rect 23891 30376 23903 30379
rect 26234 30376 26240 30388
rect 23891 30348 26240 30376
rect 23891 30345 23903 30348
rect 23845 30339 23903 30345
rect 26234 30336 26240 30348
rect 26292 30336 26298 30388
rect 26418 30336 26424 30388
rect 26476 30376 26482 30388
rect 26605 30379 26663 30385
rect 26605 30376 26617 30379
rect 26476 30348 26617 30376
rect 26476 30336 26482 30348
rect 26605 30345 26617 30348
rect 26651 30345 26663 30379
rect 26605 30339 26663 30345
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 27617 30379 27675 30385
rect 27617 30376 27629 30379
rect 27580 30348 27629 30376
rect 27580 30336 27586 30348
rect 27617 30345 27629 30348
rect 27663 30345 27675 30379
rect 27617 30339 27675 30345
rect 28626 30336 28632 30388
rect 28684 30336 28690 30388
rect 34790 30376 34796 30388
rect 33796 30348 34796 30376
rect 20165 30311 20223 30317
rect 20165 30277 20177 30311
rect 20211 30277 20223 30311
rect 20165 30271 20223 30277
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20714 30308 20720 30320
rect 20395 30280 20720 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 18046 30200 18052 30252
rect 18104 30240 18110 30252
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 18104 30212 18153 30240
rect 18104 30200 18110 30212
rect 18141 30209 18153 30212
rect 18187 30209 18199 30243
rect 18141 30203 18199 30209
rect 18417 30243 18475 30249
rect 18417 30209 18429 30243
rect 18463 30240 18475 30243
rect 18506 30240 18512 30252
rect 18463 30212 18512 30240
rect 18463 30209 18475 30212
rect 18417 30203 18475 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 18601 30243 18659 30249
rect 18601 30209 18613 30243
rect 18647 30240 18659 30243
rect 19426 30240 19432 30252
rect 18647 30212 19432 30240
rect 18647 30209 18659 30212
rect 18601 30203 18659 30209
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20364 30240 20392 30271
rect 20714 30268 20720 30280
rect 20772 30268 20778 30320
rect 27062 30308 27068 30320
rect 25976 30280 27068 30308
rect 19751 30212 20392 30240
rect 20441 30243 20499 30249
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 20441 30209 20453 30243
rect 20487 30240 20499 30243
rect 20530 30240 20536 30252
rect 20487 30212 20536 30240
rect 20487 30209 20499 30212
rect 20441 30203 20499 30209
rect 20530 30200 20536 30212
rect 20588 30200 20594 30252
rect 20898 30240 20904 30252
rect 20859 30212 20904 30240
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 20990 30200 20996 30252
rect 21048 30240 21054 30252
rect 21048 30212 21093 30240
rect 21048 30200 21054 30212
rect 22554 30200 22560 30252
rect 22612 30240 22618 30252
rect 22741 30243 22799 30249
rect 22741 30240 22753 30243
rect 22612 30212 22753 30240
rect 22612 30200 22618 30212
rect 22741 30209 22753 30212
rect 22787 30209 22799 30243
rect 22741 30203 22799 30209
rect 23934 30200 23940 30252
rect 23992 30240 23998 30252
rect 24029 30243 24087 30249
rect 24029 30240 24041 30243
rect 23992 30212 24041 30240
rect 23992 30200 23998 30212
rect 24029 30209 24041 30212
rect 24075 30240 24087 30243
rect 24210 30240 24216 30252
rect 24075 30212 24216 30240
rect 24075 30209 24087 30212
rect 24029 30203 24087 30209
rect 24210 30200 24216 30212
rect 24268 30200 24274 30252
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 24673 30243 24731 30249
rect 24673 30240 24685 30243
rect 24636 30212 24685 30240
rect 24636 30200 24642 30212
rect 24673 30209 24685 30212
rect 24719 30209 24731 30243
rect 24673 30203 24731 30209
rect 24762 30200 24768 30252
rect 24820 30240 24826 30252
rect 24857 30243 24915 30249
rect 24857 30240 24869 30243
rect 24820 30212 24869 30240
rect 24820 30200 24826 30212
rect 24857 30209 24869 30212
rect 24903 30209 24915 30243
rect 24857 30203 24915 30209
rect 20806 30132 20812 30184
rect 20864 30172 20870 30184
rect 21177 30175 21235 30181
rect 21177 30172 21189 30175
rect 20864 30144 21189 30172
rect 20864 30132 20870 30144
rect 21177 30141 21189 30144
rect 21223 30141 21235 30175
rect 22646 30172 22652 30184
rect 22607 30144 22652 30172
rect 21177 30135 21235 30141
rect 22646 30132 22652 30144
rect 22704 30132 22710 30184
rect 25976 30181 26004 30280
rect 27062 30268 27068 30280
rect 27120 30268 27126 30320
rect 26326 30200 26332 30252
rect 26384 30240 26390 30252
rect 26602 30240 26608 30252
rect 26384 30212 26608 30240
rect 26384 30200 26390 30212
rect 26602 30200 26608 30212
rect 26660 30240 26666 30252
rect 27525 30243 27583 30249
rect 27525 30240 27537 30243
rect 26660 30212 27537 30240
rect 26660 30200 26666 30212
rect 27525 30209 27537 30212
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 25961 30175 26019 30181
rect 25961 30141 25973 30175
rect 26007 30141 26019 30175
rect 25961 30135 26019 30141
rect 26145 30175 26203 30181
rect 26145 30141 26157 30175
rect 26191 30172 26203 30175
rect 26191 30144 27200 30172
rect 26191 30141 26203 30144
rect 26145 30135 26203 30141
rect 20162 30104 20168 30116
rect 20123 30076 20168 30104
rect 20162 30064 20168 30076
rect 20220 30064 20226 30116
rect 23750 30064 23756 30116
rect 23808 30104 23814 30116
rect 27172 30113 27200 30144
rect 27614 30132 27620 30184
rect 27672 30172 27678 30184
rect 27709 30175 27767 30181
rect 27709 30172 27721 30175
rect 27672 30144 27721 30172
rect 27672 30132 27678 30144
rect 27709 30141 27721 30144
rect 27755 30141 27767 30175
rect 28368 30172 28396 30203
rect 28442 30200 28448 30252
rect 28500 30240 28506 30252
rect 28644 30249 28672 30336
rect 29362 30308 29368 30320
rect 29323 30280 29368 30308
rect 29362 30268 29368 30280
rect 29420 30268 29426 30320
rect 33796 30308 33824 30348
rect 34790 30336 34796 30348
rect 34848 30376 34854 30388
rect 34848 30348 36308 30376
rect 34848 30336 34854 30348
rect 33962 30308 33968 30320
rect 33244 30280 33824 30308
rect 33923 30280 33968 30308
rect 28629 30243 28687 30249
rect 28500 30212 28545 30240
rect 28500 30200 28506 30212
rect 28629 30209 28641 30243
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 28718 30200 28724 30252
rect 28776 30240 28782 30252
rect 28776 30212 28821 30240
rect 28776 30200 28782 30212
rect 28994 30172 29000 30184
rect 28368 30144 29000 30172
rect 27709 30135 27767 30141
rect 28994 30132 29000 30144
rect 29052 30172 29058 30184
rect 29380 30172 29408 30268
rect 31570 30240 31576 30252
rect 31531 30212 31576 30240
rect 31570 30200 31576 30212
rect 31628 30200 31634 30252
rect 32766 30240 32772 30252
rect 32727 30212 32772 30240
rect 32766 30200 32772 30212
rect 32824 30200 32830 30252
rect 29052 30144 29408 30172
rect 31665 30175 31723 30181
rect 29052 30132 29058 30144
rect 31665 30141 31677 30175
rect 31711 30172 31723 30175
rect 32122 30172 32128 30184
rect 31711 30144 32128 30172
rect 31711 30141 31723 30144
rect 31665 30135 31723 30141
rect 32122 30132 32128 30144
rect 32180 30132 32186 30184
rect 33244 30181 33272 30280
rect 33962 30268 33968 30280
rect 34020 30268 34026 30320
rect 34146 30308 34152 30320
rect 34204 30317 34210 30320
rect 34204 30311 34239 30317
rect 34091 30280 34152 30308
rect 34146 30268 34152 30280
rect 34227 30308 34239 30311
rect 34885 30311 34943 30317
rect 34885 30308 34897 30311
rect 34227 30280 34897 30308
rect 34227 30277 34239 30280
rect 34204 30271 34239 30277
rect 34885 30277 34897 30280
rect 34931 30277 34943 30311
rect 34885 30271 34943 30277
rect 34204 30268 34210 30271
rect 35434 30268 35440 30320
rect 35492 30308 35498 30320
rect 35713 30311 35771 30317
rect 35713 30308 35725 30311
rect 35492 30280 35725 30308
rect 35492 30268 35498 30280
rect 35713 30277 35725 30280
rect 35759 30277 35771 30311
rect 35713 30271 35771 30277
rect 35986 30268 35992 30320
rect 36044 30308 36050 30320
rect 36044 30280 36216 30308
rect 36044 30268 36050 30280
rect 34054 30200 34060 30252
rect 34112 30240 34118 30252
rect 34793 30243 34851 30249
rect 34793 30240 34805 30243
rect 34112 30212 34805 30240
rect 34112 30200 34118 30212
rect 34793 30209 34805 30212
rect 34839 30209 34851 30243
rect 34793 30203 34851 30209
rect 34977 30243 35035 30249
rect 34977 30209 34989 30243
rect 35023 30209 35035 30243
rect 35894 30240 35900 30252
rect 35807 30212 35900 30240
rect 34977 30203 35035 30209
rect 33229 30175 33287 30181
rect 33229 30141 33241 30175
rect 33275 30141 33287 30175
rect 33229 30135 33287 30141
rect 34330 30132 34336 30184
rect 34388 30172 34394 30184
rect 34992 30172 35020 30203
rect 35894 30200 35900 30212
rect 35952 30200 35958 30252
rect 36078 30240 36084 30252
rect 36039 30212 36084 30240
rect 36078 30200 36084 30212
rect 36136 30200 36142 30252
rect 36188 30249 36216 30280
rect 36173 30243 36231 30249
rect 36173 30209 36185 30243
rect 36219 30209 36231 30243
rect 36173 30203 36231 30209
rect 34388 30144 35020 30172
rect 34388 30132 34394 30144
rect 27157 30107 27215 30113
rect 23808 30076 25452 30104
rect 23808 30064 23814 30076
rect 21082 29996 21088 30048
rect 21140 30036 21146 30048
rect 21140 30008 21185 30036
rect 21140 29996 21146 30008
rect 21726 29996 21732 30048
rect 21784 30036 21790 30048
rect 22465 30039 22523 30045
rect 22465 30036 22477 30039
rect 21784 30008 22477 30036
rect 21784 29996 21790 30008
rect 22465 30005 22477 30008
rect 22511 30005 22523 30039
rect 22465 29999 22523 30005
rect 25041 30039 25099 30045
rect 25041 30005 25053 30039
rect 25087 30036 25099 30039
rect 25314 30036 25320 30048
rect 25087 30008 25320 30036
rect 25087 30005 25099 30008
rect 25041 29999 25099 30005
rect 25314 29996 25320 30008
rect 25372 29996 25378 30048
rect 25424 30036 25452 30076
rect 27157 30073 27169 30107
rect 27203 30073 27215 30107
rect 31205 30107 31263 30113
rect 31205 30104 31217 30107
rect 27157 30067 27215 30073
rect 27264 30076 31217 30104
rect 27264 30036 27292 30076
rect 31205 30073 31217 30076
rect 31251 30073 31263 30107
rect 35912 30104 35940 30200
rect 36280 30172 36308 30348
rect 36725 30311 36783 30317
rect 36725 30277 36737 30311
rect 36771 30308 36783 30311
rect 37274 30308 37280 30320
rect 36771 30280 37280 30308
rect 36771 30277 36783 30280
rect 36725 30271 36783 30277
rect 37274 30268 37280 30280
rect 37332 30268 37338 30320
rect 36630 30240 36636 30252
rect 36591 30212 36636 30240
rect 36630 30200 36636 30212
rect 36688 30200 36694 30252
rect 36817 30243 36875 30249
rect 36817 30209 36829 30243
rect 36863 30209 36875 30243
rect 36817 30203 36875 30209
rect 36832 30172 36860 30203
rect 36280 30144 36860 30172
rect 31205 30067 31263 30073
rect 34348 30076 35940 30104
rect 28902 30036 28908 30048
rect 25424 30008 27292 30036
rect 28863 30008 28908 30036
rect 28902 29996 28908 30008
rect 28960 29996 28966 30048
rect 32490 29996 32496 30048
rect 32548 30036 32554 30048
rect 32861 30039 32919 30045
rect 32861 30036 32873 30039
rect 32548 30008 32873 30036
rect 32548 29996 32554 30008
rect 32861 30005 32873 30008
rect 32907 30005 32919 30039
rect 32861 29999 32919 30005
rect 33594 29996 33600 30048
rect 33652 30036 33658 30048
rect 34348 30045 34376 30076
rect 36078 30064 36084 30116
rect 36136 30104 36142 30116
rect 36630 30104 36636 30116
rect 36136 30076 36636 30104
rect 36136 30064 36142 30076
rect 36630 30064 36636 30076
rect 36688 30064 36694 30116
rect 34149 30039 34207 30045
rect 34149 30036 34161 30039
rect 33652 30008 34161 30036
rect 33652 29996 33658 30008
rect 34149 30005 34161 30008
rect 34195 30005 34207 30039
rect 34149 29999 34207 30005
rect 34333 30039 34391 30045
rect 34333 30005 34345 30039
rect 34379 30005 34391 30039
rect 34333 29999 34391 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 20809 29835 20867 29841
rect 20809 29801 20821 29835
rect 20855 29832 20867 29835
rect 20990 29832 20996 29844
rect 20855 29804 20996 29832
rect 20855 29801 20867 29804
rect 20809 29795 20867 29801
rect 20990 29792 20996 29804
rect 21048 29792 21054 29844
rect 22094 29792 22100 29844
rect 22152 29832 22158 29844
rect 22557 29835 22615 29841
rect 22557 29832 22569 29835
rect 22152 29804 22569 29832
rect 22152 29792 22158 29804
rect 22557 29801 22569 29804
rect 22603 29801 22615 29835
rect 22557 29795 22615 29801
rect 27522 29792 27528 29844
rect 27580 29832 27586 29844
rect 27617 29835 27675 29841
rect 27617 29832 27629 29835
rect 27580 29804 27629 29832
rect 27580 29792 27586 29804
rect 27617 29801 27629 29804
rect 27663 29801 27675 29835
rect 27617 29795 27675 29801
rect 28629 29835 28687 29841
rect 28629 29801 28641 29835
rect 28675 29832 28687 29835
rect 29086 29832 29092 29844
rect 28675 29804 29092 29832
rect 28675 29801 28687 29804
rect 28629 29795 28687 29801
rect 29086 29792 29092 29804
rect 29144 29792 29150 29844
rect 31294 29792 31300 29844
rect 31352 29832 31358 29844
rect 33686 29832 33692 29844
rect 31352 29804 33692 29832
rect 31352 29792 31358 29804
rect 33686 29792 33692 29804
rect 33744 29792 33750 29844
rect 18506 29724 18512 29776
rect 18564 29764 18570 29776
rect 19705 29767 19763 29773
rect 19705 29764 19717 29767
rect 18564 29736 19717 29764
rect 18564 29724 18570 29736
rect 19705 29733 19717 29736
rect 19751 29733 19763 29767
rect 21082 29764 21088 29776
rect 19705 29727 19763 29733
rect 20088 29736 21088 29764
rect 20088 29640 20116 29736
rect 21082 29724 21088 29736
rect 21140 29724 21146 29776
rect 24762 29724 24768 29776
rect 24820 29764 24826 29776
rect 26145 29767 26203 29773
rect 24820 29736 24900 29764
rect 24820 29724 24826 29736
rect 20717 29699 20775 29705
rect 20717 29665 20729 29699
rect 20763 29696 20775 29699
rect 20898 29696 20904 29708
rect 20763 29668 20904 29696
rect 20763 29665 20775 29668
rect 20717 29659 20775 29665
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 21818 29696 21824 29708
rect 21779 29668 21824 29696
rect 21818 29656 21824 29668
rect 21876 29656 21882 29708
rect 24872 29705 24900 29736
rect 26145 29733 26157 29767
rect 26191 29764 26203 29767
rect 32953 29767 33011 29773
rect 26191 29736 26648 29764
rect 26191 29733 26203 29736
rect 26145 29727 26203 29733
rect 24857 29699 24915 29705
rect 24857 29665 24869 29699
rect 24903 29665 24915 29699
rect 24857 29659 24915 29665
rect 25038 29656 25044 29708
rect 25096 29696 25102 29708
rect 26620 29705 26648 29736
rect 32953 29733 32965 29767
rect 32999 29764 33011 29767
rect 34054 29764 34060 29776
rect 32999 29736 34060 29764
rect 32999 29733 33011 29736
rect 32953 29727 33011 29733
rect 34054 29724 34060 29736
rect 34112 29724 34118 29776
rect 25133 29699 25191 29705
rect 25133 29696 25145 29699
rect 25096 29668 25145 29696
rect 25096 29656 25102 29668
rect 25133 29665 25145 29668
rect 25179 29665 25191 29699
rect 25133 29659 25191 29665
rect 26605 29699 26663 29705
rect 26605 29665 26617 29699
rect 26651 29665 26663 29699
rect 28994 29696 29000 29708
rect 26605 29659 26663 29665
rect 28552 29668 29000 29696
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19484 29600 19625 29628
rect 19484 29588 19490 29600
rect 19613 29597 19625 29600
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29597 19855 29631
rect 19797 29591 19855 29597
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 20070 29628 20076 29640
rect 19935 29600 20076 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 19812 29560 19840 29591
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20806 29628 20812 29640
rect 20767 29600 20812 29628
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 21726 29628 21732 29640
rect 21687 29600 21732 29628
rect 21726 29588 21732 29600
rect 21784 29588 21790 29640
rect 22373 29631 22431 29637
rect 22373 29597 22385 29631
rect 22419 29628 22431 29631
rect 22462 29628 22468 29640
rect 22419 29600 22468 29628
rect 22419 29597 22431 29600
rect 22373 29591 22431 29597
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22557 29631 22615 29637
rect 22557 29597 22569 29631
rect 22603 29628 22615 29631
rect 22646 29628 22652 29640
rect 22603 29600 22652 29628
rect 22603 29597 22615 29600
rect 22557 29591 22615 29597
rect 22646 29588 22652 29600
rect 22704 29588 22710 29640
rect 24578 29588 24584 29640
rect 24636 29628 24642 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24636 29600 24777 29628
rect 24636 29588 24642 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 25958 29628 25964 29640
rect 25919 29600 25964 29628
rect 24765 29591 24823 29597
rect 25958 29588 25964 29600
rect 26016 29588 26022 29640
rect 26878 29628 26884 29640
rect 26839 29600 26884 29628
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 28552 29637 28580 29668
rect 28994 29656 29000 29668
rect 29052 29656 29058 29708
rect 29270 29656 29276 29708
rect 29328 29696 29334 29708
rect 33410 29696 33416 29708
rect 29328 29668 31754 29696
rect 29328 29656 29334 29668
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28902 29588 28908 29640
rect 28960 29628 28966 29640
rect 29638 29628 29644 29640
rect 28960 29600 29644 29628
rect 28960 29588 28966 29600
rect 29638 29588 29644 29600
rect 29696 29628 29702 29640
rect 29825 29631 29883 29637
rect 29825 29628 29837 29631
rect 29696 29600 29837 29628
rect 29696 29588 29702 29600
rect 29825 29597 29837 29600
rect 29871 29597 29883 29631
rect 29825 29591 29883 29597
rect 30098 29588 30104 29640
rect 30156 29588 30162 29640
rect 20622 29560 20628 29572
rect 19812 29532 20628 29560
rect 20622 29520 20628 29532
rect 20680 29520 20686 29572
rect 30834 29560 30840 29572
rect 30795 29532 30840 29560
rect 30834 29520 30840 29532
rect 30892 29520 30898 29572
rect 31570 29560 31576 29572
rect 30944 29532 31576 29560
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19392 29464 19441 29492
rect 19392 29452 19398 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20441 29495 20499 29501
rect 20441 29492 20453 29495
rect 20036 29464 20453 29492
rect 20036 29452 20042 29464
rect 20441 29461 20453 29464
rect 20487 29461 20499 29495
rect 20441 29455 20499 29461
rect 20806 29452 20812 29504
rect 20864 29492 20870 29504
rect 21361 29495 21419 29501
rect 21361 29492 21373 29495
rect 20864 29464 21373 29492
rect 20864 29452 20870 29464
rect 21361 29461 21373 29464
rect 21407 29461 21419 29495
rect 23842 29492 23848 29504
rect 23803 29464 23848 29492
rect 21361 29455 21419 29461
rect 23842 29452 23848 29464
rect 23900 29452 23906 29504
rect 24118 29452 24124 29504
rect 24176 29492 24182 29504
rect 30944 29492 30972 29532
rect 31570 29520 31576 29532
rect 31628 29520 31634 29572
rect 31726 29560 31754 29668
rect 32692 29668 33416 29696
rect 32692 29637 32720 29668
rect 33410 29656 33416 29668
rect 33468 29656 33474 29708
rect 32217 29631 32275 29637
rect 32217 29597 32229 29631
rect 32263 29628 32275 29631
rect 32677 29631 32735 29637
rect 32677 29628 32689 29631
rect 32263 29600 32689 29628
rect 32263 29597 32275 29600
rect 32217 29591 32275 29597
rect 32677 29597 32689 29600
rect 32723 29597 32735 29631
rect 32677 29591 32735 29597
rect 32953 29631 33011 29637
rect 32953 29597 32965 29631
rect 32999 29628 33011 29631
rect 33042 29628 33048 29640
rect 32999 29600 33048 29628
rect 32999 29597 33011 29600
rect 32953 29591 33011 29597
rect 33042 29588 33048 29600
rect 33100 29588 33106 29640
rect 33505 29631 33563 29637
rect 33505 29597 33517 29631
rect 33551 29597 33563 29631
rect 33505 29591 33563 29597
rect 33520 29560 33548 29591
rect 34149 29563 34207 29569
rect 34149 29560 34161 29563
rect 31726 29532 34161 29560
rect 34149 29529 34161 29532
rect 34195 29529 34207 29563
rect 34149 29523 34207 29529
rect 31294 29492 31300 29504
rect 24176 29464 30972 29492
rect 31255 29464 31300 29492
rect 24176 29452 24182 29464
rect 31294 29452 31300 29464
rect 31352 29452 31358 29504
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 32769 29495 32827 29501
rect 32769 29492 32781 29495
rect 32456 29464 32781 29492
rect 32456 29452 32462 29464
rect 32769 29461 32781 29464
rect 32815 29492 32827 29495
rect 33505 29495 33563 29501
rect 33505 29492 33517 29495
rect 32815 29464 33517 29492
rect 32815 29461 32827 29464
rect 32769 29455 32827 29461
rect 33505 29461 33517 29464
rect 33551 29461 33563 29495
rect 33505 29455 33563 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 2409 29291 2467 29297
rect 2409 29257 2421 29291
rect 2455 29288 2467 29291
rect 24118 29288 24124 29300
rect 2455 29260 24124 29288
rect 2455 29257 2467 29260
rect 2409 29251 2467 29257
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29152 1915 29155
rect 2424 29152 2452 29251
rect 24118 29248 24124 29260
rect 24176 29248 24182 29300
rect 25958 29248 25964 29300
rect 26016 29288 26022 29300
rect 27157 29291 27215 29297
rect 27157 29288 27169 29291
rect 26016 29260 27169 29288
rect 26016 29248 26022 29260
rect 27157 29257 27169 29260
rect 27203 29257 27215 29291
rect 27157 29251 27215 29257
rect 28445 29291 28503 29297
rect 28445 29257 28457 29291
rect 28491 29288 28503 29291
rect 28994 29288 29000 29300
rect 28491 29260 29000 29288
rect 28491 29257 28503 29260
rect 28445 29251 28503 29257
rect 28994 29248 29000 29260
rect 29052 29248 29058 29300
rect 30653 29291 30711 29297
rect 30653 29288 30665 29291
rect 30208 29260 30665 29288
rect 16942 29220 16948 29232
rect 16903 29192 16948 29220
rect 16942 29180 16948 29192
rect 17000 29180 17006 29232
rect 18506 29220 18512 29232
rect 18156 29192 18512 29220
rect 1903 29124 2452 29152
rect 1903 29121 1915 29124
rect 1857 29115 1915 29121
rect 17405 29087 17463 29093
rect 17405 29053 17417 29087
rect 17451 29084 17463 29087
rect 18046 29084 18052 29096
rect 17451 29056 18052 29084
rect 17451 29053 17463 29056
rect 17405 29047 17463 29053
rect 18046 29044 18052 29056
rect 18104 29044 18110 29096
rect 18156 29093 18184 29192
rect 18506 29180 18512 29192
rect 18564 29180 18570 29232
rect 20898 29220 20904 29232
rect 19168 29192 20024 29220
rect 20859 29192 20904 29220
rect 19168 29161 19196 29192
rect 19996 29164 20024 29192
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 25130 29180 25136 29232
rect 25188 29180 25194 29232
rect 30208 29229 30236 29260
rect 30653 29257 30665 29260
rect 30699 29257 30711 29291
rect 30653 29251 30711 29257
rect 31757 29291 31815 29297
rect 31757 29257 31769 29291
rect 31803 29288 31815 29291
rect 33134 29288 33140 29300
rect 31803 29260 33140 29288
rect 31803 29257 31815 29260
rect 31757 29251 31815 29257
rect 33134 29248 33140 29260
rect 33192 29248 33198 29300
rect 30193 29223 30251 29229
rect 30193 29189 30205 29223
rect 30239 29189 30251 29223
rect 30193 29183 30251 29189
rect 30745 29223 30803 29229
rect 30745 29189 30757 29223
rect 30791 29220 30803 29223
rect 30834 29220 30840 29232
rect 30791 29192 30840 29220
rect 30791 29189 30803 29192
rect 30745 29183 30803 29189
rect 30834 29180 30840 29192
rect 30892 29180 30898 29232
rect 30926 29180 30932 29232
rect 30984 29220 30990 29232
rect 31389 29223 31447 29229
rect 30984 29192 31029 29220
rect 30984 29180 30990 29192
rect 31389 29189 31401 29223
rect 31435 29189 31447 29223
rect 31389 29183 31447 29189
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29121 19211 29155
rect 19153 29115 19211 29121
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29152 19395 29155
rect 19978 29152 19984 29164
rect 19383 29124 19748 29152
rect 19939 29124 19984 29152
rect 19383 29121 19395 29124
rect 19337 29115 19395 29121
rect 18141 29087 18199 29093
rect 18141 29053 18153 29087
rect 18187 29053 18199 29087
rect 18248 29084 18276 29115
rect 19426 29084 19432 29096
rect 18248 29056 19432 29084
rect 18141 29047 18199 29053
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 19720 29084 19748 29124
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20070 29112 20076 29164
rect 20128 29152 20134 29164
rect 20625 29155 20683 29161
rect 20128 29124 20173 29152
rect 20128 29112 20134 29124
rect 20625 29121 20637 29155
rect 20671 29152 20683 29155
rect 20806 29152 20812 29164
rect 20671 29124 20812 29152
rect 20671 29121 20683 29124
rect 20625 29115 20683 29121
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 21358 29112 21364 29164
rect 21416 29152 21422 29164
rect 23569 29155 23627 29161
rect 23569 29152 23581 29155
rect 21416 29124 23581 29152
rect 21416 29112 21422 29124
rect 23569 29121 23581 29124
rect 23615 29121 23627 29155
rect 23750 29152 23756 29164
rect 23711 29124 23756 29152
rect 23569 29115 23627 29121
rect 20088 29084 20116 29112
rect 19720 29056 20116 29084
rect 20717 29087 20775 29093
rect 20717 29053 20729 29087
rect 20763 29084 20775 29087
rect 20990 29084 20996 29096
rect 20763 29056 20996 29084
rect 20763 29053 20775 29056
rect 20717 29047 20775 29053
rect 20990 29044 20996 29056
rect 21048 29044 21054 29096
rect 1670 29016 1676 29028
rect 1631 28988 1676 29016
rect 1670 28976 1676 28988
rect 1728 28976 1734 29028
rect 17313 29019 17371 29025
rect 17313 28985 17325 29019
rect 17359 29016 17371 29019
rect 18064 29016 18092 29044
rect 18874 29016 18880 29028
rect 17359 28988 17908 29016
rect 18064 28988 18880 29016
rect 17359 28985 17371 28988
rect 17313 28979 17371 28985
rect 17880 28960 17908 28988
rect 18874 28976 18880 28988
rect 18932 28976 18938 29028
rect 19245 29019 19303 29025
rect 19245 28985 19257 29019
rect 19291 29016 19303 29019
rect 19610 29016 19616 29028
rect 19291 28988 19616 29016
rect 19291 28985 19303 28988
rect 19245 28979 19303 28985
rect 19610 28976 19616 28988
rect 19668 28976 19674 29028
rect 19797 29019 19855 29025
rect 19797 28985 19809 29019
rect 19843 29016 19855 29019
rect 20254 29016 20260 29028
rect 19843 28988 20260 29016
rect 19843 28985 19855 28988
rect 19797 28979 19855 28985
rect 17862 28948 17868 28960
rect 17823 28920 17868 28948
rect 17862 28908 17868 28920
rect 17920 28908 17926 28960
rect 19426 28908 19432 28960
rect 19484 28948 19490 28960
rect 19812 28948 19840 28979
rect 20254 28976 20260 28988
rect 20312 28976 20318 29028
rect 20622 29016 20628 29028
rect 20583 28988 20628 29016
rect 20622 28976 20628 28988
rect 20680 28976 20686 29028
rect 23584 29016 23612 29115
rect 23750 29112 23756 29124
rect 23808 29152 23814 29164
rect 24923 29155 24981 29161
rect 24923 29152 24935 29155
rect 23808 29124 24935 29152
rect 23808 29112 23814 29124
rect 24923 29121 24935 29124
rect 24969 29121 24981 29155
rect 24923 29115 24981 29121
rect 25019 29155 25077 29161
rect 25019 29121 25031 29155
rect 25065 29152 25077 29155
rect 25148 29152 25176 29180
rect 25065 29124 25176 29152
rect 25225 29155 25283 29161
rect 25065 29121 25077 29124
rect 25019 29115 25077 29121
rect 25225 29121 25237 29155
rect 25271 29152 25283 29155
rect 25314 29152 25320 29164
rect 25271 29124 25320 29152
rect 25271 29121 25283 29124
rect 25225 29115 25283 29121
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29152 26111 29155
rect 26605 29155 26663 29161
rect 26605 29152 26617 29155
rect 26099 29124 26617 29152
rect 26099 29121 26111 29124
rect 26053 29115 26111 29121
rect 26605 29121 26617 29124
rect 26651 29152 26663 29155
rect 27341 29155 27399 29161
rect 27341 29152 27353 29155
rect 26651 29124 27353 29152
rect 26651 29121 26663 29124
rect 26605 29115 26663 29121
rect 27341 29121 27353 29124
rect 27387 29152 27399 29155
rect 27430 29152 27436 29164
rect 27387 29124 27436 29152
rect 27387 29121 27399 29124
rect 27341 29115 27399 29121
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 28261 29155 28319 29161
rect 28261 29152 28273 29155
rect 27724 29124 28273 29152
rect 24302 29084 24308 29096
rect 24215 29056 24308 29084
rect 24302 29044 24308 29056
rect 24360 29084 24366 29096
rect 25133 29087 25191 29093
rect 25133 29084 25145 29087
rect 24360 29056 25145 29084
rect 24360 29044 24366 29056
rect 25133 29053 25145 29056
rect 25179 29084 25191 29087
rect 26970 29084 26976 29096
rect 25179 29056 26976 29084
rect 25179 29053 25191 29056
rect 25133 29047 25191 29053
rect 26970 29044 26976 29056
rect 27028 29044 27034 29096
rect 27522 29084 27528 29096
rect 27483 29056 27528 29084
rect 27522 29044 27528 29056
rect 27580 29044 27586 29096
rect 27614 29044 27620 29096
rect 27672 29084 27678 29096
rect 27724 29084 27752 29124
rect 28261 29121 28273 29124
rect 28307 29121 28319 29155
rect 28534 29152 28540 29164
rect 28495 29124 28540 29152
rect 28261 29115 28319 29121
rect 28534 29112 28540 29124
rect 28592 29112 28598 29164
rect 29638 29152 29644 29164
rect 29599 29124 29644 29152
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29152 29883 29155
rect 30098 29152 30104 29164
rect 29871 29124 30104 29152
rect 29871 29121 29883 29124
rect 29825 29115 29883 29121
rect 30098 29112 30104 29124
rect 30156 29112 30162 29164
rect 30653 29155 30711 29161
rect 30653 29121 30665 29155
rect 30699 29152 30711 29155
rect 31294 29152 31300 29164
rect 30699 29124 31300 29152
rect 30699 29121 30711 29124
rect 30653 29115 30711 29121
rect 27672 29056 27752 29084
rect 27672 29044 27678 29056
rect 28166 29044 28172 29096
rect 28224 29084 28230 29096
rect 30668 29084 30696 29115
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 31404 29152 31432 29183
rect 31478 29180 31484 29232
rect 31536 29220 31542 29232
rect 31589 29223 31647 29229
rect 31589 29220 31601 29223
rect 31536 29192 31601 29220
rect 31536 29180 31542 29192
rect 31589 29189 31601 29192
rect 31635 29220 31647 29223
rect 34054 29220 34060 29232
rect 31635 29192 32720 29220
rect 34015 29192 34060 29220
rect 31635 29189 31647 29192
rect 31589 29183 31647 29189
rect 32692 29161 32720 29192
rect 34054 29180 34060 29192
rect 34112 29180 34118 29232
rect 37182 29220 37188 29232
rect 35282 29192 37188 29220
rect 37182 29180 37188 29192
rect 37240 29180 37246 29232
rect 32492 29155 32550 29161
rect 32492 29152 32504 29155
rect 31404 29124 32504 29152
rect 28224 29056 30696 29084
rect 28224 29044 28230 29056
rect 23842 29016 23848 29028
rect 23584 28988 23848 29016
rect 23842 28976 23848 28988
rect 23900 29016 23906 29028
rect 26234 29016 26240 29028
rect 23900 28988 26240 29016
rect 23900 28976 23906 28988
rect 26234 28976 26240 28988
rect 26292 28976 26298 29028
rect 29822 28976 29828 29028
rect 29880 29016 29886 29028
rect 31404 29016 31432 29124
rect 32492 29121 32504 29124
rect 32538 29121 32550 29155
rect 32492 29115 32550 29121
rect 32677 29155 32735 29161
rect 32677 29121 32689 29155
rect 32723 29121 32735 29155
rect 36078 29152 36084 29164
rect 32677 29115 32735 29121
rect 35452 29124 36084 29152
rect 32306 29044 32312 29096
rect 32364 29084 32370 29096
rect 32401 29087 32459 29093
rect 32401 29084 32413 29087
rect 32364 29056 32413 29084
rect 32364 29044 32370 29056
rect 32401 29053 32413 29056
rect 32447 29053 32459 29087
rect 32401 29047 32459 29053
rect 32585 29087 32643 29093
rect 32585 29053 32597 29087
rect 32631 29053 32643 29087
rect 33778 29084 33784 29096
rect 33739 29056 33784 29084
rect 32585 29047 32643 29053
rect 29880 28988 31432 29016
rect 32600 29016 32628 29047
rect 33778 29044 33784 29056
rect 33836 29044 33842 29096
rect 35452 29084 35480 29124
rect 36078 29112 36084 29124
rect 36136 29112 36142 29164
rect 58069 29155 58127 29161
rect 58069 29121 58081 29155
rect 58115 29121 58127 29155
rect 58069 29115 58127 29121
rect 33888 29056 35480 29084
rect 32674 29016 32680 29028
rect 32600 28988 32680 29016
rect 29880 28976 29886 28988
rect 32674 28976 32680 28988
rect 32732 28976 32738 29028
rect 32861 29019 32919 29025
rect 32861 28985 32873 29019
rect 32907 29016 32919 29019
rect 33888 29016 33916 29056
rect 35526 29044 35532 29096
rect 35584 29084 35590 29096
rect 35805 29087 35863 29093
rect 35805 29084 35817 29087
rect 35584 29056 35817 29084
rect 35584 29044 35590 29056
rect 35805 29053 35817 29056
rect 35851 29084 35863 29087
rect 57425 29087 57483 29093
rect 57425 29084 57437 29087
rect 35851 29056 57437 29084
rect 35851 29053 35863 29056
rect 35805 29047 35863 29053
rect 57425 29053 57437 29056
rect 57471 29084 57483 29087
rect 58084 29084 58112 29115
rect 57471 29056 58112 29084
rect 57471 29053 57483 29056
rect 57425 29047 57483 29053
rect 32907 28988 33916 29016
rect 32907 28985 32919 28988
rect 32861 28979 32919 28985
rect 57882 28976 57888 29028
rect 57940 29016 57946 29028
rect 58253 29019 58311 29025
rect 58253 29016 58265 29019
rect 57940 28988 58265 29016
rect 57940 28976 57946 28988
rect 58253 28985 58265 28988
rect 58299 28985 58311 29019
rect 58253 28979 58311 28985
rect 19484 28920 19840 28948
rect 19484 28908 19490 28920
rect 23566 28908 23572 28960
rect 23624 28948 23630 28960
rect 23661 28951 23719 28957
rect 23661 28948 23673 28951
rect 23624 28920 23673 28948
rect 23624 28908 23630 28920
rect 23661 28917 23673 28920
rect 23707 28917 23719 28951
rect 23661 28911 23719 28917
rect 24765 28951 24823 28957
rect 24765 28917 24777 28951
rect 24811 28948 24823 28951
rect 25130 28948 25136 28960
rect 24811 28920 25136 28948
rect 24811 28917 24823 28920
rect 24765 28911 24823 28917
rect 25130 28908 25136 28920
rect 25188 28908 25194 28960
rect 30098 28948 30104 28960
rect 30059 28920 30104 28948
rect 30098 28908 30104 28920
rect 30156 28908 30162 28960
rect 30374 28908 30380 28960
rect 30432 28948 30438 28960
rect 31573 28951 31631 28957
rect 31573 28948 31585 28951
rect 30432 28920 31585 28948
rect 30432 28908 30438 28920
rect 31573 28917 31585 28920
rect 31619 28948 31631 28951
rect 32582 28948 32588 28960
rect 31619 28920 32588 28948
rect 31619 28917 31631 28920
rect 31573 28911 31631 28917
rect 32582 28908 32588 28920
rect 32640 28908 32646 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 19610 28744 19616 28756
rect 19571 28716 19616 28744
rect 19610 28704 19616 28716
rect 19668 28704 19674 28756
rect 20165 28747 20223 28753
rect 20165 28713 20177 28747
rect 20211 28744 20223 28747
rect 20211 28716 30788 28744
rect 20211 28713 20223 28716
rect 20165 28707 20223 28713
rect 16942 28636 16948 28688
rect 17000 28676 17006 28688
rect 17865 28679 17923 28685
rect 17865 28676 17877 28679
rect 17000 28648 17877 28676
rect 17000 28636 17006 28648
rect 17865 28645 17877 28648
rect 17911 28676 17923 28679
rect 25501 28679 25559 28685
rect 17911 28648 19380 28676
rect 17911 28645 17923 28648
rect 17865 28639 17923 28645
rect 18049 28611 18107 28617
rect 18049 28577 18061 28611
rect 18095 28608 18107 28611
rect 18095 28580 18644 28608
rect 18095 28577 18107 28580
rect 18049 28571 18107 28577
rect 18616 28549 18644 28580
rect 18601 28543 18659 28549
rect 18601 28509 18613 28543
rect 18647 28509 18659 28543
rect 18874 28540 18880 28552
rect 18787 28512 18880 28540
rect 18601 28503 18659 28509
rect 18874 28500 18880 28512
rect 18932 28540 18938 28552
rect 19242 28540 19248 28552
rect 18932 28512 19248 28540
rect 18932 28500 18938 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 19352 28540 19380 28648
rect 25501 28645 25513 28679
rect 25547 28676 25559 28679
rect 25590 28676 25596 28688
rect 25547 28648 25596 28676
rect 25547 28645 25559 28648
rect 25501 28639 25559 28645
rect 25590 28636 25596 28648
rect 25648 28676 25654 28688
rect 30760 28676 30788 28716
rect 31478 28676 31484 28688
rect 25648 28648 29960 28676
rect 30760 28648 31484 28676
rect 25648 28636 25654 28648
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28608 19947 28611
rect 20622 28608 20628 28620
rect 19935 28580 20628 28608
rect 19935 28577 19947 28580
rect 19889 28571 19947 28577
rect 20622 28568 20628 28580
rect 20680 28568 20686 28620
rect 23109 28611 23167 28617
rect 23109 28577 23121 28611
rect 23155 28577 23167 28611
rect 23566 28608 23572 28620
rect 23527 28580 23572 28608
rect 23109 28571 23167 28577
rect 19981 28543 20039 28549
rect 19981 28540 19993 28543
rect 19352 28512 19993 28540
rect 19981 28509 19993 28512
rect 20027 28509 20039 28543
rect 22278 28540 22284 28552
rect 22239 28512 22284 28540
rect 19981 28503 20039 28509
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 22462 28540 22468 28552
rect 22423 28512 22468 28540
rect 22462 28500 22468 28512
rect 22520 28540 22526 28552
rect 23124 28540 23152 28571
rect 23566 28568 23572 28580
rect 23624 28568 23630 28620
rect 26234 28608 26240 28620
rect 26195 28580 26240 28608
rect 26234 28568 26240 28580
rect 26292 28568 26298 28620
rect 29932 28617 29960 28648
rect 31478 28636 31484 28648
rect 31536 28636 31542 28688
rect 28261 28611 28319 28617
rect 28261 28577 28273 28611
rect 28307 28608 28319 28611
rect 29917 28611 29975 28617
rect 28307 28580 28856 28608
rect 28307 28577 28319 28580
rect 28261 28571 28319 28577
rect 22520 28512 23152 28540
rect 23477 28543 23535 28549
rect 22520 28500 22526 28512
rect 23477 28509 23489 28543
rect 23523 28540 23535 28543
rect 25038 28540 25044 28552
rect 23523 28512 25044 28540
rect 23523 28509 23535 28512
rect 23477 28503 23535 28509
rect 25038 28500 25044 28512
rect 25096 28500 25102 28552
rect 26252 28540 26280 28568
rect 26789 28543 26847 28549
rect 26789 28540 26801 28543
rect 26252 28512 26801 28540
rect 26789 28509 26801 28512
rect 26835 28540 26847 28543
rect 27614 28540 27620 28552
rect 26835 28512 27620 28540
rect 26835 28509 26847 28512
rect 26789 28503 26847 28509
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 28166 28540 28172 28552
rect 28079 28512 28172 28540
rect 17589 28475 17647 28481
rect 17589 28441 17601 28475
rect 17635 28472 17647 28475
rect 17862 28472 17868 28484
rect 17635 28444 17868 28472
rect 17635 28441 17647 28444
rect 17589 28435 17647 28441
rect 17862 28432 17868 28444
rect 17920 28472 17926 28484
rect 19521 28475 19579 28481
rect 19521 28472 19533 28475
rect 17920 28444 19533 28472
rect 17920 28432 17926 28444
rect 19521 28441 19533 28444
rect 19567 28441 19579 28475
rect 19521 28435 19579 28441
rect 20809 28475 20867 28481
rect 20809 28441 20821 28475
rect 20855 28472 20867 28475
rect 20898 28472 20904 28484
rect 20855 28444 20904 28472
rect 20855 28441 20867 28444
rect 20809 28435 20867 28441
rect 20898 28432 20904 28444
rect 20956 28432 20962 28484
rect 20990 28432 20996 28484
rect 21048 28472 21054 28484
rect 25130 28472 25136 28484
rect 21048 28444 21093 28472
rect 25091 28444 25136 28472
rect 21048 28432 21054 28444
rect 25130 28432 25136 28444
rect 25188 28432 25194 28484
rect 28092 28472 28120 28512
rect 28166 28500 28172 28512
rect 28224 28500 28230 28552
rect 28353 28543 28411 28549
rect 28353 28509 28365 28543
rect 28399 28540 28411 28543
rect 28534 28540 28540 28552
rect 28399 28512 28540 28540
rect 28399 28509 28411 28512
rect 28353 28503 28411 28509
rect 28534 28500 28540 28512
rect 28592 28500 28598 28552
rect 28828 28549 28856 28580
rect 29917 28577 29929 28611
rect 29963 28577 29975 28611
rect 29917 28571 29975 28577
rect 28813 28543 28871 28549
rect 28813 28509 28825 28543
rect 28859 28509 28871 28543
rect 28813 28503 28871 28509
rect 28997 28543 29055 28549
rect 28997 28509 29009 28543
rect 29043 28540 29055 28543
rect 29086 28540 29092 28552
rect 29043 28512 29092 28540
rect 29043 28509 29055 28512
rect 28997 28503 29055 28509
rect 29086 28500 29092 28512
rect 29144 28500 29150 28552
rect 30742 28500 30748 28552
rect 30800 28500 30806 28552
rect 30926 28500 30932 28552
rect 30984 28540 30990 28552
rect 32490 28540 32496 28552
rect 30984 28512 31029 28540
rect 32451 28512 32496 28540
rect 30984 28500 30990 28512
rect 32490 28500 32496 28512
rect 32548 28500 32554 28552
rect 32766 28540 32772 28552
rect 32727 28512 32772 28540
rect 32766 28500 32772 28512
rect 32824 28500 32830 28552
rect 33778 28500 33784 28552
rect 33836 28540 33842 28552
rect 33962 28540 33968 28552
rect 33836 28512 33968 28540
rect 33836 28500 33842 28512
rect 33962 28500 33968 28512
rect 34020 28540 34026 28552
rect 35253 28543 35311 28549
rect 35253 28540 35265 28543
rect 34020 28512 35265 28540
rect 34020 28500 34026 28512
rect 35253 28509 35265 28512
rect 35299 28509 35311 28543
rect 35253 28503 35311 28509
rect 29178 28472 29184 28484
rect 26988 28444 28120 28472
rect 28920 28444 29184 28472
rect 26988 28416 27016 28444
rect 18598 28404 18604 28416
rect 18559 28376 18604 28404
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 22373 28407 22431 28413
rect 22373 28404 22385 28407
rect 22336 28376 22385 28404
rect 22336 28364 22342 28376
rect 22373 28373 22385 28376
rect 22419 28373 22431 28407
rect 22373 28367 22431 28373
rect 25406 28364 25412 28416
rect 25464 28404 25470 28416
rect 25593 28407 25651 28413
rect 25593 28404 25605 28407
rect 25464 28376 25605 28404
rect 25464 28364 25470 28376
rect 25593 28373 25605 28376
rect 25639 28373 25651 28407
rect 26970 28404 26976 28416
rect 26931 28376 26976 28404
rect 25593 28367 25651 28373
rect 26970 28364 26976 28376
rect 27028 28364 27034 28416
rect 27522 28364 27528 28416
rect 27580 28404 27586 28416
rect 28920 28404 28948 28444
rect 29178 28432 29184 28444
rect 29236 28432 29242 28484
rect 30098 28432 30104 28484
rect 30156 28472 30162 28484
rect 32784 28472 32812 28500
rect 30156 28444 32812 28472
rect 33600 28484 33652 28490
rect 30156 28432 30162 28444
rect 35526 28472 35532 28484
rect 35487 28444 35532 28472
rect 35526 28432 35532 28444
rect 35584 28432 35590 28484
rect 37182 28472 37188 28484
rect 36754 28444 37188 28472
rect 37182 28432 37188 28444
rect 37240 28432 37246 28484
rect 37277 28475 37335 28481
rect 37277 28441 37289 28475
rect 37323 28472 37335 28475
rect 39482 28472 39488 28484
rect 37323 28444 39488 28472
rect 37323 28441 37335 28444
rect 37277 28435 37335 28441
rect 33600 28426 33652 28432
rect 27580 28376 28948 28404
rect 28997 28407 29055 28413
rect 27580 28364 27586 28376
rect 28997 28373 29009 28407
rect 29043 28404 29055 28407
rect 31110 28404 31116 28416
rect 29043 28376 31116 28404
rect 29043 28373 29055 28376
rect 28997 28367 29055 28373
rect 31110 28364 31116 28376
rect 31168 28364 31174 28416
rect 36538 28364 36544 28416
rect 36596 28404 36602 28416
rect 37292 28404 37320 28435
rect 39482 28432 39488 28444
rect 39540 28432 39546 28484
rect 36596 28376 37320 28404
rect 36596 28364 36602 28376
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 24857 28203 24915 28209
rect 24857 28169 24869 28203
rect 24903 28169 24915 28203
rect 24857 28163 24915 28169
rect 18877 28135 18935 28141
rect 18877 28101 18889 28135
rect 18923 28132 18935 28135
rect 19334 28132 19340 28144
rect 18923 28104 19340 28132
rect 18923 28101 18935 28104
rect 18877 28095 18935 28101
rect 19334 28092 19340 28104
rect 19392 28092 19398 28144
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 22244 28104 22416 28132
rect 22244 28092 22250 28104
rect 9858 28024 9864 28076
rect 9916 28064 9922 28076
rect 20073 28067 20131 28073
rect 20073 28064 20085 28067
rect 9916 28036 20085 28064
rect 9916 28024 9922 28036
rect 20073 28033 20085 28036
rect 20119 28033 20131 28067
rect 20898 28064 20904 28076
rect 20859 28036 20904 28064
rect 20073 28027 20131 28033
rect 20898 28024 20904 28036
rect 20956 28024 20962 28076
rect 22278 28064 22284 28076
rect 22239 28036 22284 28064
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22388 28064 22416 28104
rect 22462 28092 22468 28144
rect 22520 28132 22526 28144
rect 23293 28135 23351 28141
rect 23293 28132 23305 28135
rect 22520 28104 23305 28132
rect 22520 28092 22526 28104
rect 23293 28101 23305 28104
rect 23339 28101 23351 28135
rect 24872 28132 24900 28163
rect 28534 28160 28540 28212
rect 28592 28200 28598 28212
rect 29641 28203 29699 28209
rect 29641 28200 29653 28203
rect 28592 28172 29653 28200
rect 28592 28160 28598 28172
rect 29641 28169 29653 28172
rect 29687 28169 29699 28203
rect 29641 28163 29699 28169
rect 27157 28135 27215 28141
rect 24872 28104 25636 28132
rect 23293 28095 23351 28101
rect 23109 28067 23167 28073
rect 23109 28064 23121 28067
rect 22388 28036 23121 28064
rect 23109 28033 23121 28036
rect 23155 28033 23167 28067
rect 23109 28027 23167 28033
rect 24397 28067 24455 28073
rect 24397 28033 24409 28067
rect 24443 28064 24455 28067
rect 25130 28064 25136 28076
rect 24443 28036 25136 28064
rect 24443 28033 24455 28036
rect 24397 28027 24455 28033
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 25406 28064 25412 28076
rect 25367 28036 25412 28064
rect 25406 28024 25412 28036
rect 25464 28024 25470 28076
rect 25608 28073 25636 28104
rect 27157 28101 27169 28135
rect 27203 28132 27215 28135
rect 27614 28132 27620 28144
rect 27203 28104 27620 28132
rect 27203 28101 27215 28104
rect 27157 28095 27215 28101
rect 27614 28092 27620 28104
rect 27672 28092 27678 28144
rect 28905 28135 28963 28141
rect 28905 28101 28917 28135
rect 28951 28132 28963 28135
rect 28994 28132 29000 28144
rect 28951 28104 29000 28132
rect 28951 28101 28963 28104
rect 28905 28095 28963 28101
rect 28994 28092 29000 28104
rect 29052 28092 29058 28144
rect 29178 28092 29184 28144
rect 29236 28132 29242 28144
rect 31110 28132 31116 28144
rect 29236 28104 29946 28132
rect 31071 28104 31116 28132
rect 29236 28092 29242 28104
rect 31110 28092 31116 28104
rect 31168 28092 31174 28144
rect 34146 28132 34152 28144
rect 33994 28104 34152 28132
rect 34146 28092 34152 28104
rect 34204 28092 34210 28144
rect 34698 28092 34704 28144
rect 34756 28132 34762 28144
rect 34756 28104 35112 28132
rect 34756 28092 34762 28104
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 27522 28024 27528 28076
rect 27580 28064 27586 28076
rect 33134 28064 33140 28076
rect 27580 28036 27830 28064
rect 33095 28036 33140 28064
rect 27580 28024 27586 28036
rect 33134 28024 33140 28036
rect 33192 28024 33198 28076
rect 33594 28064 33600 28076
rect 33555 28036 33600 28064
rect 33594 28024 33600 28036
rect 33652 28024 33658 28076
rect 34790 28064 34796 28076
rect 34751 28036 34796 28064
rect 34790 28024 34796 28036
rect 34848 28024 34854 28076
rect 35084 28073 35112 28104
rect 34977 28067 35035 28073
rect 34977 28033 34989 28067
rect 35023 28033 35035 28067
rect 34977 28027 35035 28033
rect 35069 28067 35127 28073
rect 35069 28033 35081 28067
rect 35115 28033 35127 28067
rect 35069 28027 35127 28033
rect 35161 28067 35219 28073
rect 35161 28033 35173 28067
rect 35207 28064 35219 28067
rect 35618 28064 35624 28076
rect 35207 28036 35624 28064
rect 35207 28033 35219 28036
rect 35161 28027 35219 28033
rect 19242 27996 19248 28008
rect 19203 27968 19248 27996
rect 19242 27956 19248 27968
rect 19300 27956 19306 28008
rect 19337 27999 19395 28005
rect 19337 27965 19349 27999
rect 19383 27996 19395 27999
rect 19426 27996 19432 28008
rect 19383 27968 19432 27996
rect 19383 27965 19395 27968
rect 19337 27959 19395 27965
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 19521 27999 19579 28005
rect 19521 27965 19533 27999
rect 19567 27996 19579 27999
rect 20993 27999 21051 28005
rect 20993 27996 21005 27999
rect 19567 27968 21005 27996
rect 19567 27965 19579 27968
rect 19521 27959 19579 27965
rect 20993 27965 21005 27968
rect 21039 27996 21051 27999
rect 22189 27999 22247 28005
rect 22189 27996 22201 27999
rect 21039 27968 22201 27996
rect 21039 27965 21051 27968
rect 20993 27959 21051 27965
rect 22189 27965 22201 27968
rect 22235 27965 22247 27999
rect 22189 27959 22247 27965
rect 22649 27999 22707 28005
rect 22649 27965 22661 27999
rect 22695 27996 22707 27999
rect 23477 27999 23535 28005
rect 23477 27996 23489 27999
rect 22695 27968 23489 27996
rect 22695 27965 22707 27968
rect 22649 27959 22707 27965
rect 23477 27965 23489 27968
rect 23523 27996 23535 27999
rect 25317 27999 25375 28005
rect 25317 27996 25329 27999
rect 23523 27968 25329 27996
rect 23523 27965 23535 27968
rect 23477 27959 23535 27965
rect 25317 27965 25329 27968
rect 25363 27965 25375 27999
rect 25317 27959 25375 27965
rect 27246 27956 27252 28008
rect 27304 27996 27310 28008
rect 29181 27999 29239 28005
rect 29181 27996 29193 27999
rect 27304 27968 29193 27996
rect 27304 27956 27310 27968
rect 29181 27965 29193 27968
rect 29227 27996 29239 27999
rect 31389 27999 31447 28005
rect 31389 27996 31401 27999
rect 29227 27968 31401 27996
rect 29227 27965 29239 27968
rect 29181 27959 29239 27965
rect 31389 27965 31401 27968
rect 31435 27996 31447 27999
rect 31754 27996 31760 28008
rect 31435 27968 31760 27996
rect 31435 27965 31447 27968
rect 31389 27959 31447 27965
rect 31754 27956 31760 27968
rect 31812 27996 31818 28008
rect 32398 27996 32404 28008
rect 31812 27968 32404 27996
rect 31812 27956 31818 27968
rect 32398 27956 32404 27968
rect 32456 27956 32462 28008
rect 34992 27996 35020 28027
rect 35618 28024 35624 28036
rect 35676 28064 35682 28076
rect 35897 28067 35955 28073
rect 35897 28064 35909 28067
rect 35676 28036 35909 28064
rect 35676 28024 35682 28036
rect 35897 28033 35909 28036
rect 35943 28033 35955 28067
rect 35897 28027 35955 28033
rect 35342 27996 35348 28008
rect 34992 27968 35348 27996
rect 35342 27956 35348 27968
rect 35400 27956 35406 28008
rect 21358 27820 21364 27872
rect 21416 27860 21422 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21416 27832 22017 27860
rect 21416 27820 21422 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 24673 27863 24731 27869
rect 24673 27829 24685 27863
rect 24719 27860 24731 27863
rect 25590 27860 25596 27872
rect 24719 27832 25596 27860
rect 24719 27829 24731 27832
rect 24673 27823 24731 27829
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 25777 27863 25835 27869
rect 25777 27829 25789 27863
rect 25823 27860 25835 27863
rect 29822 27860 29828 27872
rect 25823 27832 29828 27860
rect 25823 27829 25835 27832
rect 25777 27823 25835 27829
rect 29822 27820 29828 27832
rect 29880 27820 29886 27872
rect 35434 27860 35440 27872
rect 35395 27832 35440 27860
rect 35434 27820 35440 27832
rect 35492 27820 35498 27872
rect 36446 27860 36452 27872
rect 36407 27832 36452 27860
rect 36446 27820 36452 27832
rect 36504 27820 36510 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 28166 27616 28172 27668
rect 28224 27656 28230 27668
rect 28353 27659 28411 27665
rect 28353 27656 28365 27659
rect 28224 27628 28365 27656
rect 28224 27616 28230 27628
rect 28353 27625 28365 27628
rect 28399 27625 28411 27659
rect 28353 27619 28411 27625
rect 35434 27616 35440 27668
rect 35492 27656 35498 27668
rect 36154 27659 36212 27665
rect 36154 27656 36166 27659
rect 35492 27628 36166 27656
rect 35492 27616 35498 27628
rect 36154 27625 36166 27628
rect 36200 27625 36212 27659
rect 36154 27619 36212 27625
rect 2866 27548 2872 27600
rect 2924 27588 2930 27600
rect 26329 27591 26387 27597
rect 26329 27588 26341 27591
rect 2924 27560 26341 27588
rect 2924 27548 2930 27560
rect 26329 27557 26341 27560
rect 26375 27557 26387 27591
rect 26329 27551 26387 27557
rect 22186 27480 22192 27532
rect 22244 27520 22250 27532
rect 22281 27523 22339 27529
rect 22281 27520 22293 27523
rect 22244 27492 22293 27520
rect 22244 27480 22250 27492
rect 22281 27489 22293 27492
rect 22327 27489 22339 27523
rect 22281 27483 22339 27489
rect 20622 27452 20628 27464
rect 20583 27424 20628 27452
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 22373 27455 22431 27461
rect 22373 27421 22385 27455
rect 22419 27452 22431 27455
rect 22462 27452 22468 27464
rect 22419 27424 22468 27452
rect 22419 27421 22431 27424
rect 22373 27415 22431 27421
rect 22462 27412 22468 27424
rect 22520 27412 22526 27464
rect 23201 27455 23259 27461
rect 23201 27421 23213 27455
rect 23247 27452 23259 27455
rect 23661 27455 23719 27461
rect 23661 27452 23673 27455
rect 23247 27424 23673 27452
rect 23247 27421 23259 27424
rect 23201 27415 23259 27421
rect 23661 27421 23673 27424
rect 23707 27452 23719 27455
rect 24026 27452 24032 27464
rect 23707 27424 24032 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 25130 27412 25136 27464
rect 25188 27412 25194 27464
rect 25590 27412 25596 27464
rect 25648 27452 25654 27464
rect 26344 27452 26372 27551
rect 26970 27548 26976 27600
rect 27028 27588 27034 27600
rect 30374 27588 30380 27600
rect 27028 27560 30380 27588
rect 27028 27548 27034 27560
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 30742 27588 30748 27600
rect 30703 27560 30748 27588
rect 30742 27548 30748 27560
rect 30800 27548 30806 27600
rect 33226 27588 33232 27600
rect 31726 27560 33232 27588
rect 26881 27523 26939 27529
rect 26881 27489 26893 27523
rect 26927 27520 26939 27523
rect 28997 27523 29055 27529
rect 28997 27520 29009 27523
rect 26927 27492 29009 27520
rect 26927 27489 26939 27492
rect 26881 27483 26939 27489
rect 28997 27489 29009 27492
rect 29043 27520 29055 27523
rect 31726 27520 31754 27560
rect 33226 27548 33232 27560
rect 33284 27548 33290 27600
rect 29043 27492 31754 27520
rect 29043 27489 29055 27492
rect 28997 27483 29055 27489
rect 27065 27455 27123 27461
rect 27065 27452 27077 27455
rect 25648 27424 25693 27452
rect 26344 27424 27077 27452
rect 25648 27412 25654 27424
rect 27065 27421 27077 27424
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 27249 27455 27307 27461
rect 27249 27421 27261 27455
rect 27295 27452 27307 27455
rect 27893 27455 27951 27461
rect 27893 27452 27905 27455
rect 27295 27424 27905 27452
rect 27295 27421 27307 27424
rect 27249 27415 27307 27421
rect 27893 27421 27905 27424
rect 27939 27421 27951 27455
rect 30653 27455 30711 27461
rect 30653 27452 30665 27455
rect 27893 27415 27951 27421
rect 30116 27424 30665 27452
rect 19334 27344 19340 27396
rect 19392 27384 19398 27396
rect 20809 27387 20867 27393
rect 20809 27384 20821 27387
rect 19392 27356 20821 27384
rect 19392 27344 19398 27356
rect 20809 27353 20821 27356
rect 20855 27353 20867 27387
rect 20809 27347 20867 27353
rect 20993 27387 21051 27393
rect 20993 27353 21005 27387
rect 21039 27384 21051 27387
rect 24578 27384 24584 27396
rect 21039 27356 24440 27384
rect 24539 27356 24584 27384
rect 21039 27353 21051 27356
rect 20993 27347 21051 27353
rect 20898 27276 20904 27328
rect 20956 27316 20962 27328
rect 22005 27319 22063 27325
rect 22005 27316 22017 27319
rect 20956 27288 22017 27316
rect 20956 27276 20962 27288
rect 22005 27285 22017 27288
rect 22051 27285 22063 27319
rect 23842 27316 23848 27328
rect 23803 27288 23848 27316
rect 22005 27279 22063 27285
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 24412 27316 24440 27356
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 26970 27316 26976 27328
rect 24412 27288 26976 27316
rect 26970 27276 26976 27288
rect 27028 27276 27034 27328
rect 27430 27276 27436 27328
rect 27488 27316 27494 27328
rect 27709 27319 27767 27325
rect 27709 27316 27721 27319
rect 27488 27288 27721 27316
rect 27488 27276 27494 27288
rect 27709 27285 27721 27288
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 28166 27276 28172 27328
rect 28224 27316 28230 27328
rect 30116 27325 30144 27424
rect 30653 27421 30665 27424
rect 30699 27421 30711 27455
rect 30653 27415 30711 27421
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27452 30895 27455
rect 31018 27452 31024 27464
rect 30883 27424 31024 27452
rect 30883 27421 30895 27424
rect 30837 27415 30895 27421
rect 31018 27412 31024 27424
rect 31076 27412 31082 27464
rect 31294 27452 31300 27464
rect 31255 27424 31300 27452
rect 31294 27412 31300 27424
rect 31352 27412 31358 27464
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 32600 27424 34161 27452
rect 30101 27319 30159 27325
rect 30101 27316 30113 27319
rect 28224 27288 30113 27316
rect 28224 27276 28230 27288
rect 30101 27285 30113 27288
rect 30147 27285 30159 27319
rect 31478 27316 31484 27328
rect 31439 27288 31484 27316
rect 30101 27279 30159 27285
rect 31478 27276 31484 27288
rect 31536 27276 31542 27328
rect 31938 27276 31944 27328
rect 31996 27316 32002 27328
rect 32600 27325 32628 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34333 27455 34391 27461
rect 34333 27421 34345 27455
rect 34379 27452 34391 27455
rect 35894 27452 35900 27464
rect 34379 27424 35296 27452
rect 35855 27424 35900 27452
rect 34379 27421 34391 27424
rect 34333 27415 34391 27421
rect 34164 27384 34192 27415
rect 35268 27393 35296 27424
rect 35894 27412 35900 27424
rect 35952 27412 35958 27464
rect 35069 27387 35127 27393
rect 35069 27384 35081 27387
rect 34164 27356 35081 27384
rect 35069 27353 35081 27356
rect 35115 27353 35127 27387
rect 35069 27347 35127 27353
rect 35253 27387 35311 27393
rect 35253 27353 35265 27387
rect 35299 27384 35311 27387
rect 35342 27384 35348 27396
rect 35299 27356 35348 27384
rect 35299 27353 35311 27356
rect 35253 27347 35311 27353
rect 32585 27319 32643 27325
rect 32585 27316 32597 27319
rect 31996 27288 32597 27316
rect 31996 27276 32002 27288
rect 32585 27285 32597 27288
rect 32631 27285 32643 27319
rect 33226 27316 33232 27328
rect 33139 27288 33232 27316
rect 32585 27279 32643 27285
rect 33226 27276 33232 27288
rect 33284 27316 33290 27328
rect 33778 27316 33784 27328
rect 33284 27288 33784 27316
rect 33284 27276 33290 27288
rect 33778 27276 33784 27288
rect 33836 27276 33842 27328
rect 34238 27316 34244 27328
rect 34199 27288 34244 27316
rect 34238 27276 34244 27288
rect 34296 27276 34302 27328
rect 34698 27276 34704 27328
rect 34756 27316 34762 27328
rect 34885 27319 34943 27325
rect 34885 27316 34897 27319
rect 34756 27288 34897 27316
rect 34756 27276 34762 27288
rect 34885 27285 34897 27288
rect 34931 27285 34943 27319
rect 35084 27316 35112 27347
rect 35342 27344 35348 27356
rect 35400 27344 35406 27396
rect 37182 27344 37188 27396
rect 37240 27344 37246 27396
rect 37918 27384 37924 27396
rect 37879 27356 37924 27384
rect 37918 27344 37924 27356
rect 37976 27344 37982 27396
rect 38378 27384 38384 27396
rect 38339 27356 38384 27384
rect 38378 27344 38384 27356
rect 38436 27344 38442 27396
rect 36446 27316 36452 27328
rect 35084 27288 36452 27316
rect 34885 27279 34943 27285
rect 36446 27276 36452 27288
rect 36504 27276 36510 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 24578 27112 24584 27124
rect 21284 27084 24584 27112
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 21284 27044 21312 27084
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 24673 27115 24731 27121
rect 24673 27081 24685 27115
rect 24719 27112 24731 27115
rect 27154 27112 27160 27124
rect 24719 27084 27160 27112
rect 24719 27081 24731 27084
rect 24673 27075 24731 27081
rect 21048 27016 21312 27044
rect 21048 27004 21054 27016
rect 21192 26985 21220 27016
rect 23382 27004 23388 27056
rect 23440 27004 23446 27056
rect 23845 27047 23903 27053
rect 23845 27013 23857 27047
rect 23891 27044 23903 27047
rect 24688 27044 24716 27075
rect 27154 27072 27160 27084
rect 27212 27112 27218 27124
rect 30009 27115 30067 27121
rect 30009 27112 30021 27115
rect 27212 27084 30021 27112
rect 27212 27072 27218 27084
rect 30009 27081 30021 27084
rect 30055 27081 30067 27115
rect 34606 27112 34612 27124
rect 30009 27075 30067 27081
rect 34072 27084 34612 27112
rect 27430 27044 27436 27056
rect 23891 27016 24716 27044
rect 27391 27016 27436 27044
rect 23891 27013 23903 27016
rect 23845 27007 23903 27013
rect 27430 27004 27436 27016
rect 27488 27004 27494 27056
rect 27522 27004 27528 27056
rect 27580 27044 27586 27056
rect 31202 27044 31208 27056
rect 27580 27016 27922 27044
rect 31050 27016 31208 27044
rect 27580 27004 27586 27016
rect 31202 27004 31208 27016
rect 31260 27004 31266 27056
rect 31478 27044 31484 27056
rect 31439 27016 31484 27044
rect 31478 27004 31484 27016
rect 31536 27004 31542 27056
rect 34072 27053 34100 27084
rect 34606 27072 34612 27084
rect 34664 27112 34670 27124
rect 35345 27115 35403 27121
rect 34664 27084 35020 27112
rect 34664 27072 34670 27084
rect 34057 27047 34115 27053
rect 34057 27013 34069 27047
rect 34103 27013 34115 27047
rect 34057 27007 34115 27013
rect 34238 27004 34244 27056
rect 34296 27044 34302 27056
rect 34296 27016 34928 27044
rect 34296 27004 34302 27016
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26945 21235 26979
rect 21358 26976 21364 26988
rect 21319 26948 21364 26976
rect 21177 26939 21235 26945
rect 21358 26936 21364 26948
rect 21416 26936 21422 26988
rect 31754 26936 31760 26988
rect 31812 26976 31818 26988
rect 32861 26979 32919 26985
rect 31812 26948 31857 26976
rect 31812 26936 31818 26948
rect 32861 26945 32873 26979
rect 32907 26976 32919 26979
rect 33778 26976 33784 26988
rect 32907 26948 33784 26976
rect 32907 26945 32919 26948
rect 32861 26939 32919 26945
rect 33778 26936 33784 26948
rect 33836 26936 33842 26988
rect 33962 26976 33968 26988
rect 33923 26948 33968 26976
rect 33962 26936 33968 26948
rect 34020 26936 34026 26988
rect 34698 26976 34704 26988
rect 34659 26948 34704 26976
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 34900 26985 34928 27016
rect 34992 26985 35020 27084
rect 35345 27081 35357 27115
rect 35391 27112 35403 27115
rect 35526 27112 35532 27124
rect 35391 27084 35532 27112
rect 35391 27081 35403 27084
rect 35345 27075 35403 27081
rect 35526 27072 35532 27084
rect 35584 27072 35590 27124
rect 36906 27072 36912 27124
rect 36964 27112 36970 27124
rect 37182 27112 37188 27124
rect 36964 27084 37188 27112
rect 36964 27072 36970 27084
rect 37182 27072 37188 27084
rect 37240 27112 37246 27124
rect 37461 27115 37519 27121
rect 37461 27112 37473 27115
rect 37240 27084 37473 27112
rect 37240 27072 37246 27084
rect 37461 27081 37473 27084
rect 37507 27081 37519 27115
rect 39482 27112 39488 27124
rect 39443 27084 39488 27112
rect 37461 27075 37519 27081
rect 39482 27072 39488 27084
rect 39540 27072 39546 27124
rect 34885 26979 34943 26985
rect 34885 26945 34897 26979
rect 34931 26945 34943 26979
rect 34885 26939 34943 26945
rect 34977 26979 35035 26985
rect 34977 26945 34989 26979
rect 35023 26945 35035 26979
rect 34977 26939 35035 26945
rect 35069 26979 35127 26985
rect 35069 26945 35081 26979
rect 35115 26976 35127 26979
rect 35434 26976 35440 26988
rect 35115 26948 35440 26976
rect 35115 26945 35127 26948
rect 35069 26939 35127 26945
rect 20438 26908 20444 26920
rect 20399 26880 20444 26908
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 24121 26911 24179 26917
rect 24121 26877 24133 26911
rect 24167 26908 24179 26911
rect 24578 26908 24584 26920
rect 24167 26880 24584 26908
rect 24167 26877 24179 26880
rect 24121 26871 24179 26877
rect 24578 26868 24584 26880
rect 24636 26868 24642 26920
rect 27154 26908 27160 26920
rect 27115 26880 27160 26908
rect 27154 26868 27160 26880
rect 27212 26868 27218 26920
rect 32677 26911 32735 26917
rect 32677 26877 32689 26911
rect 32723 26908 32735 26911
rect 33980 26908 34008 26936
rect 32723 26880 34008 26908
rect 34992 26908 35020 26939
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 36265 26979 36323 26985
rect 36265 26945 36277 26979
rect 36311 26976 36323 26979
rect 36924 26976 36952 27072
rect 36311 26948 36952 26976
rect 36311 26945 36323 26948
rect 36265 26939 36323 26945
rect 38378 26936 38384 26988
rect 38436 26976 38442 26988
rect 38473 26979 38531 26985
rect 38473 26976 38485 26979
rect 38436 26948 38485 26976
rect 38436 26936 38442 26948
rect 38473 26945 38485 26948
rect 38519 26945 38531 26979
rect 38473 26939 38531 26945
rect 35526 26908 35532 26920
rect 34992 26880 35532 26908
rect 32723 26877 32735 26880
rect 32677 26871 32735 26877
rect 35526 26868 35532 26880
rect 35584 26868 35590 26920
rect 38289 26911 38347 26917
rect 38289 26877 38301 26911
rect 38335 26908 38347 26911
rect 38838 26908 38844 26920
rect 38335 26880 38844 26908
rect 38335 26877 38347 26880
rect 38289 26871 38347 26877
rect 38838 26868 38844 26880
rect 38896 26868 38902 26920
rect 43990 26868 43996 26920
rect 44048 26908 44054 26920
rect 57606 26908 57612 26920
rect 44048 26880 57612 26908
rect 44048 26868 44054 26880
rect 57606 26868 57612 26880
rect 57664 26868 57670 26920
rect 33778 26800 33784 26852
rect 33836 26840 33842 26852
rect 34054 26840 34060 26852
rect 33836 26812 34060 26840
rect 33836 26800 33842 26812
rect 34054 26800 34060 26812
rect 34112 26840 34118 26852
rect 34112 26812 36860 26840
rect 34112 26800 34118 26812
rect 36832 26784 36860 26812
rect 39482 26800 39488 26852
rect 39540 26840 39546 26852
rect 57146 26840 57152 26852
rect 39540 26812 57152 26840
rect 39540 26800 39546 26812
rect 57146 26800 57152 26812
rect 57204 26800 57210 26852
rect 22373 26775 22431 26781
rect 22373 26741 22385 26775
rect 22419 26772 22431 26775
rect 24210 26772 24216 26784
rect 22419 26744 24216 26772
rect 22419 26741 22431 26744
rect 22373 26735 22431 26741
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 28905 26775 28963 26781
rect 28905 26741 28917 26775
rect 28951 26772 28963 26775
rect 29454 26772 29460 26784
rect 28951 26744 29460 26772
rect 28951 26741 28963 26744
rect 28905 26735 28963 26741
rect 29454 26732 29460 26744
rect 29512 26732 29518 26784
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33226 26772 33232 26784
rect 33091 26744 33232 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33226 26732 33232 26744
rect 33284 26732 33290 26784
rect 35894 26732 35900 26784
rect 35952 26772 35958 26784
rect 36081 26775 36139 26781
rect 36081 26772 36093 26775
rect 35952 26744 36093 26772
rect 35952 26732 35958 26744
rect 36081 26741 36093 26744
rect 36127 26741 36139 26775
rect 36814 26772 36820 26784
rect 36775 26744 36820 26772
rect 36081 26735 36139 26741
rect 36814 26732 36820 26744
rect 36872 26732 36878 26784
rect 38746 26732 38752 26784
rect 38804 26772 38810 26784
rect 38933 26775 38991 26781
rect 38933 26772 38945 26775
rect 38804 26744 38945 26772
rect 38804 26732 38810 26744
rect 38933 26741 38945 26744
rect 38979 26741 38991 26775
rect 41874 26772 41880 26784
rect 41835 26744 41880 26772
rect 38933 26735 38991 26741
rect 41874 26732 41880 26744
rect 41932 26772 41938 26784
rect 42797 26775 42855 26781
rect 42797 26772 42809 26775
rect 41932 26744 42809 26772
rect 41932 26732 41938 26744
rect 42797 26741 42809 26744
rect 42843 26741 42855 26775
rect 42797 26735 42855 26741
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 23382 26528 23388 26580
rect 23440 26568 23446 26580
rect 23661 26571 23719 26577
rect 23661 26568 23673 26571
rect 23440 26540 23673 26568
rect 23440 26528 23446 26540
rect 23661 26537 23673 26540
rect 23707 26537 23719 26571
rect 23661 26531 23719 26537
rect 23676 26296 23704 26531
rect 23842 26528 23848 26580
rect 23900 26568 23906 26580
rect 30009 26571 30067 26577
rect 23900 26540 28948 26568
rect 23900 26528 23906 26540
rect 23952 26373 23980 26540
rect 27430 26460 27436 26512
rect 27488 26460 27494 26512
rect 24578 26432 24584 26444
rect 24491 26404 24584 26432
rect 24578 26392 24584 26404
rect 24636 26432 24642 26444
rect 26326 26432 26332 26444
rect 24636 26404 26332 26432
rect 24636 26392 24642 26404
rect 26326 26392 26332 26404
rect 26384 26392 26390 26444
rect 26605 26435 26663 26441
rect 26605 26401 26617 26435
rect 26651 26432 26663 26435
rect 26786 26432 26792 26444
rect 26651 26404 26792 26432
rect 26651 26401 26663 26404
rect 26605 26395 26663 26401
rect 26786 26392 26792 26404
rect 26844 26392 26850 26444
rect 27448 26432 27476 26460
rect 27709 26435 27767 26441
rect 27709 26432 27721 26435
rect 27448 26404 27721 26432
rect 27709 26401 27721 26404
rect 27755 26401 27767 26435
rect 27709 26395 27767 26401
rect 23937 26367 23995 26373
rect 23937 26333 23949 26367
rect 23983 26364 23995 26367
rect 24118 26364 24124 26376
rect 23983 26336 24124 26364
rect 23983 26333 23995 26336
rect 23937 26327 23995 26333
rect 24118 26324 24124 26336
rect 24176 26324 24182 26376
rect 27062 26324 27068 26376
rect 27120 26364 27126 26376
rect 27433 26367 27491 26373
rect 27433 26364 27445 26367
rect 27120 26336 27445 26364
rect 27120 26324 27126 26336
rect 27433 26333 27445 26336
rect 27479 26333 27491 26367
rect 28920 26364 28948 26540
rect 30009 26537 30021 26571
rect 30055 26568 30067 26571
rect 31294 26568 31300 26580
rect 30055 26540 31300 26568
rect 30055 26537 30067 26540
rect 30009 26531 30067 26537
rect 31294 26528 31300 26540
rect 31352 26528 31358 26580
rect 33410 26568 33416 26580
rect 33371 26540 33416 26568
rect 33410 26528 33416 26540
rect 33468 26528 33474 26580
rect 34149 26571 34207 26577
rect 34149 26537 34161 26571
rect 34195 26568 34207 26571
rect 34790 26568 34796 26580
rect 34195 26540 34796 26568
rect 34195 26537 34207 26540
rect 34149 26531 34207 26537
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 35253 26571 35311 26577
rect 35253 26537 35265 26571
rect 35299 26568 35311 26571
rect 35342 26568 35348 26580
rect 35299 26540 35348 26568
rect 35299 26537 35311 26540
rect 35253 26531 35311 26537
rect 35342 26528 35348 26540
rect 35400 26528 35406 26580
rect 36170 26568 36176 26580
rect 35452 26540 36176 26568
rect 29181 26503 29239 26509
rect 29181 26469 29193 26503
rect 29227 26500 29239 26503
rect 30101 26503 30159 26509
rect 30101 26500 30113 26503
rect 29227 26472 30113 26500
rect 29227 26469 29239 26472
rect 29181 26463 29239 26469
rect 30101 26469 30113 26472
rect 30147 26469 30159 26503
rect 31941 26503 31999 26509
rect 31941 26500 31953 26503
rect 30101 26463 30159 26469
rect 31726 26472 31953 26500
rect 30466 26432 30472 26444
rect 30427 26404 30472 26432
rect 30466 26392 30472 26404
rect 30524 26392 30530 26444
rect 31021 26367 31079 26373
rect 31021 26364 31033 26367
rect 28920 26336 31033 26364
rect 27433 26327 27491 26333
rect 31021 26333 31033 26336
rect 31067 26364 31079 26367
rect 31726 26364 31754 26472
rect 31941 26469 31953 26472
rect 31987 26500 31999 26503
rect 35452 26500 35480 26540
rect 36170 26528 36176 26540
rect 36228 26528 36234 26580
rect 37182 26528 37188 26580
rect 37240 26568 37246 26580
rect 58158 26568 58164 26580
rect 37240 26540 58164 26568
rect 37240 26528 37246 26540
rect 58158 26528 58164 26540
rect 58216 26528 58222 26580
rect 31987 26472 35480 26500
rect 39393 26503 39451 26509
rect 31987 26469 31999 26472
rect 31941 26463 31999 26469
rect 39393 26469 39405 26503
rect 39439 26500 39451 26503
rect 40218 26500 40224 26512
rect 39439 26472 40224 26500
rect 39439 26469 39451 26472
rect 39393 26463 39451 26469
rect 40218 26460 40224 26472
rect 40276 26460 40282 26512
rect 33962 26392 33968 26444
rect 34020 26432 34026 26444
rect 35805 26435 35863 26441
rect 35805 26432 35817 26435
rect 34020 26404 35817 26432
rect 34020 26392 34026 26404
rect 35805 26401 35817 26404
rect 35851 26401 35863 26435
rect 35805 26395 35863 26401
rect 33226 26364 33232 26376
rect 31067 26336 31754 26364
rect 33187 26336 33232 26364
rect 31067 26333 31079 26336
rect 31021 26327 31079 26333
rect 33226 26324 33232 26336
rect 33284 26324 33290 26376
rect 34057 26367 34115 26373
rect 34057 26333 34069 26367
rect 34103 26333 34115 26367
rect 34057 26327 34115 26333
rect 34241 26367 34299 26373
rect 34241 26333 34253 26367
rect 34287 26364 34299 26367
rect 34330 26364 34336 26376
rect 34287 26336 34336 26364
rect 34287 26333 34299 26336
rect 34241 26327 34299 26333
rect 23676 26268 24164 26296
rect 24136 26228 24164 26268
rect 24210 26256 24216 26308
rect 24268 26296 24274 26308
rect 24857 26299 24915 26305
rect 24857 26296 24869 26299
rect 24268 26268 24869 26296
rect 24268 26256 24274 26268
rect 24857 26265 24869 26268
rect 24903 26265 24915 26299
rect 27338 26296 27344 26308
rect 24857 26259 24915 26265
rect 24964 26268 25346 26296
rect 26160 26268 27344 26296
rect 24964 26228 24992 26268
rect 24136 26200 24992 26228
rect 25240 26228 25268 26268
rect 26160 26228 26188 26268
rect 27338 26256 27344 26268
rect 27396 26296 27402 26308
rect 27396 26268 28198 26296
rect 27396 26256 27402 26268
rect 31202 26256 31208 26308
rect 31260 26296 31266 26308
rect 31389 26299 31447 26305
rect 31389 26296 31401 26299
rect 31260 26268 31401 26296
rect 31260 26256 31266 26268
rect 31389 26265 31401 26268
rect 31435 26296 31447 26299
rect 32582 26296 32588 26308
rect 31435 26268 32588 26296
rect 31435 26265 31447 26268
rect 31389 26259 31447 26265
rect 32582 26256 32588 26268
rect 32640 26256 32646 26308
rect 32677 26299 32735 26305
rect 32677 26265 32689 26299
rect 32723 26265 32735 26299
rect 34072 26296 34100 26327
rect 34330 26324 34336 26336
rect 34388 26364 34394 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34388 26336 34897 26364
rect 34388 26324 34394 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 34790 26296 34796 26308
rect 34072 26268 34796 26296
rect 32677 26259 32735 26265
rect 25240 26200 26188 26228
rect 30650 26188 30656 26240
rect 30708 26228 30714 26240
rect 32692 26228 32720 26259
rect 34790 26256 34796 26268
rect 34848 26296 34854 26308
rect 35069 26299 35127 26305
rect 35069 26296 35081 26299
rect 34848 26268 35081 26296
rect 34848 26256 34854 26268
rect 35069 26265 35081 26268
rect 35115 26265 35127 26299
rect 35820 26296 35848 26395
rect 37274 26392 37280 26444
rect 37332 26392 37338 26444
rect 37829 26435 37887 26441
rect 37829 26401 37841 26435
rect 37875 26432 37887 26435
rect 38378 26432 38384 26444
rect 37875 26404 38384 26432
rect 37875 26401 37887 26404
rect 37829 26395 37887 26401
rect 38378 26392 38384 26404
rect 38436 26432 38442 26444
rect 40129 26435 40187 26441
rect 40129 26432 40141 26435
rect 38436 26404 40141 26432
rect 38436 26392 38442 26404
rect 40129 26401 40141 26404
rect 40175 26401 40187 26435
rect 40129 26395 40187 26401
rect 37292 26364 37320 26392
rect 39206 26364 39212 26376
rect 37214 26336 37320 26364
rect 39167 26336 39212 26364
rect 39206 26324 39212 26336
rect 39264 26324 39270 26376
rect 40034 26324 40040 26376
rect 40092 26364 40098 26376
rect 41141 26367 41199 26373
rect 41141 26364 41153 26367
rect 40092 26336 41153 26364
rect 40092 26324 40098 26336
rect 41141 26333 41153 26336
rect 41187 26333 41199 26367
rect 41141 26327 41199 26333
rect 41874 26324 41880 26376
rect 41932 26364 41938 26376
rect 42521 26367 42579 26373
rect 42521 26364 42533 26367
rect 41932 26336 42533 26364
rect 41932 26324 41938 26336
rect 42521 26333 42533 26336
rect 42567 26364 42579 26367
rect 42981 26367 43039 26373
rect 42981 26364 42993 26367
rect 42567 26336 42993 26364
rect 42567 26333 42579 26336
rect 42521 26327 42579 26333
rect 42981 26333 42993 26336
rect 43027 26333 43039 26367
rect 42981 26327 43039 26333
rect 36078 26296 36084 26308
rect 35820 26268 35940 26296
rect 36039 26268 36084 26296
rect 35069 26259 35127 26265
rect 35912 26240 35940 26268
rect 36078 26256 36084 26268
rect 36136 26256 36142 26308
rect 38010 26256 38016 26308
rect 38068 26296 38074 26308
rect 38289 26299 38347 26305
rect 38289 26296 38301 26299
rect 38068 26268 38301 26296
rect 38068 26256 38074 26268
rect 38289 26265 38301 26268
rect 38335 26265 38347 26299
rect 38289 26259 38347 26265
rect 38657 26299 38715 26305
rect 38657 26265 38669 26299
rect 38703 26296 38715 26299
rect 38746 26296 38752 26308
rect 38703 26268 38752 26296
rect 38703 26265 38715 26268
rect 38657 26259 38715 26265
rect 38746 26256 38752 26268
rect 38804 26256 38810 26308
rect 41046 26256 41052 26308
rect 41104 26296 41110 26308
rect 42245 26299 42303 26305
rect 42245 26296 42257 26299
rect 41104 26268 42257 26296
rect 41104 26256 41110 26268
rect 42245 26265 42257 26268
rect 42291 26296 42303 26299
rect 43257 26299 43315 26305
rect 42291 26268 43116 26296
rect 42291 26265 42303 26268
rect 42245 26259 42303 26265
rect 33870 26228 33876 26240
rect 30708 26200 33876 26228
rect 30708 26188 30714 26200
rect 33870 26188 33876 26200
rect 33928 26188 33934 26240
rect 35894 26188 35900 26240
rect 35952 26188 35958 26240
rect 40126 26188 40132 26240
rect 40184 26228 40190 26240
rect 40589 26231 40647 26237
rect 40589 26228 40601 26231
rect 40184 26200 40601 26228
rect 40184 26188 40190 26200
rect 40589 26197 40601 26200
rect 40635 26197 40647 26231
rect 43088 26228 43116 26268
rect 43257 26265 43269 26299
rect 43303 26296 43315 26299
rect 43438 26296 43444 26308
rect 43303 26268 43444 26296
rect 43303 26265 43315 26268
rect 43257 26259 43315 26265
rect 43438 26256 43444 26268
rect 43496 26256 43502 26308
rect 44818 26228 44824 26240
rect 43088 26200 44824 26228
rect 40589 26191 40647 26197
rect 44818 26188 44824 26200
rect 44876 26188 44882 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 24118 26024 24124 26036
rect 24079 25996 24124 26024
rect 24118 25984 24124 25996
rect 24176 25984 24182 26036
rect 26605 26027 26663 26033
rect 26605 25993 26617 26027
rect 26651 26024 26663 26027
rect 27154 26024 27160 26036
rect 26651 25996 27160 26024
rect 26651 25993 26663 25996
rect 26605 25987 26663 25993
rect 27154 25984 27160 25996
rect 27212 25984 27218 26036
rect 30466 25984 30472 26036
rect 30524 26024 30530 26036
rect 31389 26027 31447 26033
rect 31389 26024 31401 26027
rect 30524 25996 31401 26024
rect 30524 25984 30530 25996
rect 31389 25993 31401 25996
rect 31435 25993 31447 26027
rect 31389 25987 31447 25993
rect 33137 26027 33195 26033
rect 33137 25993 33149 26027
rect 33183 26024 33195 26027
rect 33410 26024 33416 26036
rect 33183 25996 33416 26024
rect 33183 25993 33195 25996
rect 33137 25987 33195 25993
rect 33410 25984 33416 25996
rect 33468 25984 33474 26036
rect 33870 25984 33876 26036
rect 33928 26024 33934 26036
rect 35434 26024 35440 26036
rect 33928 25996 34652 26024
rect 33928 25984 33934 25996
rect 29454 25956 29460 25968
rect 29415 25928 29460 25956
rect 29454 25916 29460 25928
rect 29512 25916 29518 25968
rect 31202 25956 31208 25968
rect 30682 25928 31208 25956
rect 31202 25916 31208 25928
rect 31260 25916 31266 25968
rect 34333 25959 34391 25965
rect 34333 25956 34345 25959
rect 33796 25928 34345 25956
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25888 26295 25891
rect 27522 25888 27528 25900
rect 26283 25860 27528 25888
rect 26283 25857 26295 25860
rect 26237 25851 26295 25857
rect 27522 25848 27528 25860
rect 27580 25848 27586 25900
rect 33594 25888 33600 25900
rect 33555 25860 33600 25888
rect 33594 25848 33600 25860
rect 33652 25848 33658 25900
rect 33796 25897 33824 25928
rect 34333 25925 34345 25928
rect 34379 25925 34391 25959
rect 34333 25919 34391 25925
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25857 33839 25891
rect 33781 25851 33839 25857
rect 34241 25891 34299 25897
rect 34241 25857 34253 25891
rect 34287 25857 34299 25891
rect 34425 25891 34483 25897
rect 34425 25888 34437 25891
rect 34241 25851 34299 25857
rect 34348 25860 34437 25888
rect 26326 25820 26332 25832
rect 26239 25792 26332 25820
rect 26326 25780 26332 25792
rect 26384 25820 26390 25832
rect 27246 25820 27252 25832
rect 26384 25792 27252 25820
rect 26384 25780 26390 25792
rect 27246 25780 27252 25792
rect 27304 25780 27310 25832
rect 29181 25823 29239 25829
rect 29181 25789 29193 25823
rect 29227 25789 29239 25823
rect 29181 25783 29239 25789
rect 28629 25755 28687 25761
rect 28629 25752 28641 25755
rect 27264 25724 28641 25752
rect 27062 25644 27068 25696
rect 27120 25684 27126 25696
rect 27264 25693 27292 25724
rect 28629 25721 28641 25724
rect 28675 25752 28687 25755
rect 29196 25752 29224 25783
rect 33410 25780 33416 25832
rect 33468 25820 33474 25832
rect 34256 25820 34284 25851
rect 33468 25792 34284 25820
rect 33468 25780 33474 25792
rect 28675 25724 29224 25752
rect 28675 25721 28687 25724
rect 28629 25715 28687 25721
rect 34238 25712 34244 25764
rect 34296 25752 34302 25764
rect 34348 25752 34376 25860
rect 34425 25857 34437 25860
rect 34471 25857 34483 25891
rect 34624 25888 34652 25996
rect 35176 25996 35440 26024
rect 35176 25897 35204 25996
rect 35434 25984 35440 25996
rect 35492 25984 35498 26036
rect 35713 26027 35771 26033
rect 35713 25993 35725 26027
rect 35759 26024 35771 26027
rect 36078 26024 36084 26036
rect 35759 25996 36084 26024
rect 35759 25993 35771 25996
rect 35713 25987 35771 25993
rect 36078 25984 36084 25996
rect 36136 25984 36142 26036
rect 38289 26027 38347 26033
rect 38289 25993 38301 26027
rect 38335 26024 38347 26027
rect 39206 26024 39212 26036
rect 38335 25996 39212 26024
rect 38335 25993 38347 25996
rect 38289 25987 38347 25993
rect 39206 25984 39212 25996
rect 39264 25984 39270 26036
rect 41046 26024 41052 26036
rect 41007 25996 41052 26024
rect 41046 25984 41052 25996
rect 41104 25984 41110 26036
rect 35345 25959 35403 25965
rect 35345 25925 35357 25959
rect 35391 25956 35403 25959
rect 36265 25959 36323 25965
rect 36265 25956 36277 25959
rect 35391 25928 36277 25956
rect 35391 25925 35403 25928
rect 35345 25919 35403 25925
rect 36265 25925 36277 25928
rect 36311 25925 36323 25959
rect 42613 25959 42671 25965
rect 42613 25956 42625 25959
rect 36265 25919 36323 25925
rect 36372 25928 42625 25956
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 34624 25860 35173 25888
rect 34425 25851 34483 25857
rect 35161 25857 35173 25860
rect 35207 25857 35219 25891
rect 35434 25888 35440 25900
rect 35395 25860 35440 25888
rect 35161 25851 35219 25857
rect 35176 25820 35204 25851
rect 35434 25848 35440 25860
rect 35492 25848 35498 25900
rect 35526 25848 35532 25900
rect 35584 25888 35590 25900
rect 36372 25897 36400 25928
rect 42613 25925 42625 25928
rect 42659 25956 42671 25959
rect 42794 25956 42800 25968
rect 42659 25928 42800 25956
rect 42659 25925 42671 25928
rect 42613 25919 42671 25925
rect 42794 25916 42800 25928
rect 42852 25916 42858 25968
rect 43622 25916 43628 25968
rect 43680 25956 43686 25968
rect 43680 25928 45402 25956
rect 43680 25916 43686 25928
rect 36173 25891 36231 25897
rect 36173 25888 36185 25891
rect 35584 25860 36185 25888
rect 35584 25848 35590 25860
rect 36173 25857 36185 25860
rect 36219 25857 36231 25891
rect 36173 25851 36231 25857
rect 36357 25891 36415 25897
rect 36357 25857 36369 25891
rect 36403 25857 36415 25891
rect 39482 25888 39488 25900
rect 39443 25860 39488 25888
rect 36357 25851 36415 25857
rect 39482 25848 39488 25860
rect 39540 25848 39546 25900
rect 40126 25888 40132 25900
rect 40087 25860 40132 25888
rect 40126 25848 40132 25860
rect 40184 25848 40190 25900
rect 41141 25891 41199 25897
rect 41141 25857 41153 25891
rect 41187 25888 41199 25891
rect 42058 25888 42064 25900
rect 41187 25860 42064 25888
rect 41187 25857 41199 25860
rect 41141 25851 41199 25857
rect 42058 25848 42064 25860
rect 42116 25848 42122 25900
rect 43438 25888 43444 25900
rect 43399 25860 43444 25888
rect 43438 25848 43444 25860
rect 43496 25848 43502 25900
rect 43530 25848 43536 25900
rect 43588 25888 43594 25900
rect 43588 25860 43633 25888
rect 43588 25848 43594 25860
rect 44818 25848 44824 25900
rect 44876 25888 44882 25900
rect 46017 25891 46075 25897
rect 46017 25888 46029 25891
rect 44876 25860 46029 25888
rect 44876 25848 44882 25860
rect 46017 25857 46029 25860
rect 46063 25857 46075 25891
rect 46017 25851 46075 25857
rect 46106 25848 46112 25900
rect 46164 25888 46170 25900
rect 46477 25891 46535 25897
rect 46477 25888 46489 25891
rect 46164 25860 46489 25888
rect 46164 25848 46170 25860
rect 46477 25857 46489 25860
rect 46523 25857 46535 25891
rect 46477 25851 46535 25857
rect 36817 25823 36875 25829
rect 36817 25820 36829 25823
rect 35176 25792 36829 25820
rect 36817 25789 36829 25792
rect 36863 25789 36875 25823
rect 36817 25783 36875 25789
rect 37829 25823 37887 25829
rect 37829 25789 37841 25823
rect 37875 25820 37887 25823
rect 38010 25820 38016 25832
rect 37875 25792 38016 25820
rect 37875 25789 37887 25792
rect 37829 25783 37887 25789
rect 38010 25780 38016 25792
rect 38068 25780 38074 25832
rect 41233 25823 41291 25829
rect 41233 25789 41245 25823
rect 41279 25789 41291 25823
rect 41233 25783 41291 25789
rect 34296 25724 34376 25752
rect 38197 25755 38255 25761
rect 34296 25712 34302 25724
rect 38197 25721 38209 25755
rect 38243 25752 38255 25755
rect 38378 25752 38384 25764
rect 38243 25724 38384 25752
rect 38243 25721 38255 25724
rect 38197 25715 38255 25721
rect 38378 25712 38384 25724
rect 38436 25712 38442 25764
rect 41138 25712 41144 25764
rect 41196 25752 41202 25764
rect 41248 25752 41276 25783
rect 41196 25724 41276 25752
rect 41196 25712 41202 25724
rect 27249 25687 27307 25693
rect 27249 25684 27261 25687
rect 27120 25656 27261 25684
rect 27120 25644 27126 25656
rect 27249 25653 27261 25656
rect 27295 25653 27307 25687
rect 27249 25647 27307 25653
rect 27522 25644 27528 25696
rect 27580 25684 27586 25696
rect 27893 25687 27951 25693
rect 27893 25684 27905 25687
rect 27580 25656 27905 25684
rect 27580 25644 27586 25656
rect 27893 25653 27905 25656
rect 27939 25684 27951 25687
rect 30650 25684 30656 25696
rect 27939 25656 30656 25684
rect 27939 25653 27951 25656
rect 27893 25647 27951 25653
rect 30650 25644 30656 25656
rect 30708 25644 30714 25696
rect 30926 25684 30932 25696
rect 30887 25656 30932 25684
rect 30926 25644 30932 25656
rect 30984 25644 30990 25696
rect 33134 25644 33140 25696
rect 33192 25684 33198 25696
rect 33597 25687 33655 25693
rect 33597 25684 33609 25687
rect 33192 25656 33609 25684
rect 33192 25644 33198 25656
rect 33597 25653 33609 25656
rect 33643 25653 33655 25687
rect 33597 25647 33655 25653
rect 39853 25687 39911 25693
rect 39853 25653 39865 25687
rect 39899 25684 39911 25687
rect 39942 25684 39948 25696
rect 39899 25656 39948 25684
rect 39899 25653 39911 25656
rect 39853 25647 39911 25653
rect 39942 25644 39948 25656
rect 40000 25644 40006 25696
rect 40681 25687 40739 25693
rect 40681 25653 40693 25687
rect 40727 25684 40739 25687
rect 41046 25684 41052 25696
rect 40727 25656 41052 25684
rect 40727 25653 40739 25656
rect 40681 25647 40739 25653
rect 41046 25644 41052 25656
rect 41104 25644 41110 25696
rect 41966 25684 41972 25696
rect 41879 25656 41972 25684
rect 41966 25644 41972 25656
rect 42024 25684 42030 25696
rect 43346 25684 43352 25696
rect 42024 25656 43352 25684
rect 42024 25644 42030 25656
rect 43346 25644 43352 25656
rect 43404 25644 43410 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 27522 25480 27528 25492
rect 27483 25452 27528 25480
rect 27522 25440 27528 25452
rect 27580 25440 27586 25492
rect 33594 25440 33600 25492
rect 33652 25480 33658 25492
rect 33870 25480 33876 25492
rect 33652 25452 33876 25480
rect 33652 25440 33658 25452
rect 33870 25440 33876 25452
rect 33928 25440 33934 25492
rect 34057 25483 34115 25489
rect 34057 25449 34069 25483
rect 34103 25449 34115 25483
rect 34057 25443 34115 25449
rect 35253 25483 35311 25489
rect 35253 25449 35265 25483
rect 35299 25480 35311 25483
rect 35802 25480 35808 25492
rect 35299 25452 35808 25480
rect 35299 25449 35311 25452
rect 35253 25443 35311 25449
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 27540 25276 27568 25440
rect 30926 25412 30932 25424
rect 30887 25384 30932 25412
rect 30926 25372 30932 25384
rect 30984 25372 30990 25424
rect 33962 25412 33968 25424
rect 33428 25384 33968 25412
rect 33134 25344 33140 25356
rect 33095 25316 33140 25344
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 33428 25288 33456 25384
rect 33962 25372 33968 25384
rect 34020 25412 34026 25424
rect 34072 25412 34100 25443
rect 35802 25440 35808 25452
rect 35860 25440 35866 25492
rect 39206 25440 39212 25492
rect 39264 25480 39270 25492
rect 39301 25483 39359 25489
rect 39301 25480 39313 25483
rect 39264 25452 39313 25480
rect 39264 25440 39270 25452
rect 39301 25449 39313 25452
rect 39347 25480 39359 25483
rect 40037 25483 40095 25489
rect 40037 25480 40049 25483
rect 39347 25452 40049 25480
rect 39347 25449 39359 25452
rect 39301 25443 39359 25449
rect 40037 25449 40049 25452
rect 40083 25449 40095 25483
rect 41046 25480 41052 25492
rect 41007 25452 41052 25480
rect 40037 25443 40095 25449
rect 41046 25440 41052 25452
rect 41104 25440 41110 25492
rect 35526 25412 35532 25424
rect 34020 25384 34100 25412
rect 35084 25384 35532 25412
rect 34020 25372 34026 25384
rect 30466 25276 30472 25288
rect 26927 25248 27568 25276
rect 30427 25248 30472 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 30466 25236 30472 25248
rect 30524 25236 30530 25288
rect 33410 25236 33416 25288
rect 33468 25276 33474 25288
rect 35084 25285 35112 25384
rect 35526 25372 35532 25384
rect 35584 25372 35590 25424
rect 38010 25372 38016 25424
rect 38068 25412 38074 25424
rect 39117 25415 39175 25421
rect 39117 25412 39129 25415
rect 38068 25384 39129 25412
rect 38068 25372 38074 25384
rect 39117 25381 39129 25384
rect 39163 25412 39175 25415
rect 41138 25412 41144 25424
rect 39163 25384 41144 25412
rect 39163 25381 39175 25384
rect 39117 25375 39175 25381
rect 41138 25372 41144 25384
rect 41196 25372 41202 25424
rect 41693 25415 41751 25421
rect 41693 25412 41705 25415
rect 41386 25384 41705 25412
rect 35434 25304 35440 25356
rect 35492 25344 35498 25356
rect 38105 25347 38163 25353
rect 38105 25344 38117 25347
rect 35492 25316 38117 25344
rect 35492 25304 35498 25316
rect 38105 25313 38117 25316
rect 38151 25313 38163 25347
rect 38105 25307 38163 25313
rect 39298 25304 39304 25356
rect 39356 25344 39362 25356
rect 40865 25347 40923 25353
rect 40865 25344 40877 25347
rect 39356 25316 40877 25344
rect 39356 25304 39362 25316
rect 40865 25313 40877 25316
rect 40911 25313 40923 25347
rect 41386 25344 41414 25384
rect 41693 25381 41705 25384
rect 41739 25412 41751 25415
rect 43990 25412 43996 25424
rect 41739 25384 43996 25412
rect 41739 25381 41751 25384
rect 41693 25375 41751 25381
rect 43990 25372 43996 25384
rect 44048 25372 44054 25424
rect 40865 25307 40923 25313
rect 40972 25316 41414 25344
rect 42337 25347 42395 25353
rect 35069 25279 35127 25285
rect 33468 25248 33513 25276
rect 33888 25248 34365 25276
rect 33468 25236 33474 25248
rect 26973 25211 27031 25217
rect 26973 25177 26985 25211
rect 27019 25208 27031 25211
rect 27062 25208 27068 25220
rect 27019 25180 27068 25208
rect 27019 25177 27031 25180
rect 26973 25171 27031 25177
rect 27062 25168 27068 25180
rect 27120 25168 27126 25220
rect 31386 25208 31392 25220
rect 31347 25180 31392 25208
rect 31386 25168 31392 25180
rect 31444 25168 31450 25220
rect 32674 25168 32680 25220
rect 32732 25208 32738 25220
rect 33888 25208 33916 25248
rect 34054 25217 34060 25220
rect 32732 25180 33916 25208
rect 34041 25211 34060 25217
rect 32732 25168 32738 25180
rect 34041 25177 34053 25211
rect 34041 25171 34060 25177
rect 34054 25168 34060 25171
rect 34112 25168 34118 25220
rect 34238 25208 34244 25220
rect 34199 25180 34244 25208
rect 34238 25168 34244 25180
rect 34296 25168 34302 25220
rect 34337 25208 34365 25248
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35250 25276 35256 25288
rect 35211 25248 35256 25276
rect 35069 25239 35127 25245
rect 35250 25236 35256 25248
rect 35308 25236 35314 25288
rect 35894 25276 35900 25288
rect 35855 25248 35900 25276
rect 35894 25236 35900 25248
rect 35952 25236 35958 25288
rect 37274 25236 37280 25288
rect 37332 25236 37338 25288
rect 40034 25276 40040 25288
rect 39995 25248 40040 25276
rect 40034 25236 40040 25248
rect 40092 25236 40098 25288
rect 40218 25236 40224 25288
rect 40276 25276 40282 25288
rect 40770 25276 40776 25288
rect 40276 25248 40776 25276
rect 40276 25236 40282 25248
rect 40770 25236 40776 25248
rect 40828 25236 40834 25288
rect 34337 25180 35664 25208
rect 28350 25100 28356 25152
rect 28408 25140 28414 25152
rect 30469 25143 30527 25149
rect 30469 25140 30481 25143
rect 28408 25112 30481 25140
rect 28408 25100 28414 25112
rect 30469 25109 30481 25112
rect 30515 25109 30527 25143
rect 30469 25103 30527 25109
rect 35437 25143 35495 25149
rect 35437 25109 35449 25143
rect 35483 25140 35495 25143
rect 35526 25140 35532 25152
rect 35483 25112 35532 25140
rect 35483 25109 35495 25112
rect 35437 25103 35495 25109
rect 35526 25100 35532 25112
rect 35584 25100 35590 25152
rect 35636 25140 35664 25180
rect 35710 25168 35716 25220
rect 35768 25208 35774 25220
rect 36173 25211 36231 25217
rect 36173 25208 36185 25211
rect 35768 25180 36185 25208
rect 35768 25168 35774 25180
rect 36173 25177 36185 25180
rect 36219 25177 36231 25211
rect 36173 25171 36231 25177
rect 37292 25140 37320 25236
rect 38838 25208 38844 25220
rect 38799 25180 38844 25208
rect 38838 25168 38844 25180
rect 38896 25168 38902 25220
rect 40126 25168 40132 25220
rect 40184 25208 40190 25220
rect 40972 25208 41000 25316
rect 42337 25313 42349 25347
rect 42383 25344 42395 25347
rect 43438 25344 43444 25356
rect 42383 25316 43444 25344
rect 42383 25313 42395 25316
rect 42337 25307 42395 25313
rect 43438 25304 43444 25316
rect 43496 25304 43502 25356
rect 41141 25279 41199 25285
rect 41141 25245 41153 25279
rect 41187 25276 41199 25279
rect 41230 25276 41236 25288
rect 41187 25248 41236 25276
rect 41187 25245 41199 25248
rect 41141 25239 41199 25245
rect 41230 25236 41236 25248
rect 41288 25276 41294 25288
rect 41966 25276 41972 25288
rect 41288 25248 41972 25276
rect 41288 25236 41294 25248
rect 41966 25236 41972 25248
rect 42024 25236 42030 25288
rect 42426 25276 42432 25288
rect 42387 25248 42432 25276
rect 42426 25236 42432 25248
rect 42484 25236 42490 25288
rect 43346 25276 43352 25288
rect 43259 25248 43352 25276
rect 43346 25236 43352 25248
rect 43404 25276 43410 25288
rect 43898 25276 43904 25288
rect 43404 25248 43904 25276
rect 43404 25236 43410 25248
rect 43898 25236 43904 25248
rect 43956 25236 43962 25288
rect 45189 25279 45247 25285
rect 45189 25245 45201 25279
rect 45235 25276 45247 25279
rect 46106 25276 46112 25288
rect 45235 25248 46112 25276
rect 45235 25245 45247 25248
rect 45189 25239 45247 25245
rect 46106 25236 46112 25248
rect 46164 25236 46170 25288
rect 40184 25180 41000 25208
rect 42797 25211 42855 25217
rect 40184 25168 40190 25180
rect 42797 25177 42809 25211
rect 42843 25208 42855 25211
rect 42978 25208 42984 25220
rect 42843 25180 42984 25208
rect 42843 25177 42855 25180
rect 42797 25171 42855 25177
rect 42978 25168 42984 25180
rect 43036 25208 43042 25220
rect 43806 25208 43812 25220
rect 43036 25180 43812 25208
rect 43036 25168 43042 25180
rect 43806 25168 43812 25180
rect 43864 25208 43870 25220
rect 44085 25211 44143 25217
rect 44085 25208 44097 25211
rect 43864 25180 44097 25208
rect 43864 25168 43870 25180
rect 44085 25177 44097 25180
rect 44131 25177 44143 25211
rect 45462 25208 45468 25220
rect 45423 25180 45468 25208
rect 44085 25171 44143 25177
rect 45462 25168 45468 25180
rect 45520 25168 45526 25220
rect 37642 25140 37648 25152
rect 35636 25112 37320 25140
rect 37603 25112 37648 25140
rect 37642 25100 37648 25112
rect 37700 25100 37706 25152
rect 38102 25100 38108 25152
rect 38160 25140 38166 25152
rect 39206 25140 39212 25152
rect 38160 25112 39212 25140
rect 38160 25100 38166 25112
rect 39206 25100 39212 25112
rect 39264 25100 39270 25152
rect 40310 25100 40316 25152
rect 40368 25140 40374 25152
rect 40405 25143 40463 25149
rect 40405 25140 40417 25143
rect 40368 25112 40417 25140
rect 40368 25100 40374 25112
rect 40405 25109 40417 25112
rect 40451 25109 40463 25143
rect 40862 25140 40868 25152
rect 40823 25112 40868 25140
rect 40405 25103 40463 25109
rect 40862 25100 40868 25112
rect 40920 25100 40926 25152
rect 42150 25140 42156 25152
rect 42111 25112 42156 25140
rect 42150 25100 42156 25112
rect 42208 25100 42214 25152
rect 43346 25100 43352 25152
rect 43404 25140 43410 25152
rect 44177 25143 44235 25149
rect 44177 25140 44189 25143
rect 43404 25112 44189 25140
rect 43404 25100 43410 25112
rect 44177 25109 44189 25112
rect 44223 25109 44235 25143
rect 44177 25103 44235 25109
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 30466 24896 30472 24948
rect 30524 24936 30530 24948
rect 31021 24939 31079 24945
rect 31021 24936 31033 24939
rect 30524 24908 31033 24936
rect 30524 24896 30530 24908
rect 31021 24905 31033 24908
rect 31067 24905 31079 24939
rect 31021 24899 31079 24905
rect 32861 24939 32919 24945
rect 32861 24905 32873 24939
rect 32907 24936 32919 24939
rect 34054 24936 34060 24948
rect 32907 24908 34060 24936
rect 32907 24905 32919 24908
rect 32861 24899 32919 24905
rect 34054 24896 34060 24908
rect 34112 24896 34118 24948
rect 35250 24896 35256 24948
rect 35308 24936 35314 24948
rect 35986 24936 35992 24948
rect 35308 24908 35992 24936
rect 35308 24896 35314 24908
rect 35986 24896 35992 24908
rect 36044 24936 36050 24948
rect 40494 24936 40500 24948
rect 36044 24908 40500 24936
rect 36044 24896 36050 24908
rect 40494 24896 40500 24908
rect 40552 24936 40558 24948
rect 41046 24936 41052 24948
rect 40552 24908 40908 24936
rect 41007 24908 41052 24936
rect 40552 24896 40558 24908
rect 33962 24828 33968 24880
rect 34020 24868 34026 24880
rect 34020 24840 34284 24868
rect 34020 24828 34026 24840
rect 24946 24760 24952 24812
rect 25004 24760 25010 24812
rect 31757 24803 31815 24809
rect 31757 24769 31769 24803
rect 31803 24800 31815 24803
rect 33318 24800 33324 24812
rect 31803 24772 33324 24800
rect 31803 24769 31815 24772
rect 31757 24763 31815 24769
rect 33318 24760 33324 24772
rect 33376 24760 33382 24812
rect 34256 24809 34284 24840
rect 37642 24828 37648 24880
rect 37700 24868 37706 24880
rect 38746 24868 38752 24880
rect 37700 24840 38752 24868
rect 37700 24828 37706 24840
rect 38746 24828 38752 24840
rect 38804 24868 38810 24880
rect 40586 24868 40592 24880
rect 38804 24840 40592 24868
rect 38804 24828 38810 24840
rect 40586 24828 40592 24840
rect 40644 24828 40650 24880
rect 40880 24868 40908 24908
rect 41046 24896 41052 24908
rect 41104 24896 41110 24948
rect 41141 24939 41199 24945
rect 41141 24905 41153 24939
rect 41187 24936 41199 24939
rect 41690 24936 41696 24948
rect 41187 24908 41696 24936
rect 41187 24905 41199 24908
rect 41141 24899 41199 24905
rect 41690 24896 41696 24908
rect 41748 24936 41754 24948
rect 42150 24936 42156 24948
rect 41748 24908 42156 24936
rect 41748 24896 41754 24908
rect 42150 24896 42156 24908
rect 42208 24896 42214 24948
rect 42978 24945 42984 24948
rect 42797 24939 42855 24945
rect 42797 24936 42809 24939
rect 42260 24908 42809 24936
rect 42260 24868 42288 24908
rect 42797 24905 42809 24908
rect 42843 24905 42855 24939
rect 42797 24899 42855 24905
rect 42965 24939 42984 24945
rect 42965 24905 42977 24939
rect 42965 24899 42984 24905
rect 42978 24896 42984 24899
rect 43036 24896 43042 24948
rect 40880 24840 42288 24868
rect 42426 24828 42432 24880
rect 42484 24868 42490 24880
rect 43165 24871 43223 24877
rect 43165 24868 43177 24871
rect 42484 24840 43177 24868
rect 42484 24828 42490 24840
rect 43165 24837 43177 24840
rect 43211 24868 43223 24871
rect 43530 24868 43536 24880
rect 43211 24840 43536 24868
rect 43211 24837 43223 24840
rect 43165 24831 43223 24837
rect 43530 24828 43536 24840
rect 43588 24868 43594 24880
rect 45462 24868 45468 24880
rect 43588 24840 45468 24868
rect 43588 24828 43594 24840
rect 34149 24803 34207 24809
rect 34149 24800 34161 24803
rect 34072 24772 34161 24800
rect 2038 24692 2044 24744
rect 2096 24732 2102 24744
rect 24213 24735 24271 24741
rect 24213 24732 24225 24735
rect 2096 24704 24225 24732
rect 2096 24692 2102 24704
rect 24213 24701 24225 24704
rect 24259 24701 24271 24735
rect 25038 24732 25044 24744
rect 24999 24704 25044 24732
rect 24213 24695 24271 24701
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 33336 24664 33364 24760
rect 33870 24732 33876 24744
rect 33831 24704 33876 24732
rect 33870 24692 33876 24704
rect 33928 24692 33934 24744
rect 34072 24732 34100 24772
rect 34149 24769 34161 24772
rect 34195 24769 34207 24803
rect 34149 24763 34207 24769
rect 34241 24803 34299 24809
rect 34241 24769 34253 24803
rect 34287 24769 34299 24803
rect 34241 24763 34299 24769
rect 34330 24760 34336 24812
rect 34388 24800 34394 24812
rect 34388 24772 34433 24800
rect 34388 24760 34394 24772
rect 34514 24760 34520 24812
rect 34572 24800 34578 24812
rect 34572 24772 34617 24800
rect 34572 24760 34578 24772
rect 34790 24760 34796 24812
rect 34848 24800 34854 24812
rect 35805 24803 35863 24809
rect 34848 24772 35756 24800
rect 34848 24760 34854 24772
rect 35342 24732 35348 24744
rect 34072 24704 35348 24732
rect 35342 24692 35348 24704
rect 35400 24692 35406 24744
rect 35526 24732 35532 24744
rect 35487 24704 35532 24732
rect 35526 24692 35532 24704
rect 35584 24692 35590 24744
rect 35728 24732 35756 24772
rect 35805 24769 35817 24803
rect 35851 24800 35863 24803
rect 35894 24800 35900 24812
rect 35851 24772 35900 24800
rect 35851 24769 35863 24772
rect 35805 24763 35863 24769
rect 35894 24760 35900 24772
rect 35952 24760 35958 24812
rect 36449 24803 36507 24809
rect 36449 24769 36461 24803
rect 36495 24800 36507 24803
rect 36538 24800 36544 24812
rect 36495 24772 36544 24800
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 36814 24760 36820 24812
rect 36872 24800 36878 24812
rect 37918 24800 37924 24812
rect 36872 24772 37924 24800
rect 36872 24760 36878 24772
rect 37918 24760 37924 24772
rect 37976 24760 37982 24812
rect 38010 24760 38016 24812
rect 38068 24800 38074 24812
rect 38105 24803 38163 24809
rect 38105 24800 38117 24803
rect 38068 24772 38117 24800
rect 38068 24760 38074 24772
rect 38105 24769 38117 24772
rect 38151 24769 38163 24803
rect 38562 24800 38568 24812
rect 38523 24772 38568 24800
rect 38105 24763 38163 24769
rect 38562 24760 38568 24772
rect 38620 24760 38626 24812
rect 38838 24760 38844 24812
rect 38896 24800 38902 24812
rect 39209 24803 39267 24809
rect 39209 24800 39221 24803
rect 38896 24772 39221 24800
rect 38896 24760 38902 24772
rect 39209 24769 39221 24772
rect 39255 24800 39267 24803
rect 39666 24800 39672 24812
rect 39255 24772 39672 24800
rect 39255 24769 39267 24772
rect 39209 24763 39267 24769
rect 39666 24760 39672 24772
rect 39724 24760 39730 24812
rect 39761 24803 39819 24809
rect 39761 24769 39773 24803
rect 39807 24800 39819 24803
rect 40954 24800 40960 24812
rect 39807 24772 40816 24800
rect 40915 24772 40960 24800
rect 39807 24769 39819 24772
rect 39761 24763 39819 24769
rect 38473 24735 38531 24741
rect 35728 24704 38424 24732
rect 35618 24664 35624 24676
rect 33336 24636 35112 24664
rect 35579 24636 35624 24664
rect 28261 24599 28319 24605
rect 28261 24565 28273 24599
rect 28307 24596 28319 24599
rect 28442 24596 28448 24608
rect 28307 24568 28448 24596
rect 28307 24565 28319 24568
rect 28261 24559 28319 24565
rect 28442 24556 28448 24568
rect 28500 24556 28506 24608
rect 33413 24599 33471 24605
rect 33413 24565 33425 24599
rect 33459 24596 33471 24599
rect 33594 24596 33600 24608
rect 33459 24568 33600 24596
rect 33459 24565 33471 24568
rect 33413 24559 33471 24565
rect 33594 24556 33600 24568
rect 33652 24596 33658 24608
rect 34238 24596 34244 24608
rect 33652 24568 34244 24596
rect 33652 24556 33658 24568
rect 34238 24556 34244 24568
rect 34296 24596 34302 24608
rect 34977 24599 35035 24605
rect 34977 24596 34989 24599
rect 34296 24568 34989 24596
rect 34296 24556 34302 24568
rect 34977 24565 34989 24568
rect 35023 24565 35035 24599
rect 35084 24596 35112 24636
rect 35618 24624 35624 24636
rect 35676 24624 35682 24676
rect 36814 24664 36820 24676
rect 36775 24636 36820 24664
rect 36814 24624 36820 24636
rect 36872 24624 36878 24676
rect 35713 24599 35771 24605
rect 35713 24596 35725 24599
rect 35084 24568 35725 24596
rect 34977 24559 35035 24565
rect 35713 24565 35725 24568
rect 35759 24565 35771 24599
rect 35713 24559 35771 24565
rect 36909 24599 36967 24605
rect 36909 24565 36921 24599
rect 36955 24596 36967 24599
rect 37274 24596 37280 24608
rect 36955 24568 37280 24596
rect 36955 24565 36967 24568
rect 36909 24559 36967 24565
rect 37274 24556 37280 24568
rect 37332 24556 37338 24608
rect 38396 24596 38424 24704
rect 38473 24701 38485 24735
rect 38519 24732 38531 24735
rect 38746 24732 38752 24744
rect 38519 24704 38752 24732
rect 38519 24701 38531 24704
rect 38473 24695 38531 24701
rect 38746 24692 38752 24704
rect 38804 24692 38810 24744
rect 40788 24732 40816 24772
rect 40954 24760 40960 24772
rect 41012 24760 41018 24812
rect 41325 24803 41383 24809
rect 41325 24769 41337 24803
rect 41371 24800 41383 24803
rect 41598 24800 41604 24812
rect 41371 24772 41604 24800
rect 41371 24769 41383 24772
rect 41325 24763 41383 24769
rect 41598 24760 41604 24772
rect 41656 24800 41662 24812
rect 43622 24800 43628 24812
rect 41656 24772 43628 24800
rect 41656 24760 41662 24772
rect 43622 24760 43628 24772
rect 43680 24760 43686 24812
rect 43809 24803 43867 24809
rect 43809 24769 43821 24803
rect 43855 24800 43867 24803
rect 44266 24800 44272 24812
rect 43855 24772 44272 24800
rect 43855 24769 43867 24772
rect 43809 24763 43867 24769
rect 44266 24760 44272 24772
rect 44324 24760 44330 24812
rect 44818 24800 44824 24812
rect 44779 24772 44824 24800
rect 44818 24760 44824 24772
rect 44876 24760 44882 24812
rect 44928 24809 44956 24840
rect 45462 24828 45468 24840
rect 45520 24828 45526 24880
rect 44913 24803 44971 24809
rect 44913 24769 44925 24803
rect 44959 24769 44971 24803
rect 44913 24763 44971 24769
rect 45280 24803 45338 24809
rect 45280 24769 45292 24803
rect 45326 24800 45338 24803
rect 45554 24800 45560 24812
rect 45326 24772 45560 24800
rect 45326 24769 45338 24772
rect 45280 24763 45338 24769
rect 45554 24760 45560 24772
rect 45612 24800 45618 24812
rect 45925 24803 45983 24809
rect 45925 24800 45937 24803
rect 45612 24772 45937 24800
rect 45612 24760 45618 24772
rect 45925 24769 45937 24772
rect 45971 24769 45983 24803
rect 45925 24763 45983 24769
rect 41230 24732 41236 24744
rect 40788 24704 41236 24732
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 41417 24735 41475 24741
rect 41417 24701 41429 24735
rect 41463 24732 41475 24735
rect 41506 24732 41512 24744
rect 41463 24704 41512 24732
rect 41463 24701 41475 24704
rect 41417 24695 41475 24701
rect 41506 24692 41512 24704
rect 41564 24692 41570 24744
rect 38562 24624 38568 24676
rect 38620 24664 38626 24676
rect 41877 24667 41935 24673
rect 41877 24664 41889 24667
rect 38620 24636 41889 24664
rect 38620 24624 38626 24636
rect 41877 24633 41889 24636
rect 41923 24664 41935 24667
rect 42610 24664 42616 24676
rect 41923 24636 42616 24664
rect 41923 24633 41935 24636
rect 41877 24627 41935 24633
rect 42610 24624 42616 24636
rect 42668 24624 42674 24676
rect 43438 24664 43444 24676
rect 42996 24636 43444 24664
rect 39206 24596 39212 24608
rect 38396 24568 39212 24596
rect 39206 24556 39212 24568
rect 39264 24556 39270 24608
rect 40037 24599 40095 24605
rect 40037 24565 40049 24599
rect 40083 24596 40095 24599
rect 40218 24596 40224 24608
rect 40083 24568 40224 24596
rect 40083 24565 40095 24568
rect 40037 24559 40095 24565
rect 40218 24556 40224 24568
rect 40276 24556 40282 24608
rect 40678 24596 40684 24608
rect 40639 24568 40684 24596
rect 40678 24556 40684 24568
rect 40736 24556 40742 24608
rect 42996 24605 43024 24636
rect 43438 24624 43444 24636
rect 43496 24664 43502 24676
rect 44082 24664 44088 24676
rect 43496 24636 44088 24664
rect 43496 24624 43502 24636
rect 44082 24624 44088 24636
rect 44140 24624 44146 24676
rect 45462 24664 45468 24676
rect 45423 24636 45468 24664
rect 45462 24624 45468 24636
rect 45520 24624 45526 24676
rect 42981 24599 43039 24605
rect 42981 24565 42993 24599
rect 43027 24565 43039 24599
rect 42981 24559 43039 24565
rect 43806 24556 43812 24608
rect 43864 24596 43870 24608
rect 43901 24599 43959 24605
rect 43901 24596 43913 24599
rect 43864 24568 43913 24596
rect 43864 24556 43870 24568
rect 43901 24565 43913 24568
rect 43947 24565 43959 24599
rect 43901 24559 43959 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 34149 24395 34207 24401
rect 34149 24361 34161 24395
rect 34195 24392 34207 24395
rect 34330 24392 34336 24404
rect 34195 24364 34336 24392
rect 34195 24361 34207 24364
rect 34149 24355 34207 24361
rect 34330 24352 34336 24364
rect 34388 24352 34394 24404
rect 35713 24395 35771 24401
rect 35713 24361 35725 24395
rect 35759 24392 35771 24395
rect 37826 24392 37832 24404
rect 35759 24364 37832 24392
rect 35759 24361 35771 24364
rect 35713 24355 35771 24361
rect 37826 24352 37832 24364
rect 37884 24352 37890 24404
rect 37918 24352 37924 24404
rect 37976 24392 37982 24404
rect 39393 24395 39451 24401
rect 39393 24392 39405 24395
rect 37976 24364 39405 24392
rect 37976 24352 37982 24364
rect 39393 24361 39405 24364
rect 39439 24392 39451 24395
rect 40126 24392 40132 24404
rect 39439 24364 40132 24392
rect 39439 24361 39451 24364
rect 39393 24355 39451 24361
rect 40126 24352 40132 24364
rect 40184 24352 40190 24404
rect 40678 24392 40684 24404
rect 40639 24364 40684 24392
rect 40678 24352 40684 24364
rect 40736 24352 40742 24404
rect 42242 24392 42248 24404
rect 40880 24364 42248 24392
rect 34514 24284 34520 24336
rect 34572 24324 34578 24336
rect 38473 24327 38531 24333
rect 38473 24324 38485 24327
rect 34572 24296 38485 24324
rect 34572 24284 34578 24296
rect 38473 24293 38485 24296
rect 38519 24293 38531 24327
rect 38746 24324 38752 24336
rect 38473 24287 38531 24293
rect 38626 24296 38752 24324
rect 28905 24259 28963 24265
rect 28905 24225 28917 24259
rect 28951 24256 28963 24259
rect 28994 24256 29000 24268
rect 28951 24228 29000 24256
rect 28951 24225 28963 24228
rect 28905 24219 28963 24225
rect 28994 24216 29000 24228
rect 29052 24216 29058 24268
rect 29181 24259 29239 24265
rect 29181 24225 29193 24259
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 30561 24259 30619 24265
rect 30561 24225 30573 24259
rect 30607 24256 30619 24259
rect 30742 24256 30748 24268
rect 30607 24228 30748 24256
rect 30607 24225 30619 24228
rect 30561 24219 30619 24225
rect 25958 24188 25964 24200
rect 25919 24160 25964 24188
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26418 24148 26424 24200
rect 26476 24188 26482 24200
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 26476 24160 26617 24188
rect 26476 24148 26482 24160
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24188 28135 24191
rect 28258 24188 28264 24200
rect 28123 24160 28264 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 27430 24120 27436 24132
rect 27391 24092 27436 24120
rect 27430 24080 27436 24092
rect 27488 24080 27494 24132
rect 27908 24120 27936 24151
rect 28258 24148 28264 24160
rect 28316 24148 28322 24200
rect 28813 24191 28871 24197
rect 28813 24157 28825 24191
rect 28859 24188 28871 24191
rect 29086 24188 29092 24200
rect 28859 24160 29092 24188
rect 28859 24157 28871 24160
rect 28813 24151 28871 24157
rect 29086 24148 29092 24160
rect 29144 24148 29150 24200
rect 29196 24188 29224 24219
rect 30742 24216 30748 24228
rect 30800 24216 30806 24268
rect 33045 24259 33103 24265
rect 33045 24225 33057 24259
rect 33091 24256 33103 24259
rect 33870 24256 33876 24268
rect 33091 24228 33876 24256
rect 33091 24225 33103 24228
rect 33045 24219 33103 24225
rect 33870 24216 33876 24228
rect 33928 24216 33934 24268
rect 33962 24216 33968 24268
rect 34020 24256 34026 24268
rect 38626 24256 38654 24296
rect 38746 24284 38752 24296
rect 38804 24284 38810 24336
rect 40034 24284 40040 24336
rect 40092 24324 40098 24336
rect 40880 24324 40908 24364
rect 42242 24352 42248 24364
rect 42300 24392 42306 24404
rect 42300 24364 43024 24392
rect 42300 24352 42306 24364
rect 40092 24296 40908 24324
rect 40092 24284 40098 24296
rect 41138 24284 41144 24336
rect 41196 24324 41202 24336
rect 42797 24327 42855 24333
rect 42797 24324 42809 24327
rect 41196 24296 42809 24324
rect 41196 24284 41202 24296
rect 42797 24293 42809 24296
rect 42843 24293 42855 24327
rect 42996 24324 43024 24364
rect 43990 24352 43996 24404
rect 44048 24392 44054 24404
rect 44453 24395 44511 24401
rect 44453 24392 44465 24395
rect 44048 24364 44465 24392
rect 44048 24352 44054 24364
rect 44453 24361 44465 24364
rect 44499 24361 44511 24395
rect 44453 24355 44511 24361
rect 45462 24324 45468 24336
rect 42996 24296 45468 24324
rect 42797 24287 42855 24293
rect 40773 24259 40831 24265
rect 34020 24228 34284 24256
rect 34020 24216 34026 24228
rect 30098 24188 30104 24200
rect 29196 24160 30104 24188
rect 30098 24148 30104 24160
rect 30156 24188 30162 24200
rect 30469 24191 30527 24197
rect 30469 24188 30481 24191
rect 30156 24160 30481 24188
rect 30156 24148 30162 24160
rect 30469 24157 30481 24160
rect 30515 24157 30527 24191
rect 30469 24151 30527 24157
rect 31297 24191 31355 24197
rect 31297 24157 31309 24191
rect 31343 24188 31355 24191
rect 31662 24188 31668 24200
rect 31343 24160 31668 24188
rect 31343 24157 31355 24160
rect 31297 24151 31355 24157
rect 31662 24148 31668 24160
rect 31720 24148 31726 24200
rect 33321 24191 33379 24197
rect 33321 24157 33333 24191
rect 33367 24188 33379 24191
rect 33410 24188 33416 24200
rect 33367 24160 33416 24188
rect 33367 24157 33379 24160
rect 33321 24151 33379 24157
rect 33410 24148 33416 24160
rect 33468 24148 33474 24200
rect 33686 24148 33692 24200
rect 33744 24188 33750 24200
rect 34256 24197 34284 24228
rect 36924 24228 38654 24256
rect 38856 24228 40540 24256
rect 34057 24191 34115 24197
rect 34057 24188 34069 24191
rect 33744 24160 34069 24188
rect 33744 24148 33750 24160
rect 34057 24157 34069 24160
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34241 24191 34299 24197
rect 34241 24157 34253 24191
rect 34287 24157 34299 24191
rect 34241 24151 34299 24157
rect 35434 24148 35440 24200
rect 35492 24188 35498 24200
rect 35529 24191 35587 24197
rect 35529 24188 35541 24191
rect 35492 24160 35541 24188
rect 35492 24148 35498 24160
rect 35529 24157 35541 24160
rect 35575 24157 35587 24191
rect 35529 24151 35587 24157
rect 35805 24191 35863 24197
rect 35805 24157 35817 24191
rect 35851 24188 35863 24191
rect 35894 24188 35900 24200
rect 35851 24160 35900 24188
rect 35851 24157 35863 24160
rect 35805 24151 35863 24157
rect 35894 24148 35900 24160
rect 35952 24188 35958 24200
rect 36538 24188 36544 24200
rect 35952 24160 36544 24188
rect 35952 24148 35958 24160
rect 36538 24148 36544 24160
rect 36596 24148 36602 24200
rect 36725 24191 36783 24197
rect 36725 24157 36737 24191
rect 36771 24188 36783 24191
rect 36814 24188 36820 24200
rect 36771 24160 36820 24188
rect 36771 24157 36783 24160
rect 36725 24151 36783 24157
rect 36814 24148 36820 24160
rect 36872 24148 36878 24200
rect 36924 24197 36952 24228
rect 36909 24191 36967 24197
rect 36909 24157 36921 24191
rect 36955 24157 36967 24191
rect 36909 24151 36967 24157
rect 37093 24191 37151 24197
rect 37093 24157 37105 24191
rect 37139 24157 37151 24191
rect 37274 24188 37280 24200
rect 37235 24160 37280 24188
rect 37093 24151 37151 24157
rect 28442 24120 28448 24132
rect 27908 24092 28448 24120
rect 28442 24080 28448 24092
rect 28500 24080 28506 24132
rect 32582 24080 32588 24132
rect 32640 24080 32646 24132
rect 37001 24123 37059 24129
rect 37001 24120 37013 24123
rect 32692 24092 37013 24120
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 27893 24055 27951 24061
rect 27893 24052 27905 24055
rect 27856 24024 27905 24052
rect 27856 24012 27862 24024
rect 27893 24021 27905 24024
rect 27939 24021 27951 24055
rect 27893 24015 27951 24021
rect 27982 24012 27988 24064
rect 28040 24052 28046 24064
rect 30101 24055 30159 24061
rect 30101 24052 30113 24055
rect 28040 24024 30113 24052
rect 28040 24012 28046 24024
rect 30101 24021 30113 24024
rect 30147 24021 30159 24055
rect 30101 24015 30159 24021
rect 32214 24012 32220 24064
rect 32272 24052 32278 24064
rect 32692 24052 32720 24092
rect 37001 24089 37013 24092
rect 37047 24089 37059 24123
rect 37108 24120 37136 24151
rect 37274 24148 37280 24160
rect 37332 24148 37338 24200
rect 38703 24191 38761 24197
rect 38703 24157 38715 24191
rect 38749 24188 38761 24191
rect 38856 24188 38884 24228
rect 38749 24160 38884 24188
rect 38933 24191 38991 24197
rect 38749 24157 38761 24160
rect 38703 24151 38761 24157
rect 38933 24157 38945 24191
rect 38979 24188 38991 24191
rect 39298 24188 39304 24200
rect 38979 24160 39304 24188
rect 38979 24157 38991 24160
rect 38933 24151 38991 24157
rect 39298 24148 39304 24160
rect 39356 24148 39362 24200
rect 40310 24191 40368 24197
rect 40310 24157 40322 24191
rect 40356 24188 40368 24191
rect 40402 24188 40408 24200
rect 40356 24160 40408 24188
rect 40356 24157 40368 24160
rect 40310 24151 40368 24157
rect 40402 24148 40408 24160
rect 40460 24148 40466 24200
rect 40512 24188 40540 24228
rect 40773 24225 40785 24259
rect 40819 24256 40831 24259
rect 40862 24256 40868 24268
rect 40819 24228 40868 24256
rect 40819 24225 40831 24228
rect 40773 24219 40831 24225
rect 40862 24216 40868 24228
rect 40920 24216 40926 24268
rect 40954 24216 40960 24268
rect 41012 24256 41018 24268
rect 42610 24256 42616 24268
rect 41012 24228 41920 24256
rect 42571 24228 42616 24256
rect 41012 24216 41018 24228
rect 40972 24188 41000 24216
rect 41506 24188 41512 24200
rect 40512 24160 41000 24188
rect 41467 24160 41512 24188
rect 41506 24148 41512 24160
rect 41564 24148 41570 24200
rect 41892 24197 41920 24228
rect 42610 24216 42616 24228
rect 42668 24216 42674 24268
rect 42812 24256 42840 24287
rect 45462 24284 45468 24296
rect 45520 24284 45526 24336
rect 44266 24256 44272 24268
rect 42812 24228 44272 24256
rect 44266 24216 44272 24228
rect 44324 24216 44330 24268
rect 41693 24191 41751 24197
rect 41598 24185 41656 24191
rect 41598 24151 41610 24185
rect 41644 24151 41656 24185
rect 41693 24178 41705 24191
rect 41739 24178 41751 24191
rect 41877 24191 41935 24197
rect 41598 24145 41656 24151
rect 37182 24120 37188 24132
rect 37108 24092 37188 24120
rect 37001 24083 37059 24089
rect 37182 24080 37188 24092
rect 37240 24080 37246 24132
rect 38838 24120 38844 24132
rect 38799 24092 38844 24120
rect 38838 24080 38844 24092
rect 38896 24080 38902 24132
rect 41616 24064 41644 24145
rect 41690 24126 41696 24178
rect 41748 24126 41754 24178
rect 41877 24157 41889 24191
rect 41923 24188 41935 24191
rect 41966 24188 41972 24200
rect 41923 24160 41972 24188
rect 41923 24157 41935 24160
rect 41877 24151 41935 24157
rect 41966 24148 41972 24160
rect 42024 24148 42030 24200
rect 42058 24148 42064 24200
rect 42116 24188 42122 24200
rect 42889 24191 42947 24197
rect 42889 24188 42901 24191
rect 42116 24160 42901 24188
rect 42116 24148 42122 24160
rect 42889 24157 42901 24160
rect 42935 24188 42947 24191
rect 43901 24191 43959 24197
rect 42935 24160 43668 24188
rect 42935 24157 42947 24160
rect 42889 24151 42947 24157
rect 43530 24120 43536 24132
rect 43491 24092 43536 24120
rect 43530 24080 43536 24092
rect 43588 24080 43594 24132
rect 43640 24120 43668 24160
rect 43901 24157 43913 24191
rect 43947 24188 43959 24191
rect 43990 24188 43996 24200
rect 43947 24160 43996 24188
rect 43947 24157 43959 24160
rect 43901 24151 43959 24157
rect 43990 24148 43996 24160
rect 44048 24148 44054 24200
rect 46106 24148 46112 24200
rect 46164 24188 46170 24200
rect 46201 24191 46259 24197
rect 46201 24188 46213 24191
rect 46164 24160 46213 24188
rect 46164 24148 46170 24160
rect 46201 24157 46213 24160
rect 46247 24157 46259 24191
rect 46201 24151 46259 24157
rect 44174 24120 44180 24132
rect 43640 24092 44180 24120
rect 44174 24080 44180 24092
rect 44232 24080 44238 24132
rect 45281 24123 45339 24129
rect 45281 24089 45293 24123
rect 45327 24089 45339 24123
rect 45281 24083 45339 24089
rect 45649 24123 45707 24129
rect 45649 24089 45661 24123
rect 45695 24120 45707 24123
rect 46014 24120 46020 24132
rect 45695 24092 46020 24120
rect 45695 24089 45707 24092
rect 45649 24083 45707 24089
rect 35342 24052 35348 24064
rect 32272 24024 32720 24052
rect 35303 24024 35348 24052
rect 32272 24012 32278 24024
rect 35342 24012 35348 24024
rect 35400 24012 35406 24064
rect 35802 24012 35808 24064
rect 35860 24052 35866 24064
rect 37921 24055 37979 24061
rect 37921 24052 37933 24055
rect 35860 24024 37933 24052
rect 35860 24012 35866 24024
rect 37921 24021 37933 24024
rect 37967 24021 37979 24055
rect 40126 24052 40132 24064
rect 40087 24024 40132 24052
rect 37921 24015 37979 24021
rect 40126 24012 40132 24024
rect 40184 24012 40190 24064
rect 40310 24052 40316 24064
rect 40271 24024 40316 24052
rect 40310 24012 40316 24024
rect 40368 24012 40374 24064
rect 41230 24052 41236 24064
rect 41191 24024 41236 24052
rect 41230 24012 41236 24024
rect 41288 24012 41294 24064
rect 41598 24012 41604 24064
rect 41656 24012 41662 24064
rect 42429 24055 42487 24061
rect 42429 24021 42441 24055
rect 42475 24052 42487 24055
rect 42610 24052 42616 24064
rect 42475 24024 42616 24052
rect 42475 24021 42487 24024
rect 42429 24015 42487 24021
rect 42610 24012 42616 24024
rect 42668 24012 42674 24064
rect 45002 24012 45008 24064
rect 45060 24052 45066 24064
rect 45296 24052 45324 24083
rect 46014 24080 46020 24092
rect 46072 24080 46078 24132
rect 46293 24055 46351 24061
rect 46293 24052 46305 24055
rect 45060 24024 46305 24052
rect 45060 24012 45066 24024
rect 46293 24021 46305 24024
rect 46339 24021 46351 24055
rect 46293 24015 46351 24021
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 29086 23848 29092 23860
rect 29047 23820 29092 23848
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 34330 23848 34336 23860
rect 32692 23820 34336 23848
rect 24397 23783 24455 23789
rect 24397 23749 24409 23783
rect 24443 23780 24455 23783
rect 25038 23780 25044 23792
rect 24443 23752 25044 23780
rect 24443 23749 24455 23752
rect 24397 23743 24455 23749
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 25406 23740 25412 23792
rect 25464 23780 25470 23792
rect 27157 23783 27215 23789
rect 27157 23780 27169 23783
rect 25464 23752 27169 23780
rect 25464 23740 25470 23752
rect 27157 23749 27169 23752
rect 27203 23749 27215 23783
rect 27157 23743 27215 23749
rect 27890 23740 27896 23792
rect 27948 23780 27954 23792
rect 28229 23783 28287 23789
rect 28229 23780 28241 23783
rect 27948 23752 28241 23780
rect 27948 23740 27954 23752
rect 28229 23749 28241 23752
rect 28275 23749 28287 23783
rect 28442 23780 28448 23792
rect 28355 23752 28448 23780
rect 28229 23743 28287 23749
rect 28442 23740 28448 23752
rect 28500 23740 28506 23792
rect 30098 23780 30104 23792
rect 30059 23752 30104 23780
rect 30098 23740 30104 23752
rect 30156 23740 30162 23792
rect 1857 23715 1915 23721
rect 1857 23681 1869 23715
rect 1903 23712 1915 23715
rect 24305 23715 24363 23721
rect 1903 23684 2452 23712
rect 1903 23681 1915 23684
rect 1857 23675 1915 23681
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 2424 23517 2452 23684
rect 24305 23681 24317 23715
rect 24351 23681 24363 23715
rect 24305 23675 24363 23681
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23681 24547 23715
rect 24489 23675 24547 23681
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2498 23508 2504 23520
rect 2455 23480 2504 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2498 23468 2504 23480
rect 2556 23468 2562 23520
rect 24320 23508 24348 23675
rect 24504 23576 24532 23675
rect 24946 23672 24952 23724
rect 25004 23712 25010 23724
rect 25225 23715 25283 23721
rect 25225 23712 25237 23715
rect 25004 23684 25237 23712
rect 25004 23672 25010 23684
rect 25225 23681 25237 23684
rect 25271 23712 25283 23715
rect 25958 23712 25964 23724
rect 25271 23684 25964 23712
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 25958 23672 25964 23684
rect 26016 23672 26022 23724
rect 26605 23715 26663 23721
rect 26605 23681 26617 23715
rect 26651 23712 26663 23715
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 26651 23684 27353 23712
rect 26651 23681 26663 23684
rect 26605 23675 26663 23681
rect 27341 23681 27353 23684
rect 27387 23712 27399 23715
rect 27982 23712 27988 23724
rect 27387 23684 27988 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 28460 23712 28488 23740
rect 28902 23712 28908 23724
rect 28460 23684 28908 23712
rect 28902 23672 28908 23684
rect 28960 23712 28966 23724
rect 29089 23715 29147 23721
rect 29089 23712 29101 23715
rect 28960 23684 29101 23712
rect 28960 23672 28966 23684
rect 29089 23681 29101 23684
rect 29135 23681 29147 23715
rect 29089 23675 29147 23681
rect 29273 23715 29331 23721
rect 29273 23681 29285 23715
rect 29319 23712 29331 23715
rect 30282 23712 30288 23724
rect 29319 23684 30288 23712
rect 29319 23681 29331 23684
rect 29273 23675 29331 23681
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 32692 23721 32720 23820
rect 34330 23808 34336 23820
rect 34388 23808 34394 23860
rect 37461 23851 37519 23857
rect 37461 23817 37473 23851
rect 37507 23817 37519 23851
rect 37461 23811 37519 23817
rect 37476 23780 37504 23811
rect 39298 23808 39304 23860
rect 39356 23848 39362 23860
rect 41506 23848 41512 23860
rect 39356 23820 41512 23848
rect 39356 23808 39362 23820
rect 41506 23808 41512 23820
rect 41564 23848 41570 23860
rect 42426 23848 42432 23860
rect 41564 23820 42432 23848
rect 41564 23808 41570 23820
rect 42426 23808 42432 23820
rect 42484 23848 42490 23860
rect 43346 23848 43352 23860
rect 42484 23820 43352 23848
rect 42484 23808 42490 23820
rect 43346 23808 43352 23820
rect 43404 23808 43410 23860
rect 44542 23857 44548 23860
rect 44520 23851 44548 23857
rect 44520 23817 44532 23851
rect 44520 23811 44548 23817
rect 44542 23808 44548 23811
rect 44600 23808 44606 23860
rect 41969 23783 42027 23789
rect 41969 23780 41981 23783
rect 32968 23752 37504 23780
rect 39684 23752 41981 23780
rect 32968 23724 32996 23752
rect 39684 23724 39712 23752
rect 41969 23749 41981 23752
rect 42015 23780 42027 23783
rect 43530 23780 43536 23792
rect 42015 23752 43536 23780
rect 42015 23749 42027 23752
rect 41969 23743 42027 23749
rect 43530 23740 43536 23752
rect 43588 23740 43594 23792
rect 43806 23740 43812 23792
rect 43864 23780 43870 23792
rect 43864 23752 44128 23780
rect 43864 23740 43870 23752
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23712 31631 23715
rect 32493 23715 32551 23721
rect 32493 23712 32505 23715
rect 31619 23684 32505 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 32493 23681 32505 23684
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23681 32735 23715
rect 32950 23712 32956 23724
rect 32863 23684 32956 23712
rect 32677 23675 32735 23681
rect 32950 23672 32956 23684
rect 33008 23672 33014 23724
rect 33137 23715 33195 23721
rect 33137 23681 33149 23715
rect 33183 23712 33195 23715
rect 33502 23712 33508 23724
rect 33183 23684 33508 23712
rect 33183 23681 33195 23684
rect 33137 23675 33195 23681
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 33686 23672 33692 23724
rect 33744 23712 33750 23724
rect 33965 23715 34023 23721
rect 33965 23712 33977 23715
rect 33744 23684 33977 23712
rect 33744 23672 33750 23684
rect 33965 23681 33977 23684
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 34793 23715 34851 23721
rect 34793 23681 34805 23715
rect 34839 23681 34851 23715
rect 34793 23675 34851 23681
rect 25130 23644 25136 23656
rect 25091 23616 25136 23644
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25317 23647 25375 23653
rect 25317 23613 25329 23647
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 25409 23647 25467 23653
rect 25409 23613 25421 23647
rect 25455 23644 25467 23647
rect 25590 23644 25596 23656
rect 25455 23616 25596 23644
rect 25455 23613 25467 23616
rect 25409 23607 25467 23613
rect 25332 23576 25360 23607
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 26329 23647 26387 23653
rect 26329 23613 26341 23647
rect 26375 23644 26387 23647
rect 27617 23647 27675 23653
rect 27617 23644 27629 23647
rect 26375 23616 27629 23644
rect 26375 23613 26387 23616
rect 26329 23607 26387 23613
rect 27617 23613 27629 23616
rect 27663 23644 27675 23647
rect 27663 23616 28120 23644
rect 27663 23613 27675 23616
rect 27617 23607 27675 23613
rect 26142 23576 26148 23588
rect 24504 23548 25268 23576
rect 25332 23548 26148 23576
rect 25240 23520 25268 23548
rect 26142 23536 26148 23548
rect 26200 23536 26206 23588
rect 26513 23579 26571 23585
rect 26513 23545 26525 23579
rect 26559 23576 26571 23579
rect 27246 23576 27252 23588
rect 26559 23548 27252 23576
rect 26559 23545 26571 23548
rect 26513 23539 26571 23545
rect 27246 23536 27252 23548
rect 27304 23576 27310 23588
rect 28092 23585 28120 23616
rect 28258 23604 28264 23656
rect 28316 23644 28322 23656
rect 31665 23647 31723 23653
rect 28316 23616 31248 23644
rect 28316 23604 28322 23616
rect 27525 23579 27583 23585
rect 27525 23576 27537 23579
rect 27304 23548 27537 23576
rect 27304 23536 27310 23548
rect 27525 23545 27537 23548
rect 27571 23545 27583 23579
rect 27525 23539 27583 23545
rect 28077 23579 28135 23585
rect 28077 23545 28089 23579
rect 28123 23545 28135 23579
rect 28077 23539 28135 23545
rect 24854 23508 24860 23520
rect 24320 23480 24860 23508
rect 24854 23468 24860 23480
rect 24912 23468 24918 23520
rect 25222 23468 25228 23520
rect 25280 23508 25286 23520
rect 28276 23517 28304 23604
rect 30469 23579 30527 23585
rect 30469 23545 30481 23579
rect 30515 23576 30527 23579
rect 30742 23576 30748 23588
rect 30515 23548 30748 23576
rect 30515 23545 30527 23548
rect 30469 23539 30527 23545
rect 30742 23536 30748 23548
rect 30800 23536 30806 23588
rect 31220 23585 31248 23616
rect 31665 23613 31677 23647
rect 31711 23644 31723 23647
rect 31754 23644 31760 23656
rect 31711 23616 31760 23644
rect 31711 23613 31723 23616
rect 31665 23607 31723 23613
rect 31754 23604 31760 23616
rect 31812 23604 31818 23656
rect 33594 23644 33600 23656
rect 33555 23616 33600 23644
rect 33594 23604 33600 23616
rect 33652 23604 33658 23656
rect 34808 23644 34836 23675
rect 35526 23672 35532 23724
rect 35584 23712 35590 23724
rect 35802 23712 35808 23724
rect 35584 23684 35808 23712
rect 35584 23672 35590 23684
rect 35802 23672 35808 23684
rect 35860 23672 35866 23724
rect 36722 23672 36728 23724
rect 36780 23712 36786 23724
rect 36817 23715 36875 23721
rect 36817 23712 36829 23715
rect 36780 23684 36829 23712
rect 36780 23672 36786 23684
rect 36817 23681 36829 23684
rect 36863 23681 36875 23715
rect 37366 23712 37372 23724
rect 36817 23675 36875 23681
rect 36924 23684 37372 23712
rect 33704 23616 34836 23644
rect 31205 23579 31263 23585
rect 31205 23545 31217 23579
rect 31251 23545 31263 23579
rect 31205 23539 31263 23545
rect 26421 23511 26479 23517
rect 26421 23508 26433 23511
rect 25280 23480 26433 23508
rect 25280 23468 25286 23480
rect 26421 23477 26433 23480
rect 26467 23477 26479 23511
rect 26421 23471 26479 23477
rect 28261 23511 28319 23517
rect 28261 23477 28273 23511
rect 28307 23477 28319 23511
rect 30558 23508 30564 23520
rect 30519 23480 30564 23508
rect 28261 23471 28319 23477
rect 30558 23468 30564 23480
rect 30616 23468 30622 23520
rect 33704 23517 33732 23616
rect 34808 23576 34836 23616
rect 35250 23604 35256 23656
rect 35308 23644 35314 23656
rect 35897 23647 35955 23653
rect 35897 23644 35909 23647
rect 35308 23616 35909 23644
rect 35308 23604 35314 23616
rect 35897 23613 35909 23616
rect 35943 23644 35955 23647
rect 36924 23644 36952 23684
rect 37366 23672 37372 23684
rect 37424 23672 37430 23724
rect 37645 23715 37703 23721
rect 37645 23681 37657 23715
rect 37691 23712 37703 23715
rect 38010 23712 38016 23724
rect 37691 23684 38016 23712
rect 37691 23681 37703 23684
rect 37645 23675 37703 23681
rect 38010 23672 38016 23684
rect 38068 23672 38074 23724
rect 38657 23715 38715 23721
rect 38657 23681 38669 23715
rect 38703 23712 38715 23715
rect 39482 23712 39488 23724
rect 38703 23684 39488 23712
rect 38703 23681 38715 23684
rect 38657 23675 38715 23681
rect 39482 23672 39488 23684
rect 39540 23672 39546 23724
rect 39666 23712 39672 23724
rect 39627 23684 39672 23712
rect 39666 23672 39672 23684
rect 39724 23672 39730 23724
rect 39758 23672 39764 23724
rect 39816 23712 39822 23724
rect 40865 23715 40923 23721
rect 40865 23712 40877 23715
rect 39816 23684 40877 23712
rect 39816 23672 39822 23684
rect 40865 23681 40877 23684
rect 40911 23681 40923 23715
rect 41138 23712 41144 23724
rect 41099 23684 41144 23712
rect 40865 23675 40923 23681
rect 35943 23616 36952 23644
rect 35943 23613 35955 23616
rect 35897 23607 35955 23613
rect 36998 23604 37004 23656
rect 37056 23644 37062 23656
rect 37737 23647 37795 23653
rect 37737 23644 37749 23647
rect 37056 23616 37749 23644
rect 37056 23604 37062 23616
rect 37737 23613 37749 23616
rect 37783 23613 37795 23647
rect 37737 23607 37795 23613
rect 37829 23647 37887 23653
rect 37829 23613 37841 23647
rect 37875 23613 37887 23647
rect 37829 23607 37887 23613
rect 37844 23576 37872 23607
rect 37918 23604 37924 23656
rect 37976 23644 37982 23656
rect 38562 23644 38568 23656
rect 37976 23616 38568 23644
rect 37976 23604 37982 23616
rect 38562 23604 38568 23616
rect 38620 23604 38626 23656
rect 39500 23644 39528 23672
rect 39850 23644 39856 23656
rect 39500 23616 39856 23644
rect 39850 23604 39856 23616
rect 39908 23604 39914 23656
rect 40678 23644 40684 23656
rect 40639 23616 40684 23644
rect 40678 23604 40684 23616
rect 40736 23604 40742 23656
rect 40880 23644 40908 23675
rect 41138 23672 41144 23684
rect 41196 23672 41202 23724
rect 43162 23712 43168 23724
rect 43123 23684 43168 23712
rect 43162 23672 43168 23684
rect 43220 23672 43226 23724
rect 43438 23712 43444 23724
rect 43351 23684 43444 23712
rect 43438 23672 43444 23684
rect 43496 23712 43502 23724
rect 43622 23712 43628 23724
rect 43496 23684 43628 23712
rect 43496 23672 43502 23684
rect 43622 23672 43628 23684
rect 43680 23672 43686 23724
rect 44100 23721 44128 23752
rect 44085 23715 44143 23721
rect 44085 23681 44097 23715
rect 44131 23681 44143 23715
rect 44085 23675 44143 23681
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44232 23684 44833 23712
rect 44232 23672 44238 23684
rect 44821 23681 44833 23684
rect 44867 23712 44879 23715
rect 46106 23712 46112 23724
rect 44867 23684 46112 23712
rect 44867 23681 44879 23684
rect 44821 23675 44879 23681
rect 46106 23672 46112 23684
rect 46164 23672 46170 23724
rect 42058 23644 42064 23656
rect 40880 23616 42064 23644
rect 42058 23604 42064 23616
rect 42116 23604 42122 23656
rect 42702 23604 42708 23656
rect 42760 23644 42766 23656
rect 44910 23644 44916 23656
rect 42760 23630 44022 23644
rect 42760 23616 44036 23630
rect 44871 23616 44916 23644
rect 42760 23604 42766 23616
rect 39758 23576 39764 23588
rect 34808 23548 36860 23576
rect 37844 23548 39764 23576
rect 36832 23520 36860 23548
rect 39758 23536 39764 23548
rect 39816 23536 39822 23588
rect 41049 23579 41107 23585
rect 41049 23545 41061 23579
rect 41095 23576 41107 23579
rect 44008 23576 44036 23616
rect 44910 23604 44916 23616
rect 44968 23604 44974 23656
rect 45554 23576 45560 23588
rect 41095 23548 43576 23576
rect 44008 23548 45560 23576
rect 41095 23545 41107 23548
rect 41049 23539 41107 23545
rect 43548 23520 43576 23548
rect 45554 23536 45560 23548
rect 45612 23576 45618 23588
rect 45741 23579 45799 23585
rect 45741 23576 45753 23579
rect 45612 23548 45753 23576
rect 45612 23536 45618 23548
rect 45741 23545 45753 23548
rect 45787 23545 45799 23579
rect 45741 23539 45799 23545
rect 33689 23511 33747 23517
rect 33689 23477 33701 23511
rect 33735 23477 33747 23511
rect 33689 23471 33747 23477
rect 33778 23468 33784 23520
rect 33836 23508 33842 23520
rect 33965 23511 34023 23517
rect 33836 23480 33881 23508
rect 33836 23468 33842 23480
rect 33965 23477 33977 23511
rect 34011 23508 34023 23511
rect 34422 23508 34428 23520
rect 34011 23480 34428 23508
rect 34011 23477 34023 23480
rect 33965 23471 34023 23477
rect 34422 23468 34428 23480
rect 34480 23468 34486 23520
rect 34514 23468 34520 23520
rect 34572 23508 34578 23520
rect 34572 23480 34617 23508
rect 34572 23468 34578 23480
rect 34698 23468 34704 23520
rect 34756 23508 34762 23520
rect 35250 23508 35256 23520
rect 34756 23480 35256 23508
rect 34756 23468 34762 23480
rect 35250 23468 35256 23480
rect 35308 23468 35314 23520
rect 35986 23508 35992 23520
rect 35947 23480 35992 23508
rect 35986 23468 35992 23480
rect 36044 23468 36050 23520
rect 36173 23511 36231 23517
rect 36173 23477 36185 23511
rect 36219 23508 36231 23511
rect 36446 23508 36452 23520
rect 36219 23480 36452 23508
rect 36219 23477 36231 23480
rect 36173 23471 36231 23477
rect 36446 23468 36452 23480
rect 36504 23468 36510 23520
rect 36538 23468 36544 23520
rect 36596 23508 36602 23520
rect 36725 23511 36783 23517
rect 36725 23508 36737 23511
rect 36596 23480 36737 23508
rect 36596 23468 36602 23480
rect 36725 23477 36737 23480
rect 36771 23477 36783 23511
rect 36725 23471 36783 23477
rect 36814 23468 36820 23520
rect 36872 23508 36878 23520
rect 38749 23511 38807 23517
rect 38749 23508 38761 23511
rect 36872 23480 38761 23508
rect 36872 23468 36878 23480
rect 38749 23477 38761 23480
rect 38795 23477 38807 23511
rect 38749 23471 38807 23477
rect 39206 23468 39212 23520
rect 39264 23508 39270 23520
rect 39485 23511 39543 23517
rect 39485 23508 39497 23511
rect 39264 23480 39497 23508
rect 39264 23468 39270 23480
rect 39485 23477 39497 23480
rect 39531 23477 39543 23511
rect 39485 23471 39543 23477
rect 40126 23468 40132 23520
rect 40184 23508 40190 23520
rect 40862 23508 40868 23520
rect 40184 23480 40868 23508
rect 40184 23468 40190 23480
rect 40862 23468 40868 23480
rect 40920 23468 40926 23520
rect 41506 23468 41512 23520
rect 41564 23508 41570 23520
rect 41693 23511 41751 23517
rect 41693 23508 41705 23511
rect 41564 23480 41705 23508
rect 41564 23468 41570 23480
rect 41693 23477 41705 23480
rect 41739 23477 41751 23511
rect 42978 23508 42984 23520
rect 42939 23480 42984 23508
rect 41693 23471 41751 23477
rect 42978 23468 42984 23480
rect 43036 23468 43042 23520
rect 43530 23468 43536 23520
rect 43588 23508 43594 23520
rect 44910 23508 44916 23520
rect 43588 23480 44916 23508
rect 43588 23468 43594 23480
rect 44910 23468 44916 23480
rect 44968 23468 44974 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23273 23535 23307
rect 23477 23267 23535 23273
rect 23492 23236 23520 23267
rect 24854 23264 24860 23316
rect 24912 23304 24918 23316
rect 25406 23304 25412 23316
rect 24912 23276 25412 23304
rect 24912 23264 24918 23276
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 33778 23264 33784 23316
rect 33836 23304 33842 23316
rect 34238 23304 34244 23316
rect 33836 23276 34244 23304
rect 33836 23264 33842 23276
rect 34238 23264 34244 23276
rect 34296 23264 34302 23316
rect 35434 23264 35440 23316
rect 35492 23304 35498 23316
rect 35897 23307 35955 23313
rect 35492 23276 35756 23304
rect 35492 23264 35498 23276
rect 35728 23248 35756 23276
rect 35897 23273 35909 23307
rect 35943 23304 35955 23307
rect 38654 23304 38660 23316
rect 35943 23276 38660 23304
rect 35943 23273 35955 23276
rect 35897 23267 35955 23273
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 38838 23264 38844 23316
rect 38896 23304 38902 23316
rect 39482 23304 39488 23316
rect 38896 23276 39488 23304
rect 38896 23264 38902 23276
rect 39482 23264 39488 23276
rect 39540 23304 39546 23316
rect 45002 23304 45008 23316
rect 39540 23276 45008 23304
rect 39540 23264 39546 23276
rect 45002 23264 45008 23276
rect 45060 23264 45066 23316
rect 23842 23236 23848 23248
rect 23492 23208 23848 23236
rect 23842 23196 23848 23208
rect 23900 23236 23906 23248
rect 31113 23239 31171 23245
rect 31113 23236 31125 23239
rect 23900 23208 31125 23236
rect 23900 23196 23906 23208
rect 31113 23205 31125 23208
rect 31159 23205 31171 23239
rect 35250 23236 35256 23248
rect 31113 23199 31171 23205
rect 33428 23208 35256 23236
rect 26418 23168 26424 23180
rect 26379 23140 26424 23168
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27433 23171 27491 23177
rect 27433 23168 27445 23171
rect 27212 23140 27445 23168
rect 27212 23128 27218 23140
rect 27433 23137 27445 23140
rect 27479 23137 27491 23171
rect 27890 23168 27896 23180
rect 27851 23140 27896 23168
rect 27433 23131 27491 23137
rect 27890 23128 27896 23140
rect 27948 23128 27954 23180
rect 28629 23171 28687 23177
rect 28629 23137 28641 23171
rect 28675 23168 28687 23171
rect 28902 23168 28908 23180
rect 28675 23140 28908 23168
rect 28675 23137 28687 23140
rect 28629 23131 28687 23137
rect 28902 23128 28908 23140
rect 28960 23168 28966 23180
rect 29181 23171 29239 23177
rect 29181 23168 29193 23171
rect 28960 23140 29193 23168
rect 28960 23128 28966 23140
rect 29181 23137 29193 23140
rect 29227 23168 29239 23171
rect 29227 23140 30420 23168
rect 29227 23137 29239 23140
rect 29181 23131 29239 23137
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 22005 23103 22063 23109
rect 22005 23069 22017 23103
rect 22051 23100 22063 23103
rect 22830 23100 22836 23112
rect 22051 23072 22836 23100
rect 22051 23069 22063 23072
rect 22005 23063 22063 23069
rect 21928 23032 21956 23063
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23100 23259 23103
rect 23566 23100 23572 23112
rect 23247 23072 23572 23100
rect 23247 23069 23259 23072
rect 23201 23063 23259 23069
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 25133 23103 25191 23109
rect 25133 23069 25145 23103
rect 25179 23100 25191 23103
rect 25222 23100 25228 23112
rect 25179 23072 25228 23100
rect 25179 23069 25191 23072
rect 25133 23063 25191 23069
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 25406 23100 25412 23112
rect 25367 23072 25412 23100
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 25590 23100 25596 23112
rect 25551 23072 25596 23100
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23069 26111 23103
rect 26053 23063 26111 23069
rect 22278 23032 22284 23044
rect 21928 23004 22284 23032
rect 22278 22992 22284 23004
rect 22336 23032 22342 23044
rect 24578 23032 24584 23044
rect 22336 23004 24584 23032
rect 22336 22992 22342 23004
rect 24578 22992 24584 23004
rect 24636 22992 24642 23044
rect 26068 23032 26096 23063
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 26200 23072 26249 23100
rect 26200 23060 26206 23072
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 27798 23100 27804 23112
rect 27759 23072 27804 23100
rect 26237 23063 26295 23069
rect 27798 23060 27804 23072
rect 27856 23060 27862 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29052 23072 29745 23100
rect 29052 23060 29058 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 30282 23100 30288 23112
rect 30195 23072 30288 23100
rect 29733 23063 29791 23069
rect 30282 23060 30288 23072
rect 30340 23060 30346 23112
rect 30392 23100 30420 23140
rect 30558 23128 30564 23180
rect 30616 23168 30622 23180
rect 30837 23171 30895 23177
rect 30837 23168 30849 23171
rect 30616 23140 30849 23168
rect 30616 23128 30622 23140
rect 30837 23137 30849 23140
rect 30883 23137 30895 23171
rect 32398 23168 32404 23180
rect 32359 23140 32404 23168
rect 30837 23131 30895 23137
rect 32398 23128 32404 23140
rect 32456 23128 32462 23180
rect 30745 23103 30803 23109
rect 30745 23100 30757 23103
rect 30392 23072 30757 23100
rect 30745 23069 30757 23072
rect 30791 23100 30803 23103
rect 31386 23100 31392 23112
rect 30791 23072 31392 23100
rect 30791 23069 30803 23072
rect 30745 23063 30803 23069
rect 31386 23060 31392 23072
rect 31444 23060 31450 23112
rect 31754 23060 31760 23112
rect 31812 23100 31818 23112
rect 32309 23103 32367 23109
rect 32309 23100 32321 23103
rect 31812 23072 32321 23100
rect 31812 23060 31818 23072
rect 32309 23069 32321 23072
rect 32355 23069 32367 23103
rect 33226 23100 33232 23112
rect 33187 23072 33232 23100
rect 32309 23063 32367 23069
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 33428 23109 33456 23208
rect 35250 23196 35256 23208
rect 35308 23196 35314 23248
rect 35710 23196 35716 23248
rect 35768 23236 35774 23248
rect 37182 23236 37188 23248
rect 35768 23208 37188 23236
rect 35768 23196 35774 23208
rect 37182 23196 37188 23208
rect 37240 23236 37246 23248
rect 39114 23236 39120 23248
rect 37240 23208 39120 23236
rect 37240 23196 37246 23208
rect 39114 23196 39120 23208
rect 39172 23196 39178 23248
rect 40586 23196 40592 23248
rect 40644 23236 40650 23248
rect 43346 23236 43352 23248
rect 40644 23208 43352 23236
rect 40644 23196 40650 23208
rect 43346 23196 43352 23208
rect 43404 23196 43410 23248
rect 43530 23236 43536 23248
rect 43491 23208 43536 23236
rect 43530 23196 43536 23208
rect 43588 23196 43594 23248
rect 34238 23128 34244 23180
rect 34296 23168 34302 23180
rect 34296 23140 34928 23168
rect 34296 23128 34302 23140
rect 33413 23103 33471 23109
rect 33413 23069 33425 23103
rect 33459 23069 33471 23103
rect 33413 23063 33471 23069
rect 34149 23103 34207 23109
rect 34149 23069 34161 23103
rect 34195 23069 34207 23103
rect 34149 23063 34207 23069
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23100 34391 23103
rect 34606 23100 34612 23112
rect 34379 23072 34612 23100
rect 34379 23069 34391 23072
rect 34333 23063 34391 23069
rect 25148 23004 26096 23032
rect 25148 22976 25176 23004
rect 21726 22964 21732 22976
rect 21687 22936 21732 22964
rect 21726 22924 21732 22936
rect 21784 22924 21790 22976
rect 22373 22967 22431 22973
rect 22373 22933 22385 22967
rect 22419 22964 22431 22967
rect 23658 22964 23664 22976
rect 22419 22936 23664 22964
rect 22419 22933 22431 22936
rect 22373 22927 22431 22933
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 24949 22967 25007 22973
rect 24949 22964 24961 22967
rect 24820 22936 24961 22964
rect 24820 22924 24826 22936
rect 24949 22933 24961 22936
rect 24995 22933 25007 22967
rect 24949 22927 25007 22933
rect 25130 22924 25136 22976
rect 25188 22924 25194 22976
rect 30300 22964 30328 23060
rect 34164 23032 34192 23063
rect 34606 23060 34612 23072
rect 34664 23060 34670 23112
rect 34900 23109 34928 23140
rect 35434 23128 35440 23180
rect 35492 23168 35498 23180
rect 36633 23171 36691 23177
rect 36633 23168 36645 23171
rect 35492 23140 36645 23168
rect 35492 23128 35498 23140
rect 36633 23137 36645 23140
rect 36679 23137 36691 23171
rect 38470 23168 38476 23180
rect 36633 23131 36691 23137
rect 36925 23140 38476 23168
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23069 34943 23103
rect 34885 23063 34943 23069
rect 35069 23103 35127 23109
rect 35069 23069 35081 23103
rect 35115 23100 35127 23103
rect 35342 23100 35348 23112
rect 35115 23072 35348 23100
rect 35115 23069 35127 23072
rect 35069 23063 35127 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 35618 23032 35624 23044
rect 34164 23004 35624 23032
rect 35618 22992 35624 23004
rect 35676 22992 35682 23044
rect 35710 22992 35716 23044
rect 35768 23032 35774 23044
rect 35929 23035 35987 23041
rect 35768 23004 35813 23032
rect 35768 22992 35774 23004
rect 35929 23001 35941 23035
rect 35975 23032 35987 23035
rect 36354 23032 36360 23044
rect 35975 23004 36360 23032
rect 35975 23001 35987 23004
rect 35929 22995 35987 23001
rect 36354 22992 36360 23004
rect 36412 22992 36418 23044
rect 36556 23032 36584 23063
rect 36722 23060 36728 23112
rect 36780 23100 36786 23112
rect 36925 23100 36953 23140
rect 38470 23128 38476 23140
rect 38528 23128 38534 23180
rect 40313 23171 40371 23177
rect 38948 23140 39896 23168
rect 36780 23072 36953 23100
rect 36780 23060 36786 23072
rect 37274 23060 37280 23112
rect 37332 23100 37338 23112
rect 38948 23109 38976 23140
rect 37553 23103 37611 23109
rect 37553 23100 37565 23103
rect 37332 23072 37565 23100
rect 37332 23060 37338 23072
rect 37553 23069 37565 23072
rect 37599 23069 37611 23103
rect 38933 23103 38991 23109
rect 38933 23100 38945 23103
rect 37553 23063 37611 23069
rect 37660 23072 38945 23100
rect 36906 23032 36912 23044
rect 36556 23004 36912 23032
rect 36906 22992 36912 23004
rect 36964 23032 36970 23044
rect 37660 23032 37688 23072
rect 38933 23069 38945 23072
rect 38979 23069 38991 23103
rect 39298 23100 39304 23112
rect 39259 23072 39304 23100
rect 38933 23063 38991 23069
rect 39298 23060 39304 23072
rect 39356 23060 39362 23112
rect 39393 23103 39451 23109
rect 39393 23069 39405 23103
rect 39439 23100 39451 23103
rect 39482 23100 39488 23112
rect 39439 23072 39488 23100
rect 39439 23069 39451 23072
rect 39393 23063 39451 23069
rect 39482 23060 39488 23072
rect 39540 23060 39546 23112
rect 38749 23035 38807 23041
rect 38749 23032 38761 23035
rect 36964 23004 37688 23032
rect 37752 23004 38761 23032
rect 36964 22992 36970 23004
rect 31665 22967 31723 22973
rect 31665 22964 31677 22967
rect 30300 22936 31677 22964
rect 31665 22933 31677 22936
rect 31711 22933 31723 22967
rect 31665 22927 31723 22933
rect 32766 22924 32772 22976
rect 32824 22964 32830 22976
rect 33321 22967 33379 22973
rect 33321 22964 33333 22967
rect 32824 22936 33333 22964
rect 32824 22924 32830 22936
rect 33321 22933 33333 22936
rect 33367 22933 33379 22967
rect 33321 22927 33379 22933
rect 33410 22924 33416 22976
rect 33468 22964 33474 22976
rect 34977 22967 35035 22973
rect 34977 22964 34989 22967
rect 33468 22936 34989 22964
rect 33468 22924 33474 22936
rect 34977 22933 34989 22936
rect 35023 22933 35035 22967
rect 36078 22964 36084 22976
rect 36039 22936 36084 22964
rect 34977 22927 35035 22933
rect 36078 22924 36084 22936
rect 36136 22924 36142 22976
rect 37182 22924 37188 22976
rect 37240 22964 37246 22976
rect 37752 22964 37780 23004
rect 38749 23001 38761 23004
rect 38795 23001 38807 23035
rect 39868 23032 39896 23140
rect 40313 23137 40325 23171
rect 40359 23168 40371 23171
rect 41877 23171 41935 23177
rect 41877 23168 41889 23171
rect 40359 23140 41889 23168
rect 40359 23137 40371 23140
rect 40313 23131 40371 23137
rect 41877 23137 41889 23140
rect 41923 23137 41935 23171
rect 42978 23168 42984 23180
rect 41877 23131 41935 23137
rect 42076 23140 42984 23168
rect 39942 23060 39948 23112
rect 40000 23100 40006 23112
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 40000 23072 40233 23100
rect 40000 23060 40006 23072
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 40221 23063 40279 23069
rect 40405 23103 40463 23109
rect 40405 23069 40417 23103
rect 40451 23069 40463 23103
rect 40405 23063 40463 23069
rect 40497 23103 40555 23109
rect 40497 23069 40509 23103
rect 40543 23100 40555 23103
rect 40586 23100 40592 23112
rect 40543 23072 40592 23100
rect 40543 23069 40555 23072
rect 40497 23063 40555 23069
rect 40420 23032 40448 23063
rect 40586 23060 40592 23072
rect 40644 23060 40650 23112
rect 40681 23103 40739 23109
rect 40681 23069 40693 23103
rect 40727 23100 40739 23103
rect 40862 23100 40868 23112
rect 40727 23072 40868 23100
rect 40727 23069 40739 23072
rect 40681 23063 40739 23069
rect 40862 23060 40868 23072
rect 40920 23060 40926 23112
rect 41230 23100 41236 23112
rect 41191 23072 41236 23100
rect 41230 23060 41236 23072
rect 41288 23060 41294 23112
rect 41414 23060 41420 23112
rect 41472 23100 41478 23112
rect 42076 23109 42104 23140
rect 42978 23128 42984 23140
rect 43036 23128 43042 23180
rect 42061 23103 42119 23109
rect 41472 23072 41517 23100
rect 41472 23060 41478 23072
rect 42061 23069 42073 23103
rect 42107 23069 42119 23103
rect 42061 23063 42119 23069
rect 42153 23103 42211 23109
rect 42153 23069 42165 23103
rect 42199 23069 42211 23103
rect 42702 23100 42708 23112
rect 42663 23072 42708 23100
rect 42153 23063 42211 23069
rect 41138 23032 41144 23044
rect 39868 23004 40265 23032
rect 40420 23004 41144 23032
rect 38749 22995 38807 23001
rect 37240 22936 37780 22964
rect 37829 22967 37887 22973
rect 37240 22924 37246 22936
rect 37829 22933 37841 22967
rect 37875 22964 37887 22967
rect 38654 22964 38660 22976
rect 37875 22936 38660 22964
rect 37875 22933 37887 22936
rect 37829 22927 37887 22933
rect 38654 22924 38660 22936
rect 38712 22924 38718 22976
rect 40034 22964 40040 22976
rect 39995 22936 40040 22964
rect 40034 22924 40040 22936
rect 40092 22924 40098 22976
rect 40237 22964 40265 23004
rect 41138 22992 41144 23004
rect 41196 22992 41202 23044
rect 41782 23032 41788 23044
rect 41432 23004 41788 23032
rect 40954 22964 40960 22976
rect 40237 22936 40960 22964
rect 40954 22924 40960 22936
rect 41012 22924 41018 22976
rect 41325 22967 41383 22973
rect 41325 22933 41337 22967
rect 41371 22964 41383 22967
rect 41432 22964 41460 23004
rect 41782 22992 41788 23004
rect 41840 23032 41846 23044
rect 42168 23032 42196 23063
rect 42702 23060 42708 23072
rect 42760 23060 42766 23112
rect 45554 23100 45560 23112
rect 45515 23072 45560 23100
rect 45554 23060 45560 23072
rect 45612 23100 45618 23112
rect 46106 23100 46112 23112
rect 45612 23072 46112 23100
rect 45612 23060 45618 23072
rect 46106 23060 46112 23072
rect 46164 23060 46170 23112
rect 43806 23032 43812 23044
rect 41840 23004 42196 23032
rect 43767 23004 43812 23032
rect 41840 22992 41846 23004
rect 43806 22992 43812 23004
rect 43864 22992 43870 23044
rect 44634 22992 44640 23044
rect 44692 23032 44698 23044
rect 45189 23035 45247 23041
rect 45189 23032 45201 23035
rect 44692 23004 45201 23032
rect 44692 22992 44698 23004
rect 45189 23001 45201 23004
rect 45235 23001 45247 23035
rect 45189 22995 45247 23001
rect 41371 22936 41460 22964
rect 41371 22933 41383 22936
rect 41325 22927 41383 22933
rect 43162 22924 43168 22976
rect 43220 22964 43226 22976
rect 43349 22967 43407 22973
rect 43349 22964 43361 22967
rect 43220 22936 43361 22964
rect 43220 22924 43226 22936
rect 43349 22933 43361 22936
rect 43395 22964 43407 22967
rect 43622 22964 43628 22976
rect 43395 22936 43628 22964
rect 43395 22933 43407 22936
rect 43349 22927 43407 22933
rect 43622 22924 43628 22936
rect 43680 22924 43686 22976
rect 43990 22924 43996 22976
rect 44048 22964 44054 22976
rect 44269 22967 44327 22973
rect 44269 22964 44281 22967
rect 44048 22936 44281 22964
rect 44048 22924 44054 22936
rect 44269 22933 44281 22936
rect 44315 22933 44327 22967
rect 44269 22927 44327 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 22830 22760 22836 22772
rect 22791 22732 22836 22760
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 24578 22760 24584 22772
rect 24539 22732 24584 22760
rect 24578 22720 24584 22732
rect 24636 22720 24642 22772
rect 24946 22760 24952 22772
rect 24907 22732 24952 22760
rect 24946 22720 24952 22732
rect 25004 22720 25010 22772
rect 27246 22760 27252 22772
rect 27207 22732 27252 22760
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 27801 22763 27859 22769
rect 27801 22729 27813 22763
rect 27847 22760 27859 22763
rect 27890 22760 27896 22772
rect 27847 22732 27896 22760
rect 27847 22729 27859 22732
rect 27801 22723 27859 22729
rect 27890 22720 27896 22732
rect 27948 22720 27954 22772
rect 32398 22760 32404 22772
rect 32359 22732 32404 22760
rect 32398 22720 32404 22732
rect 32456 22720 32462 22772
rect 32766 22760 32772 22772
rect 32727 22732 32772 22760
rect 32766 22720 32772 22732
rect 32824 22720 32830 22772
rect 34054 22760 34060 22772
rect 32876 22732 34060 22760
rect 26142 22692 26148 22704
rect 24872 22664 26148 22692
rect 24872 22636 24900 22664
rect 26142 22652 26148 22664
rect 26200 22652 26206 22704
rect 28994 22692 29000 22704
rect 28955 22664 29000 22692
rect 28994 22652 29000 22664
rect 29052 22652 29058 22704
rect 30745 22695 30803 22701
rect 30745 22661 30757 22695
rect 30791 22692 30803 22695
rect 32306 22692 32312 22704
rect 30791 22664 32312 22692
rect 30791 22661 30803 22664
rect 30745 22655 30803 22661
rect 32306 22652 32312 22664
rect 32364 22652 32370 22704
rect 23566 22624 23572 22636
rect 23527 22596 23572 22624
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 23842 22624 23848 22636
rect 23803 22596 23848 22624
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 24762 22624 24768 22636
rect 24723 22596 24768 22624
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 24854 22584 24860 22636
rect 24912 22624 24918 22636
rect 24912 22596 25005 22624
rect 24912 22584 24918 22596
rect 25038 22584 25044 22636
rect 25096 22624 25102 22636
rect 25225 22627 25283 22633
rect 25225 22624 25237 22627
rect 25096 22596 25237 22624
rect 25096 22584 25102 22596
rect 25225 22593 25237 22596
rect 25271 22593 25283 22627
rect 27154 22624 27160 22636
rect 27115 22596 27160 22624
rect 25225 22587 25283 22593
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22593 27399 22627
rect 28166 22624 28172 22636
rect 28127 22596 28172 22624
rect 27341 22587 27399 22593
rect 25130 22556 25136 22568
rect 25091 22528 25136 22556
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 26970 22516 26976 22568
rect 27028 22556 27034 22568
rect 27356 22556 27384 22587
rect 28166 22584 28172 22596
rect 28224 22584 28230 22636
rect 28261 22627 28319 22633
rect 28261 22593 28273 22627
rect 28307 22624 28319 22627
rect 30929 22627 30987 22633
rect 28307 22596 29316 22624
rect 28307 22593 28319 22596
rect 28261 22587 28319 22593
rect 27028 22528 27384 22556
rect 28445 22559 28503 22565
rect 27028 22516 27034 22528
rect 28445 22525 28457 22559
rect 28491 22525 28503 22559
rect 29288 22556 29316 22596
rect 29822 22556 29828 22568
rect 29288 22528 29828 22556
rect 28445 22519 28503 22525
rect 28460 22488 28488 22519
rect 29822 22516 29828 22528
rect 29880 22516 29886 22568
rect 29932 22556 29960 22610
rect 30929 22593 30941 22627
rect 30975 22624 30987 22627
rect 31846 22624 31852 22636
rect 30975 22596 31852 22624
rect 30975 22593 30987 22596
rect 30929 22587 30987 22593
rect 31846 22584 31852 22596
rect 31904 22624 31910 22636
rect 32214 22624 32220 22636
rect 31904 22596 32220 22624
rect 31904 22584 31910 22596
rect 32214 22584 32220 22596
rect 32272 22584 32278 22636
rect 32582 22624 32588 22636
rect 32543 22596 32588 22624
rect 32582 22584 32588 22596
rect 32640 22584 32646 22636
rect 32876 22633 32904 22732
rect 34054 22720 34060 22732
rect 34112 22720 34118 22772
rect 34238 22720 34244 22772
rect 34296 22760 34302 22772
rect 34606 22760 34612 22772
rect 34296 22732 34612 22760
rect 34296 22720 34302 22732
rect 34606 22720 34612 22732
rect 34664 22720 34670 22772
rect 35161 22763 35219 22769
rect 35161 22729 35173 22763
rect 35207 22760 35219 22763
rect 36262 22760 36268 22772
rect 35207 22732 36268 22760
rect 35207 22729 35219 22732
rect 35161 22723 35219 22729
rect 36262 22720 36268 22732
rect 36320 22760 36326 22772
rect 39482 22760 39488 22772
rect 36320 22732 38654 22760
rect 39443 22732 39488 22760
rect 36320 22720 36326 22732
rect 35713 22695 35771 22701
rect 35713 22692 35725 22695
rect 33704 22664 35725 22692
rect 32861 22627 32919 22633
rect 32861 22593 32873 22627
rect 32907 22593 32919 22627
rect 32861 22587 32919 22593
rect 33704 22556 33732 22664
rect 35713 22661 35725 22664
rect 35759 22661 35771 22695
rect 37182 22692 37188 22704
rect 35713 22655 35771 22661
rect 36142 22664 37188 22692
rect 34149 22627 34207 22633
rect 34149 22593 34161 22627
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34241 22627 34299 22633
rect 34241 22593 34253 22627
rect 34287 22593 34299 22627
rect 34422 22624 34428 22636
rect 34383 22596 34428 22624
rect 34241 22587 34299 22593
rect 29932 22528 33732 22556
rect 29270 22488 29276 22500
rect 28460 22460 29276 22488
rect 29270 22448 29276 22460
rect 29328 22448 29334 22500
rect 30834 22448 30840 22500
rect 30892 22488 30898 22500
rect 33965 22491 34023 22497
rect 33965 22488 33977 22491
rect 30892 22460 33977 22488
rect 30892 22448 30898 22460
rect 33965 22457 33977 22460
rect 34011 22457 34023 22491
rect 33965 22451 34023 22457
rect 30561 22423 30619 22429
rect 30561 22389 30573 22423
rect 30607 22420 30619 22423
rect 31202 22420 31208 22432
rect 30607 22392 31208 22420
rect 30607 22389 30619 22392
rect 30561 22383 30619 22389
rect 31202 22380 31208 22392
rect 31260 22380 31266 22432
rect 31386 22420 31392 22432
rect 31347 22392 31392 22420
rect 31386 22380 31392 22392
rect 31444 22380 31450 22432
rect 33413 22423 33471 22429
rect 33413 22389 33425 22423
rect 33459 22420 33471 22423
rect 33594 22420 33600 22432
rect 33459 22392 33600 22420
rect 33459 22389 33471 22392
rect 33413 22383 33471 22389
rect 33594 22380 33600 22392
rect 33652 22420 33658 22432
rect 33870 22420 33876 22432
rect 33652 22392 33876 22420
rect 33652 22380 33658 22392
rect 33870 22380 33876 22392
rect 33928 22380 33934 22432
rect 34164 22420 34192 22587
rect 34256 22488 34284 22587
rect 34422 22584 34428 22596
rect 34480 22584 34486 22636
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22593 34575 22627
rect 34517 22587 34575 22593
rect 34532 22556 34560 22587
rect 34606 22584 34612 22636
rect 34664 22624 34670 22636
rect 34977 22627 35035 22633
rect 34977 22624 34989 22627
rect 34664 22596 34989 22624
rect 34664 22584 34670 22596
rect 34977 22593 34989 22596
rect 35023 22593 35035 22627
rect 35250 22624 35256 22636
rect 35163 22596 35256 22624
rect 34977 22587 35035 22593
rect 35250 22584 35256 22596
rect 35308 22624 35314 22636
rect 35308 22596 35848 22624
rect 35308 22584 35314 22596
rect 34532 22528 35020 22556
rect 34514 22488 34520 22500
rect 34256 22460 34520 22488
rect 34514 22448 34520 22460
rect 34572 22448 34578 22500
rect 34992 22497 35020 22528
rect 34977 22491 35035 22497
rect 34977 22457 34989 22491
rect 35023 22457 35035 22491
rect 34977 22451 35035 22457
rect 35710 22420 35716 22432
rect 34164 22392 35716 22420
rect 35710 22380 35716 22392
rect 35768 22380 35774 22432
rect 35820 22420 35848 22596
rect 35894 22584 35900 22636
rect 35952 22624 35958 22636
rect 36142 22633 36170 22664
rect 37182 22652 37188 22664
rect 37240 22652 37246 22704
rect 38626 22692 38654 22732
rect 39482 22720 39488 22732
rect 39540 22720 39546 22772
rect 41138 22720 41144 22772
rect 41196 22760 41202 22772
rect 41877 22763 41935 22769
rect 41877 22760 41889 22763
rect 41196 22732 41889 22760
rect 41196 22720 41202 22732
rect 41877 22729 41889 22732
rect 41923 22729 41935 22763
rect 41877 22723 41935 22729
rect 39298 22692 39304 22704
rect 38626 22664 39304 22692
rect 39298 22652 39304 22664
rect 39356 22652 39362 22704
rect 39758 22652 39764 22704
rect 39816 22692 39822 22704
rect 39942 22692 39948 22704
rect 39816 22664 39948 22692
rect 39816 22652 39822 22664
rect 39942 22652 39948 22664
rect 40000 22692 40006 22704
rect 40000 22664 40448 22692
rect 40000 22652 40006 22664
rect 36127 22627 36185 22633
rect 35952 22596 35997 22624
rect 35952 22584 35958 22596
rect 36127 22593 36139 22627
rect 36173 22593 36185 22627
rect 36127 22587 36185 22593
rect 36357 22627 36415 22633
rect 36357 22593 36369 22627
rect 36403 22624 36415 22627
rect 36446 22624 36452 22636
rect 36403 22596 36452 22624
rect 36403 22593 36415 22596
rect 36357 22587 36415 22593
rect 36446 22584 36452 22596
rect 36504 22584 36510 22636
rect 36630 22584 36636 22636
rect 36688 22624 36694 22636
rect 36817 22627 36875 22633
rect 36817 22624 36829 22627
rect 36688 22596 36829 22624
rect 36688 22584 36694 22596
rect 36817 22593 36829 22596
rect 36863 22593 36875 22627
rect 38010 22624 38016 22636
rect 37971 22596 38016 22624
rect 36817 22587 36875 22593
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 38289 22627 38347 22633
rect 38289 22593 38301 22627
rect 38335 22624 38347 22627
rect 38654 22624 38660 22636
rect 38335 22596 38660 22624
rect 38335 22593 38347 22596
rect 38289 22587 38347 22593
rect 38654 22584 38660 22596
rect 38712 22624 38718 22636
rect 39574 22624 39580 22636
rect 38712 22596 39580 22624
rect 38712 22584 38718 22596
rect 39574 22584 39580 22596
rect 39632 22584 39638 22636
rect 40420 22633 40448 22664
rect 40862 22652 40868 22704
rect 40920 22692 40926 22704
rect 41233 22695 41291 22701
rect 41233 22692 41245 22695
rect 40920 22664 41245 22692
rect 40920 22652 40926 22664
rect 41233 22661 41245 22664
rect 41279 22661 41291 22695
rect 42978 22692 42984 22704
rect 41233 22655 41291 22661
rect 41984 22664 42984 22692
rect 40313 22627 40371 22633
rect 40313 22624 40325 22627
rect 39960 22596 40325 22624
rect 39960 22568 39988 22596
rect 40313 22593 40325 22596
rect 40359 22593 40371 22627
rect 40313 22587 40371 22593
rect 40405 22627 40463 22633
rect 40405 22593 40417 22627
rect 40451 22593 40463 22627
rect 41138 22624 41144 22636
rect 41099 22596 41144 22624
rect 40405 22587 40463 22593
rect 41138 22584 41144 22596
rect 41196 22584 41202 22636
rect 41325 22627 41383 22633
rect 41325 22593 41337 22627
rect 41371 22593 41383 22627
rect 41782 22624 41788 22636
rect 41743 22596 41788 22624
rect 41325 22587 41383 22593
rect 35986 22556 35992 22568
rect 35947 22528 35992 22556
rect 35986 22516 35992 22528
rect 36044 22516 36050 22568
rect 36265 22559 36323 22565
rect 36265 22525 36277 22559
rect 36311 22525 36323 22559
rect 36265 22519 36323 22525
rect 36170 22448 36176 22500
rect 36228 22488 36234 22500
rect 36280 22488 36308 22519
rect 37550 22516 37556 22568
rect 37608 22556 37614 22568
rect 37921 22559 37979 22565
rect 37921 22556 37933 22559
rect 37608 22528 37933 22556
rect 37608 22516 37614 22528
rect 37921 22525 37933 22528
rect 37967 22525 37979 22559
rect 37921 22519 37979 22525
rect 38381 22559 38439 22565
rect 38381 22525 38393 22559
rect 38427 22556 38439 22559
rect 38841 22559 38899 22565
rect 38841 22556 38853 22559
rect 38427 22528 38853 22556
rect 38427 22525 38439 22528
rect 38381 22519 38439 22525
rect 38841 22525 38853 22528
rect 38887 22525 38899 22559
rect 39022 22556 39028 22568
rect 38983 22528 39028 22556
rect 38841 22519 38899 22525
rect 39022 22516 39028 22528
rect 39080 22516 39086 22568
rect 39114 22516 39120 22568
rect 39172 22556 39178 22568
rect 39172 22528 39217 22556
rect 39172 22516 39178 22528
rect 39942 22516 39948 22568
rect 40000 22516 40006 22568
rect 40126 22556 40132 22568
rect 40087 22528 40132 22556
rect 40126 22516 40132 22528
rect 40184 22516 40190 22568
rect 40218 22516 40224 22568
rect 40276 22556 40282 22568
rect 40276 22528 40321 22556
rect 40276 22516 40282 22528
rect 39482 22488 39488 22500
rect 36228 22460 36308 22488
rect 36372 22460 39488 22488
rect 36228 22448 36234 22460
rect 36372 22420 36400 22460
rect 39482 22448 39488 22460
rect 39540 22448 39546 22500
rect 40586 22448 40592 22500
rect 40644 22488 40650 22500
rect 41046 22488 41052 22500
rect 40644 22460 41052 22488
rect 40644 22448 40650 22460
rect 41046 22448 41052 22460
rect 41104 22448 41110 22500
rect 41340 22488 41368 22587
rect 41782 22584 41788 22596
rect 41840 22584 41846 22636
rect 41984 22633 42012 22664
rect 42978 22652 42984 22664
rect 43036 22652 43042 22704
rect 43346 22652 43352 22704
rect 43404 22692 43410 22704
rect 57425 22695 57483 22701
rect 57425 22692 57437 22695
rect 43404 22664 57437 22692
rect 43404 22652 43410 22664
rect 57425 22661 57437 22664
rect 57471 22661 57483 22695
rect 57425 22655 57483 22661
rect 41969 22627 42027 22633
rect 41969 22593 41981 22627
rect 42015 22593 42027 22627
rect 41969 22587 42027 22593
rect 42334 22584 42340 22636
rect 42392 22624 42398 22636
rect 42889 22627 42947 22633
rect 42889 22624 42901 22627
rect 42392 22596 42901 22624
rect 42392 22584 42398 22596
rect 42889 22593 42901 22596
rect 42935 22593 42947 22627
rect 42889 22587 42947 22593
rect 43625 22627 43683 22633
rect 43625 22593 43637 22627
rect 43671 22624 43683 22627
rect 44634 22624 44640 22636
rect 43671 22596 44640 22624
rect 43671 22593 43683 22596
rect 43625 22587 43683 22593
rect 41690 22488 41696 22500
rect 41340 22460 41696 22488
rect 41690 22448 41696 22460
rect 41748 22448 41754 22500
rect 41800 22488 41828 22584
rect 42610 22556 42616 22568
rect 42571 22528 42616 22556
rect 42610 22516 42616 22528
rect 42668 22516 42674 22568
rect 42794 22516 42800 22568
rect 42852 22556 42858 22568
rect 43640 22556 43668 22587
rect 44634 22584 44640 22596
rect 44692 22584 44698 22636
rect 45002 22624 45008 22636
rect 44963 22596 45008 22624
rect 45002 22584 45008 22596
rect 45060 22584 45066 22636
rect 45557 22627 45615 22633
rect 45557 22593 45569 22627
rect 45603 22593 45615 22627
rect 45557 22587 45615 22593
rect 42852 22528 43668 22556
rect 42852 22516 42858 22528
rect 44082 22516 44088 22568
rect 44140 22556 44146 22568
rect 44545 22559 44603 22565
rect 44545 22556 44557 22559
rect 44140 22528 44557 22556
rect 44140 22516 44146 22528
rect 44545 22525 44557 22528
rect 44591 22525 44603 22559
rect 44545 22519 44603 22525
rect 45462 22516 45468 22568
rect 45520 22556 45526 22568
rect 45572 22556 45600 22587
rect 45738 22584 45744 22636
rect 45796 22624 45802 22636
rect 46109 22627 46167 22633
rect 46109 22624 46121 22627
rect 45796 22596 46121 22624
rect 45796 22584 45802 22596
rect 46109 22593 46121 22596
rect 46155 22593 46167 22627
rect 57440 22624 57468 22655
rect 58069 22627 58127 22633
rect 58069 22624 58081 22627
rect 57440 22596 58081 22624
rect 46109 22587 46167 22593
rect 58069 22593 58081 22596
rect 58115 22593 58127 22627
rect 58069 22587 58127 22593
rect 46385 22559 46443 22565
rect 46385 22556 46397 22559
rect 45520 22528 46397 22556
rect 45520 22516 45526 22528
rect 46385 22525 46397 22528
rect 46431 22525 46443 22559
rect 46385 22519 46443 22525
rect 42705 22491 42763 22497
rect 42705 22488 42717 22491
rect 41800 22460 42717 22488
rect 42705 22457 42717 22460
rect 42751 22457 42763 22491
rect 42705 22451 42763 22457
rect 45094 22448 45100 22500
rect 45152 22488 45158 22500
rect 45281 22491 45339 22497
rect 45281 22488 45293 22491
rect 45152 22460 45293 22488
rect 45152 22448 45158 22460
rect 45281 22457 45293 22460
rect 45327 22457 45339 22491
rect 58250 22488 58256 22500
rect 58211 22460 58256 22488
rect 45281 22451 45339 22457
rect 58250 22448 58256 22460
rect 58308 22448 58314 22500
rect 35820 22392 36400 22420
rect 37737 22423 37795 22429
rect 37737 22389 37749 22423
rect 37783 22420 37795 22423
rect 38286 22420 38292 22432
rect 37783 22392 38292 22420
rect 37783 22389 37795 22392
rect 37737 22383 37795 22389
rect 38286 22380 38292 22392
rect 38344 22380 38350 22432
rect 39114 22380 39120 22432
rect 39172 22420 39178 22432
rect 39945 22423 40003 22429
rect 39945 22420 39957 22423
rect 39172 22392 39957 22420
rect 39172 22380 39178 22392
rect 39945 22389 39957 22392
rect 39991 22389 40003 22423
rect 43070 22420 43076 22432
rect 43031 22392 43076 22420
rect 39945 22383 40003 22389
rect 43070 22380 43076 22392
rect 43128 22380 43134 22432
rect 43901 22423 43959 22429
rect 43901 22389 43913 22423
rect 43947 22420 43959 22423
rect 43990 22420 43996 22432
rect 43947 22392 43996 22420
rect 43947 22389 43959 22392
rect 43901 22383 43959 22389
rect 43990 22380 43996 22392
rect 44048 22380 44054 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 24854 22176 24860 22228
rect 24912 22216 24918 22228
rect 25041 22219 25099 22225
rect 25041 22216 25053 22219
rect 24912 22188 25053 22216
rect 24912 22176 24918 22188
rect 25041 22185 25053 22188
rect 25087 22185 25099 22219
rect 25041 22179 25099 22185
rect 32582 22176 32588 22228
rect 32640 22216 32646 22228
rect 33042 22216 33048 22228
rect 32640 22188 33048 22216
rect 32640 22176 32646 22188
rect 33042 22176 33048 22188
rect 33100 22216 33106 22228
rect 35069 22219 35127 22225
rect 35069 22216 35081 22219
rect 33100 22188 35081 22216
rect 33100 22176 33106 22188
rect 35069 22185 35081 22188
rect 35115 22216 35127 22219
rect 35986 22216 35992 22228
rect 35115 22188 35992 22216
rect 35115 22185 35127 22188
rect 35069 22179 35127 22185
rect 35986 22176 35992 22188
rect 36044 22176 36050 22228
rect 37734 22216 37740 22228
rect 36096 22188 37740 22216
rect 25869 22151 25927 22157
rect 25869 22117 25881 22151
rect 25915 22148 25927 22151
rect 25958 22148 25964 22160
rect 25915 22120 25964 22148
rect 25915 22117 25927 22120
rect 25869 22111 25927 22117
rect 25958 22108 25964 22120
rect 26016 22108 26022 22160
rect 32953 22151 33011 22157
rect 32953 22117 32965 22151
rect 32999 22148 33011 22151
rect 33410 22148 33416 22160
rect 32999 22120 33416 22148
rect 32999 22117 33011 22120
rect 32953 22111 33011 22117
rect 33410 22108 33416 22120
rect 33468 22108 33474 22160
rect 34606 22108 34612 22160
rect 34664 22148 34670 22160
rect 36096 22148 36124 22188
rect 37734 22176 37740 22188
rect 37792 22176 37798 22228
rect 38010 22176 38016 22228
rect 38068 22216 38074 22228
rect 38197 22219 38255 22225
rect 38197 22216 38209 22219
rect 38068 22188 38209 22216
rect 38068 22176 38074 22188
rect 38197 22185 38209 22188
rect 38243 22185 38255 22219
rect 38197 22179 38255 22185
rect 38608 22176 38614 22228
rect 38666 22176 38672 22228
rect 39482 22176 39488 22228
rect 39540 22216 39546 22228
rect 42889 22219 42947 22225
rect 42889 22216 42901 22219
rect 39540 22188 42901 22216
rect 39540 22176 39546 22188
rect 42889 22185 42901 22188
rect 42935 22185 42947 22219
rect 42889 22179 42947 22185
rect 43162 22176 43168 22228
rect 43220 22216 43226 22228
rect 44177 22219 44235 22225
rect 44177 22216 44189 22219
rect 43220 22188 44189 22216
rect 43220 22176 43226 22188
rect 44177 22185 44189 22188
rect 44223 22185 44235 22219
rect 44177 22179 44235 22185
rect 34664 22120 36124 22148
rect 34664 22108 34670 22120
rect 36170 22108 36176 22160
rect 36228 22108 36234 22160
rect 38378 22108 38384 22160
rect 38436 22148 38442 22160
rect 38626 22148 38654 22176
rect 41690 22148 41696 22160
rect 38436 22120 38516 22148
rect 38626 22120 41696 22148
rect 38436 22108 38442 22120
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 22888 22052 23612 22080
rect 22888 22040 22894 22052
rect 21726 21972 21732 22024
rect 21784 21972 21790 22024
rect 22189 22015 22247 22021
rect 22189 21981 22201 22015
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 1946 21904 1952 21956
rect 2004 21944 2010 21956
rect 21177 21947 21235 21953
rect 21177 21944 21189 21947
rect 2004 21916 21189 21944
rect 2004 21904 2010 21916
rect 21177 21913 21189 21916
rect 21223 21913 21235 21947
rect 22204 21944 22232 21975
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22336 21984 23520 22012
rect 22336 21972 22342 21984
rect 23382 21944 23388 21956
rect 22204 21916 23388 21944
rect 21177 21907 21235 21913
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 23492 21888 23520 21984
rect 23290 21876 23296 21888
rect 23251 21848 23296 21876
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 23474 21876 23480 21888
rect 23435 21848 23480 21876
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23584 21885 23612 22052
rect 25682 22040 25688 22092
rect 25740 22080 25746 22092
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 25740 22052 26525 22080
rect 25740 22040 25746 22052
rect 26513 22049 26525 22052
rect 26559 22049 26571 22083
rect 26970 22080 26976 22092
rect 26931 22052 26976 22080
rect 26513 22043 26571 22049
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 29270 22040 29276 22092
rect 29328 22080 29334 22092
rect 32677 22083 32735 22089
rect 32677 22080 32689 22083
rect 29328 22052 32689 22080
rect 29328 22040 29334 22052
rect 32677 22049 32689 22052
rect 32723 22049 32735 22083
rect 32677 22043 32735 22049
rect 33045 22083 33103 22089
rect 33045 22049 33057 22083
rect 33091 22080 33103 22083
rect 33226 22080 33232 22092
rect 33091 22052 33232 22080
rect 33091 22049 33103 22052
rect 33045 22043 33103 22049
rect 33226 22040 33232 22052
rect 33284 22040 33290 22092
rect 35434 22080 35440 22092
rect 33888 22052 35440 22080
rect 25133 22015 25191 22021
rect 25133 21981 25145 22015
rect 25179 21981 25191 22015
rect 25590 22012 25596 22024
rect 25551 21984 25596 22012
rect 25133 21975 25191 21981
rect 23750 21944 23756 21956
rect 23711 21916 23756 21944
rect 23750 21904 23756 21916
rect 23808 21904 23814 21956
rect 25148 21944 25176 21975
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 25774 22012 25780 22024
rect 25735 21984 25780 22012
rect 25774 21972 25780 21984
rect 25832 21972 25838 22024
rect 26881 22015 26939 22021
rect 26881 21981 26893 22015
rect 26927 22012 26939 22015
rect 27154 22012 27160 22024
rect 26927 21984 27160 22012
rect 26927 21981 26939 21984
rect 26881 21975 26939 21981
rect 27154 21972 27160 21984
rect 27212 21972 27218 22024
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30650 22012 30656 22024
rect 30607 21984 30656 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 30650 21972 30656 21984
rect 30708 21972 30714 22024
rect 30837 22015 30895 22021
rect 30837 21981 30849 22015
rect 30883 22012 30895 22015
rect 31018 22012 31024 22024
rect 30883 21984 31024 22012
rect 30883 21981 30895 21984
rect 30837 21975 30895 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 31478 22012 31484 22024
rect 31439 21984 31484 22012
rect 31478 21972 31484 21984
rect 31536 21972 31542 22024
rect 31573 22015 31631 22021
rect 31573 21981 31585 22015
rect 31619 21981 31631 22015
rect 31573 21975 31631 21981
rect 31665 22015 31723 22021
rect 31665 21981 31677 22015
rect 31711 21981 31723 22015
rect 31665 21975 31723 21981
rect 31757 22015 31815 22021
rect 31757 21981 31769 22015
rect 31803 22012 31815 22015
rect 31846 22012 31852 22024
rect 31803 21984 31852 22012
rect 31803 21981 31815 21984
rect 31757 21975 31815 21981
rect 26510 21944 26516 21956
rect 25148 21916 26516 21944
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21845 23627 21879
rect 23569 21839 23627 21845
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 30524 21848 31309 21876
rect 30524 21836 30530 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 31588 21876 31616 21975
rect 31680 21944 31708 21975
rect 31846 21972 31852 21984
rect 31904 21972 31910 22024
rect 32829 22015 32887 22021
rect 32829 22012 32841 22015
rect 32600 21984 32841 22012
rect 32600 21956 32628 21984
rect 32829 21981 32841 21984
rect 32875 21981 32887 22015
rect 32829 21975 32887 21981
rect 33134 21972 33140 22024
rect 33192 22012 33198 22024
rect 33192 21984 33237 22012
rect 33192 21972 33198 21984
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 33888 22021 33916 22052
rect 35434 22040 35440 22052
rect 35492 22040 35498 22092
rect 35710 22080 35716 22092
rect 35671 22052 35716 22080
rect 35710 22040 35716 22052
rect 35768 22040 35774 22092
rect 36188 22080 36216 22108
rect 35912 22052 36216 22080
rect 33873 22015 33931 22021
rect 33873 22012 33885 22015
rect 33376 21984 33885 22012
rect 33376 21972 33382 21984
rect 33873 21981 33885 21984
rect 33919 21981 33931 22015
rect 33873 21975 33931 21981
rect 34057 22015 34115 22021
rect 34057 21981 34069 22015
rect 34103 22012 34115 22015
rect 34698 22012 34704 22024
rect 34103 21984 34704 22012
rect 34103 21981 34115 21984
rect 34057 21975 34115 21981
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 34885 22015 34943 22021
rect 34885 21981 34897 22015
rect 34931 22012 34943 22015
rect 35066 22012 35072 22024
rect 34931 21984 35072 22012
rect 34931 21981 34943 21984
rect 34885 21975 34943 21981
rect 32582 21944 32588 21956
rect 31680 21916 32588 21944
rect 32582 21904 32588 21916
rect 32640 21904 32646 21956
rect 33336 21944 33364 21972
rect 33152 21916 33364 21944
rect 33152 21876 33180 21916
rect 34514 21904 34520 21956
rect 34572 21944 34578 21956
rect 34900 21944 34928 21975
rect 35066 21972 35072 21984
rect 35124 21972 35130 22024
rect 35912 22021 35940 22052
rect 36446 22040 36452 22092
rect 36504 22080 36510 22092
rect 36725 22083 36783 22089
rect 36725 22080 36737 22083
rect 36504 22052 36737 22080
rect 36504 22040 36510 22052
rect 36725 22049 36737 22052
rect 36771 22080 36783 22083
rect 36998 22080 37004 22092
rect 36771 22052 37004 22080
rect 36771 22049 36783 22052
rect 36725 22043 36783 22049
rect 36998 22040 37004 22052
rect 37056 22040 37062 22092
rect 38488 22089 38516 22120
rect 41690 22108 41696 22120
rect 41748 22108 41754 22160
rect 41782 22108 41788 22160
rect 41840 22148 41846 22160
rect 45922 22148 45928 22160
rect 41840 22120 45928 22148
rect 41840 22108 41846 22120
rect 45922 22108 45928 22120
rect 45980 22108 45986 22160
rect 38473 22083 38531 22089
rect 38473 22049 38485 22083
rect 38519 22049 38531 22083
rect 38473 22043 38531 22049
rect 38654 22040 38660 22092
rect 38712 22080 38718 22092
rect 39298 22080 39304 22092
rect 38712 22052 39160 22080
rect 39259 22052 39304 22080
rect 38712 22040 38718 22052
rect 35897 22015 35955 22021
rect 35897 21981 35909 22015
rect 35943 21981 35955 22015
rect 35897 21975 35955 21981
rect 35989 22015 36047 22021
rect 35989 21981 36001 22015
rect 36035 21981 36047 22015
rect 35989 21975 36047 21981
rect 36117 22015 36175 22021
rect 36117 21981 36129 22015
rect 36163 22012 36175 22015
rect 36814 22012 36820 22024
rect 36163 21984 36820 22012
rect 36163 21981 36175 21984
rect 36117 21975 36175 21981
rect 34572 21916 34928 21944
rect 36004 21944 36032 21975
rect 36814 21972 36820 21984
rect 36872 21972 36878 22024
rect 37369 22015 37427 22021
rect 37369 21981 37381 22015
rect 37415 22012 37427 22015
rect 38010 22012 38016 22024
rect 37415 21984 38016 22012
rect 37415 21981 37427 21984
rect 37369 21975 37427 21981
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 38194 21972 38200 22024
rect 38252 22012 38258 22024
rect 38381 22015 38439 22021
rect 38381 22012 38393 22015
rect 38252 21984 38393 22012
rect 38252 21972 38258 21984
rect 38381 21981 38393 21984
rect 38427 21981 38439 22015
rect 38381 21975 38439 21981
rect 38565 22015 38623 22021
rect 38565 21981 38577 22015
rect 38611 21981 38623 22015
rect 39132 22012 39160 22052
rect 39298 22040 39304 22052
rect 39356 22040 39362 22092
rect 39942 22040 39948 22092
rect 40000 22080 40006 22092
rect 40681 22083 40739 22089
rect 40681 22080 40693 22083
rect 40000 22052 40693 22080
rect 40000 22040 40006 22052
rect 40681 22049 40693 22052
rect 40727 22049 40739 22083
rect 40681 22043 40739 22049
rect 40954 22040 40960 22092
rect 41012 22080 41018 22092
rect 41012 22052 41920 22080
rect 41012 22040 41018 22052
rect 39758 22012 39764 22024
rect 39132 21984 39764 22012
rect 38565 21975 38623 21981
rect 36262 21944 36268 21956
rect 36004 21916 36268 21944
rect 34572 21904 34578 21916
rect 36262 21904 36268 21916
rect 36320 21904 36326 21956
rect 36722 21904 36728 21956
rect 36780 21944 36786 21956
rect 37185 21947 37243 21953
rect 37185 21944 37197 21947
rect 36780 21916 37197 21944
rect 36780 21904 36786 21916
rect 37185 21913 37197 21916
rect 37231 21913 37243 21947
rect 37734 21944 37740 21956
rect 37695 21916 37740 21944
rect 37185 21907 37243 21913
rect 37734 21904 37740 21916
rect 37792 21904 37798 21956
rect 38581 21944 38609 21975
rect 39758 21972 39764 21984
rect 39816 21972 39822 22024
rect 40034 22012 40040 22024
rect 39995 21984 40040 22012
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 40218 21972 40224 22024
rect 40276 22012 40282 22024
rect 40276 21984 40321 22012
rect 40276 21972 40282 21984
rect 41138 21972 41144 22024
rect 41196 22012 41202 22024
rect 41892 22012 41920 22052
rect 41966 22040 41972 22092
rect 42024 22080 42030 22092
rect 42337 22083 42395 22089
rect 42337 22080 42349 22083
rect 42024 22052 42349 22080
rect 42024 22040 42030 22052
rect 42337 22049 42349 22052
rect 42383 22049 42395 22083
rect 43622 22080 43628 22092
rect 42337 22043 42395 22049
rect 43364 22052 43628 22080
rect 43364 22024 43392 22052
rect 43622 22040 43628 22052
rect 43680 22040 43686 22092
rect 45738 22080 45744 22092
rect 44376 22052 45744 22080
rect 42794 22012 42800 22024
rect 41196 21984 41736 22012
rect 41196 21972 41202 21984
rect 40310 21944 40316 21956
rect 38581 21916 40316 21944
rect 31588 21848 33180 21876
rect 31297 21839 31355 21845
rect 33226 21836 33232 21888
rect 33284 21876 33290 21888
rect 33689 21879 33747 21885
rect 33689 21876 33701 21879
rect 33284 21848 33701 21876
rect 33284 21836 33290 21848
rect 33689 21845 33701 21848
rect 33735 21876 33747 21879
rect 33870 21876 33876 21888
rect 33735 21848 33876 21876
rect 33735 21845 33747 21848
rect 33689 21839 33747 21845
rect 33870 21836 33876 21848
rect 33928 21836 33934 21888
rect 35526 21836 35532 21888
rect 35584 21876 35590 21888
rect 35802 21876 35808 21888
rect 35584 21848 35808 21876
rect 35584 21836 35590 21848
rect 35802 21836 35808 21848
rect 35860 21876 35866 21888
rect 36446 21876 36452 21888
rect 35860 21848 36452 21876
rect 35860 21836 35866 21848
rect 36446 21836 36452 21848
rect 36504 21836 36510 21888
rect 37366 21836 37372 21888
rect 37424 21876 37430 21888
rect 38581 21876 38609 21916
rect 40310 21904 40316 21916
rect 40368 21944 40374 21956
rect 40954 21944 40960 21956
rect 40368 21916 40960 21944
rect 40368 21904 40374 21916
rect 40954 21904 40960 21916
rect 41012 21904 41018 21956
rect 37424 21848 38609 21876
rect 37424 21836 37430 21848
rect 39022 21836 39028 21888
rect 39080 21876 39086 21888
rect 39850 21876 39856 21888
rect 39080 21848 39856 21876
rect 39080 21836 39086 21848
rect 39850 21836 39856 21848
rect 39908 21876 39914 21888
rect 40037 21879 40095 21885
rect 40037 21876 40049 21879
rect 39908 21848 40049 21876
rect 39908 21836 39914 21848
rect 40037 21845 40049 21848
rect 40083 21845 40095 21879
rect 40037 21839 40095 21845
rect 40126 21836 40132 21888
rect 40184 21876 40190 21888
rect 41230 21876 41236 21888
rect 40184 21848 41236 21876
rect 40184 21836 40190 21848
rect 41230 21836 41236 21848
rect 41288 21836 41294 21888
rect 41708 21876 41736 21984
rect 41892 21984 42800 22012
rect 41892 21944 41920 21984
rect 42794 21972 42800 21984
rect 42852 21972 42858 22024
rect 43165 22015 43223 22021
rect 43076 21993 43134 21999
rect 43076 21959 43088 21993
rect 43122 21959 43134 21993
rect 43165 21981 43177 22015
rect 43211 21981 43223 22015
rect 43346 22012 43352 22024
rect 43307 21984 43352 22012
rect 43165 21975 43223 21981
rect 43076 21956 43134 21959
rect 42061 21947 42119 21953
rect 42061 21944 42073 21947
rect 41892 21916 42073 21944
rect 42061 21913 42073 21916
rect 42107 21913 42119 21947
rect 42061 21907 42119 21913
rect 43070 21904 43076 21956
rect 43128 21904 43134 21956
rect 43180 21944 43208 21975
rect 43346 21972 43352 21984
rect 43404 21972 43410 22024
rect 43441 22015 43499 22021
rect 43441 21981 43453 22015
rect 43487 22012 43499 22015
rect 43990 22012 43996 22024
rect 43487 21984 43996 22012
rect 43487 21981 43499 21984
rect 43441 21975 43499 21981
rect 43990 21972 43996 21984
rect 44048 21972 44054 22024
rect 44085 22015 44143 22021
rect 44085 21981 44097 22015
rect 44131 21981 44143 22015
rect 44085 21975 44143 21981
rect 44177 22015 44235 22021
rect 44177 21981 44189 22015
rect 44223 22012 44235 22015
rect 44266 22012 44272 22024
rect 44223 21984 44272 22012
rect 44223 21981 44235 21984
rect 44177 21975 44235 21981
rect 43714 21944 43720 21956
rect 43180 21916 43720 21944
rect 43714 21904 43720 21916
rect 43772 21904 43778 21956
rect 44100 21944 44128 21975
rect 44266 21972 44272 21984
rect 44324 22012 44330 22024
rect 44376 22012 44404 22052
rect 45738 22040 45744 22052
rect 45796 22040 45802 22092
rect 45370 22012 45376 22024
rect 44324 21984 44417 22012
rect 45331 21984 45376 22012
rect 44324 21978 44404 21984
rect 44324 21972 44330 21978
rect 45370 21972 45376 21984
rect 45428 21972 45434 22024
rect 45462 21972 45468 22024
rect 45520 22012 45526 22024
rect 45649 22015 45707 22021
rect 45649 22012 45661 22015
rect 45520 21984 45661 22012
rect 45520 21972 45526 21984
rect 45649 21981 45661 21984
rect 45695 21981 45707 22015
rect 45830 22012 45836 22024
rect 45791 21984 45836 22012
rect 45649 21975 45707 21981
rect 45830 21972 45836 21984
rect 45888 21972 45894 22024
rect 44450 21944 44456 21956
rect 44100 21916 44456 21944
rect 44450 21904 44456 21916
rect 44508 21944 44514 21956
rect 45388 21944 45416 21972
rect 44508 21916 45416 21944
rect 44508 21904 44514 21916
rect 45189 21879 45247 21885
rect 45189 21876 45201 21879
rect 41708 21848 45201 21876
rect 45189 21845 45201 21848
rect 45235 21845 45247 21879
rect 45189 21839 45247 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 23658 21672 23664 21684
rect 23619 21644 23664 21672
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 23750 21632 23756 21684
rect 23808 21672 23814 21684
rect 25501 21675 25559 21681
rect 23808 21644 23853 21672
rect 23808 21632 23814 21644
rect 25501 21641 25513 21675
rect 25547 21672 25559 21675
rect 25590 21672 25596 21684
rect 25547 21644 25596 21672
rect 25547 21641 25559 21644
rect 25501 21635 25559 21641
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 28166 21672 28172 21684
rect 27948 21644 28172 21672
rect 27948 21632 27954 21644
rect 28166 21632 28172 21644
rect 28224 21672 28230 21684
rect 28997 21675 29055 21681
rect 28997 21672 29009 21675
rect 28224 21644 29009 21672
rect 28224 21632 28230 21644
rect 28997 21641 29009 21644
rect 29043 21672 29055 21675
rect 30193 21675 30251 21681
rect 30193 21672 30205 21675
rect 29043 21644 30205 21672
rect 29043 21641 29055 21644
rect 28997 21635 29055 21641
rect 30193 21641 30205 21644
rect 30239 21641 30251 21675
rect 31018 21672 31024 21684
rect 30979 21644 31024 21672
rect 30193 21635 30251 21641
rect 31018 21632 31024 21644
rect 31076 21632 31082 21684
rect 32401 21675 32459 21681
rect 32401 21641 32413 21675
rect 32447 21672 32459 21675
rect 33318 21672 33324 21684
rect 32447 21644 33324 21672
rect 32447 21641 32459 21644
rect 32401 21635 32459 21641
rect 33318 21632 33324 21644
rect 33376 21632 33382 21684
rect 34054 21632 34060 21684
rect 34112 21672 34118 21684
rect 34517 21675 34575 21681
rect 34517 21672 34529 21675
rect 34112 21644 34529 21672
rect 34112 21632 34118 21644
rect 34517 21641 34529 21644
rect 34563 21641 34575 21675
rect 34517 21635 34575 21641
rect 34698 21632 34704 21684
rect 34756 21672 34762 21684
rect 35434 21672 35440 21684
rect 34756 21644 35440 21672
rect 34756 21632 34762 21644
rect 35434 21632 35440 21644
rect 35492 21632 35498 21684
rect 35713 21675 35771 21681
rect 35713 21641 35725 21675
rect 35759 21672 35771 21675
rect 36170 21672 36176 21684
rect 35759 21644 36176 21672
rect 35759 21641 35771 21644
rect 35713 21635 35771 21641
rect 36170 21632 36176 21644
rect 36228 21632 36234 21684
rect 36814 21632 36820 21684
rect 36872 21672 36878 21684
rect 37550 21672 37556 21684
rect 36872 21644 37556 21672
rect 36872 21632 36878 21644
rect 37550 21632 37556 21644
rect 37608 21672 37614 21684
rect 37826 21672 37832 21684
rect 37608 21644 37832 21672
rect 37608 21632 37614 21644
rect 37826 21632 37832 21644
rect 37884 21632 37890 21684
rect 38194 21632 38200 21684
rect 38252 21672 38258 21684
rect 39298 21672 39304 21684
rect 38252 21644 39304 21672
rect 38252 21632 38258 21644
rect 39298 21632 39304 21644
rect 39356 21632 39362 21684
rect 44818 21672 44824 21684
rect 44779 21644 44824 21672
rect 44818 21632 44824 21644
rect 44876 21632 44882 21684
rect 45830 21672 45836 21684
rect 45204 21644 45836 21672
rect 23290 21564 23296 21616
rect 23348 21604 23354 21616
rect 23934 21604 23940 21616
rect 23348 21576 23940 21604
rect 23348 21564 23354 21576
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 29822 21604 29828 21616
rect 29104 21576 29828 21604
rect 23474 21536 23480 21548
rect 22954 21508 23480 21536
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23842 21536 23848 21548
rect 23615 21508 23848 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 25682 21536 25688 21548
rect 25643 21508 25688 21536
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 27893 21539 27951 21545
rect 27893 21505 27905 21539
rect 27939 21536 27951 21539
rect 28350 21536 28356 21548
rect 27939 21508 28356 21536
rect 27939 21505 27951 21508
rect 27893 21499 27951 21505
rect 28350 21496 28356 21508
rect 28408 21496 28414 21548
rect 29104 21480 29132 21576
rect 29822 21564 29828 21576
rect 29880 21604 29886 21616
rect 30285 21607 30343 21613
rect 30285 21604 30297 21607
rect 29880 21576 30297 21604
rect 29880 21564 29886 21576
rect 30285 21573 30297 21576
rect 30331 21573 30343 21607
rect 32582 21604 32588 21616
rect 32543 21576 32588 21604
rect 30285 21567 30343 21573
rect 32582 21564 32588 21576
rect 32640 21564 32646 21616
rect 33873 21607 33931 21613
rect 33873 21573 33885 21607
rect 33919 21604 33931 21607
rect 34977 21607 35035 21613
rect 34977 21604 34989 21607
rect 33919 21576 34989 21604
rect 33919 21573 33931 21576
rect 33873 21567 33931 21573
rect 34532 21548 34560 21576
rect 34977 21573 34989 21576
rect 35023 21573 35035 21607
rect 34977 21567 35035 21573
rect 35066 21564 35072 21616
rect 35124 21604 35130 21616
rect 36078 21604 36084 21616
rect 35124 21576 36084 21604
rect 35124 21564 35130 21576
rect 36078 21564 36084 21576
rect 36136 21564 36142 21616
rect 36630 21604 36636 21616
rect 36188 21576 36636 21604
rect 31202 21536 31208 21548
rect 31163 21508 31208 21536
rect 31202 21496 31208 21508
rect 31260 21496 31266 21548
rect 31389 21539 31447 21545
rect 31389 21505 31401 21539
rect 31435 21505 31447 21539
rect 31389 21499 31447 21505
rect 22097 21471 22155 21477
rect 22097 21437 22109 21471
rect 22143 21468 22155 21471
rect 22186 21468 22192 21480
rect 22143 21440 22192 21468
rect 22143 21437 22155 21440
rect 22097 21431 22155 21437
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 22830 21468 22836 21480
rect 22791 21440 22836 21468
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 23750 21428 23756 21480
rect 23808 21468 23814 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23808 21440 24041 21468
rect 23808 21428 23814 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 25961 21471 26019 21477
rect 25961 21437 25973 21471
rect 26007 21468 26019 21471
rect 26050 21468 26056 21480
rect 26007 21440 26056 21468
rect 26007 21437 26019 21440
rect 25961 21431 26019 21437
rect 26050 21428 26056 21440
rect 26108 21428 26114 21480
rect 29086 21468 29092 21480
rect 29047 21440 29092 21468
rect 29086 21428 29092 21440
rect 29144 21428 29150 21480
rect 29273 21471 29331 21477
rect 29273 21437 29285 21471
rect 29319 21437 29331 21471
rect 30466 21468 30472 21480
rect 30427 21440 30472 21468
rect 29273 21431 29331 21437
rect 25038 21360 25044 21412
rect 25096 21400 25102 21412
rect 29288 21400 29316 21431
rect 30466 21428 30472 21440
rect 30524 21428 30530 21480
rect 31404 21468 31432 21499
rect 31478 21496 31484 21548
rect 31536 21536 31542 21548
rect 32214 21536 32220 21548
rect 31536 21508 32220 21536
rect 31536 21496 31542 21508
rect 32214 21496 32220 21508
rect 32272 21536 32278 21548
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 32272 21508 32321 21536
rect 32272 21496 32278 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 32398 21496 32404 21548
rect 32456 21536 32462 21548
rect 33781 21539 33839 21545
rect 33781 21536 33793 21539
rect 32456 21508 33793 21536
rect 32456 21496 32462 21508
rect 33781 21505 33793 21508
rect 33827 21505 33839 21539
rect 33962 21536 33968 21548
rect 33923 21508 33968 21536
rect 33781 21499 33839 21505
rect 32766 21468 32772 21480
rect 31404 21440 32772 21468
rect 32766 21428 32772 21440
rect 32824 21428 32830 21480
rect 33796 21468 33824 21499
rect 33962 21496 33968 21508
rect 34020 21496 34026 21548
rect 34514 21496 34520 21548
rect 34572 21496 34578 21548
rect 34698 21536 34704 21548
rect 34659 21508 34704 21536
rect 34698 21496 34704 21508
rect 34756 21496 34762 21548
rect 34793 21539 34851 21545
rect 34793 21505 34805 21539
rect 34839 21536 34851 21539
rect 35434 21536 35440 21548
rect 34839 21508 35440 21536
rect 34839 21505 34851 21508
rect 34793 21499 34851 21505
rect 35434 21496 35440 21508
rect 35492 21496 35498 21548
rect 35529 21539 35587 21545
rect 35529 21505 35541 21539
rect 35575 21536 35587 21539
rect 35618 21536 35624 21548
rect 35575 21508 35624 21536
rect 35575 21505 35587 21508
rect 35529 21499 35587 21505
rect 35618 21496 35624 21508
rect 35676 21496 35682 21548
rect 35710 21496 35716 21548
rect 35768 21536 35774 21548
rect 36188 21545 36216 21576
rect 36630 21564 36636 21576
rect 36688 21564 36694 21616
rect 36998 21564 37004 21616
rect 37056 21604 37062 21616
rect 37056 21576 38976 21604
rect 37056 21564 37062 21576
rect 36173 21539 36231 21545
rect 35768 21508 35813 21536
rect 35768 21496 35774 21508
rect 36173 21505 36185 21539
rect 36219 21505 36231 21539
rect 36173 21499 36231 21505
rect 36265 21539 36323 21545
rect 36265 21505 36277 21539
rect 36311 21536 36323 21539
rect 37182 21536 37188 21548
rect 36311 21508 37188 21536
rect 36311 21505 36323 21508
rect 36265 21499 36323 21505
rect 37182 21496 37188 21508
rect 37240 21536 37246 21548
rect 37553 21539 37611 21545
rect 37240 21508 37504 21536
rect 37240 21496 37246 21508
rect 36449 21471 36507 21477
rect 33796 21440 36032 21468
rect 36004 21412 36032 21440
rect 36449 21437 36461 21471
rect 36495 21468 36507 21471
rect 37274 21468 37280 21480
rect 36495 21440 37280 21468
rect 36495 21437 36507 21440
rect 36449 21431 36507 21437
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 37476 21468 37504 21508
rect 37553 21505 37565 21539
rect 37599 21536 37611 21539
rect 37642 21536 37648 21548
rect 37599 21508 37648 21536
rect 37599 21505 37611 21508
rect 37553 21499 37611 21505
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 37737 21539 37795 21545
rect 37737 21505 37749 21539
rect 37783 21536 37795 21539
rect 38194 21536 38200 21548
rect 37783 21508 38200 21536
rect 37783 21505 37795 21508
rect 37737 21499 37795 21505
rect 38194 21496 38200 21508
rect 38252 21496 38258 21548
rect 38562 21536 38568 21548
rect 38523 21508 38568 21536
rect 38562 21496 38568 21508
rect 38620 21496 38626 21548
rect 38749 21539 38807 21545
rect 38749 21505 38761 21539
rect 38795 21536 38807 21539
rect 38838 21536 38844 21548
rect 38795 21508 38844 21536
rect 38795 21505 38807 21508
rect 38749 21499 38807 21505
rect 38838 21496 38844 21508
rect 38896 21496 38902 21548
rect 38948 21536 38976 21576
rect 39758 21564 39764 21616
rect 39816 21604 39822 21616
rect 41966 21604 41972 21616
rect 39816 21576 41972 21604
rect 39816 21564 39822 21576
rect 39206 21536 39212 21548
rect 38948 21508 39212 21536
rect 39206 21496 39212 21508
rect 39264 21496 39270 21548
rect 39577 21539 39635 21545
rect 39577 21505 39589 21539
rect 39623 21505 39635 21539
rect 39850 21536 39856 21548
rect 39811 21508 39856 21536
rect 39577 21499 39635 21505
rect 37918 21468 37924 21480
rect 37476 21440 37924 21468
rect 37918 21428 37924 21440
rect 37976 21428 37982 21480
rect 38470 21428 38476 21480
rect 38528 21468 38534 21480
rect 39482 21468 39488 21480
rect 38528 21440 39488 21468
rect 38528 21428 38534 21440
rect 39482 21428 39488 21440
rect 39540 21468 39546 21480
rect 39592 21468 39620 21499
rect 39850 21496 39856 21508
rect 39908 21496 39914 21548
rect 40402 21496 40408 21548
rect 40460 21536 40466 21548
rect 40788 21545 40816 21576
rect 41966 21564 41972 21576
rect 42024 21564 42030 21616
rect 42061 21607 42119 21613
rect 42061 21573 42073 21607
rect 42107 21604 42119 21607
rect 42705 21607 42763 21613
rect 42705 21604 42717 21607
rect 42107 21576 42717 21604
rect 42107 21573 42119 21576
rect 42061 21567 42119 21573
rect 42705 21573 42717 21576
rect 42751 21604 42763 21607
rect 43530 21604 43536 21616
rect 42751 21576 43536 21604
rect 42751 21573 42763 21576
rect 42705 21567 42763 21573
rect 43530 21564 43536 21576
rect 43588 21564 43594 21616
rect 44082 21564 44088 21616
rect 44140 21604 44146 21616
rect 45204 21604 45232 21644
rect 45830 21632 45836 21644
rect 45888 21632 45894 21684
rect 45922 21632 45928 21684
rect 45980 21672 45986 21684
rect 45980 21644 46025 21672
rect 45980 21632 45986 21644
rect 45462 21604 45468 21616
rect 44140 21576 45232 21604
rect 45296 21576 45468 21604
rect 44140 21564 44146 21576
rect 40589 21539 40647 21545
rect 40589 21536 40601 21539
rect 40460 21508 40601 21536
rect 40460 21496 40466 21508
rect 40589 21505 40601 21508
rect 40635 21505 40647 21539
rect 40589 21499 40647 21505
rect 40773 21539 40831 21545
rect 40773 21505 40785 21539
rect 40819 21505 40831 21539
rect 40773 21499 40831 21505
rect 40862 21496 40868 21548
rect 40920 21536 40926 21548
rect 41049 21539 41107 21545
rect 40920 21508 40965 21536
rect 40920 21496 40926 21508
rect 41049 21505 41061 21539
rect 41095 21536 41107 21539
rect 41322 21536 41328 21548
rect 41095 21508 41328 21536
rect 41095 21505 41107 21508
rect 41049 21499 41107 21505
rect 41322 21496 41328 21508
rect 41380 21496 41386 21548
rect 43254 21496 43260 21548
rect 43312 21536 43318 21548
rect 43625 21539 43683 21545
rect 43625 21536 43637 21539
rect 43312 21508 43637 21536
rect 43312 21496 43318 21508
rect 43625 21505 43637 21508
rect 43671 21536 43683 21539
rect 43806 21536 43812 21548
rect 43671 21508 43812 21536
rect 43671 21505 43683 21508
rect 43625 21499 43683 21505
rect 43806 21496 43812 21508
rect 43864 21496 43870 21548
rect 43901 21539 43959 21545
rect 43901 21505 43913 21539
rect 43947 21536 43959 21539
rect 44174 21536 44180 21548
rect 43947 21508 44180 21536
rect 43947 21505 43959 21508
rect 43901 21499 43959 21505
rect 44174 21496 44180 21508
rect 44232 21536 44238 21548
rect 44450 21536 44456 21548
rect 44232 21508 44456 21536
rect 44232 21496 44238 21508
rect 44450 21496 44456 21508
rect 44508 21496 44514 21548
rect 44652 21545 44680 21576
rect 45296 21548 45324 21576
rect 45462 21564 45468 21576
rect 45520 21604 45526 21616
rect 45520 21576 46520 21604
rect 45520 21564 45526 21576
rect 44637 21539 44695 21545
rect 44637 21505 44649 21539
rect 44683 21505 44695 21539
rect 45002 21536 45008 21548
rect 44963 21508 45008 21536
rect 44637 21499 44695 21505
rect 45002 21496 45008 21508
rect 45060 21496 45066 21548
rect 45278 21536 45284 21548
rect 45239 21508 45284 21536
rect 45278 21496 45284 21508
rect 45336 21496 45342 21548
rect 46492 21545 46520 21576
rect 45741 21539 45799 21545
rect 45741 21505 45753 21539
rect 45787 21505 45799 21539
rect 45741 21499 45799 21505
rect 46477 21539 46535 21545
rect 46477 21505 46489 21539
rect 46523 21505 46535 21539
rect 46477 21499 46535 21505
rect 39540 21440 39620 21468
rect 39669 21471 39727 21477
rect 39540 21428 39546 21440
rect 39669 21437 39681 21471
rect 39715 21468 39727 21471
rect 40494 21468 40500 21480
rect 39715 21440 40500 21468
rect 39715 21437 39727 21440
rect 39669 21431 39727 21437
rect 40494 21428 40500 21440
rect 40552 21428 40558 21480
rect 40880 21468 40908 21496
rect 43533 21471 43591 21477
rect 43533 21468 43545 21471
rect 40880 21440 43545 21468
rect 43533 21437 43545 21440
rect 43579 21468 43591 21471
rect 43579 21440 43668 21468
rect 43579 21437 43591 21440
rect 43533 21431 43591 21437
rect 43640 21412 43668 21440
rect 43714 21428 43720 21480
rect 43772 21468 43778 21480
rect 44082 21468 44088 21480
rect 43772 21440 44088 21468
rect 43772 21428 43778 21440
rect 44082 21428 44088 21440
rect 44140 21428 44146 21480
rect 45756 21468 45784 21499
rect 45020 21440 45784 21468
rect 31846 21400 31852 21412
rect 25096 21372 29040 21400
rect 29288 21372 31852 21400
rect 25096 21360 25102 21372
rect 25869 21335 25927 21341
rect 25869 21301 25881 21335
rect 25915 21332 25927 21335
rect 25958 21332 25964 21344
rect 25915 21304 25964 21332
rect 25915 21301 25927 21304
rect 25869 21295 25927 21301
rect 25958 21292 25964 21304
rect 26016 21292 26022 21344
rect 27890 21292 27896 21344
rect 27948 21332 27954 21344
rect 28077 21335 28135 21341
rect 28077 21332 28089 21335
rect 27948 21304 28089 21332
rect 27948 21292 27954 21304
rect 28077 21301 28089 21304
rect 28123 21301 28135 21335
rect 28077 21295 28135 21301
rect 28629 21335 28687 21341
rect 28629 21301 28641 21335
rect 28675 21332 28687 21335
rect 28902 21332 28908 21344
rect 28675 21304 28908 21332
rect 28675 21301 28687 21304
rect 28629 21295 28687 21301
rect 28902 21292 28908 21304
rect 28960 21292 28966 21344
rect 29012 21332 29040 21372
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 32306 21360 32312 21412
rect 32364 21400 32370 21412
rect 32585 21403 32643 21409
rect 32585 21400 32597 21403
rect 32364 21372 32597 21400
rect 32364 21360 32370 21372
rect 32585 21369 32597 21372
rect 32631 21369 32643 21403
rect 32585 21363 32643 21369
rect 35986 21360 35992 21412
rect 36044 21400 36050 21412
rect 36044 21372 36492 21400
rect 36044 21360 36050 21372
rect 29825 21335 29883 21341
rect 29825 21332 29837 21335
rect 29012 21304 29837 21332
rect 29825 21301 29837 21304
rect 29871 21301 29883 21335
rect 29825 21295 29883 21301
rect 34977 21335 35035 21341
rect 34977 21301 34989 21335
rect 35023 21332 35035 21335
rect 35710 21332 35716 21344
rect 35023 21304 35716 21332
rect 35023 21301 35035 21304
rect 34977 21295 35035 21301
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 35894 21292 35900 21344
rect 35952 21332 35958 21344
rect 36357 21335 36415 21341
rect 36357 21332 36369 21335
rect 35952 21304 36369 21332
rect 35952 21292 35958 21304
rect 36357 21301 36369 21304
rect 36403 21301 36415 21335
rect 36464 21332 36492 21372
rect 37182 21360 37188 21412
rect 37240 21400 37246 21412
rect 38289 21403 38347 21409
rect 38289 21400 38301 21403
rect 37240 21372 38301 21400
rect 37240 21360 37246 21372
rect 38289 21369 38301 21372
rect 38335 21369 38347 21403
rect 38289 21363 38347 21369
rect 39761 21403 39819 21409
rect 39761 21369 39773 21403
rect 39807 21400 39819 21403
rect 39942 21400 39948 21412
rect 39807 21372 39948 21400
rect 39807 21369 39819 21372
rect 39761 21363 39819 21369
rect 39942 21360 39948 21372
rect 40000 21360 40006 21412
rect 40957 21403 41015 21409
rect 40052 21372 40908 21400
rect 37553 21335 37611 21341
rect 37553 21332 37565 21335
rect 36464 21304 37565 21332
rect 36357 21295 36415 21301
rect 37553 21301 37565 21304
rect 37599 21301 37611 21335
rect 39390 21332 39396 21344
rect 39351 21304 39396 21332
rect 37553 21295 37611 21301
rect 39390 21292 39396 21304
rect 39448 21292 39454 21344
rect 39850 21292 39856 21344
rect 39908 21332 39914 21344
rect 40052 21332 40080 21372
rect 39908 21304 40080 21332
rect 39908 21292 39914 21304
rect 40126 21292 40132 21344
rect 40184 21332 40190 21344
rect 40770 21332 40776 21344
rect 40184 21304 40776 21332
rect 40184 21292 40190 21304
rect 40770 21292 40776 21304
rect 40828 21292 40834 21344
rect 40880 21332 40908 21372
rect 40957 21369 40969 21403
rect 41003 21400 41015 21403
rect 41046 21400 41052 21412
rect 41003 21372 41052 21400
rect 41003 21369 41015 21372
rect 40957 21363 41015 21369
rect 41046 21360 41052 21372
rect 41104 21400 41110 21412
rect 41601 21403 41659 21409
rect 41601 21400 41613 21403
rect 41104 21372 41613 21400
rect 41104 21360 41110 21372
rect 41601 21369 41613 21372
rect 41647 21369 41659 21403
rect 41601 21363 41659 21369
rect 41690 21360 41696 21412
rect 41748 21400 41754 21412
rect 43254 21400 43260 21412
rect 41748 21372 43260 21400
rect 41748 21360 41754 21372
rect 43254 21360 43260 21372
rect 43312 21360 43318 21412
rect 43622 21360 43628 21412
rect 43680 21360 43686 21412
rect 42702 21332 42708 21344
rect 40880 21304 42708 21332
rect 42702 21292 42708 21304
rect 42760 21292 42766 21344
rect 42797 21335 42855 21341
rect 42797 21301 42809 21335
rect 42843 21332 42855 21335
rect 42886 21332 42892 21344
rect 42843 21304 42892 21332
rect 42843 21301 42855 21304
rect 42797 21295 42855 21301
rect 42886 21292 42892 21304
rect 42944 21292 42950 21344
rect 44634 21292 44640 21344
rect 44692 21332 44698 21344
rect 45020 21341 45048 21440
rect 45005 21335 45063 21341
rect 45005 21332 45017 21335
rect 44692 21304 45017 21332
rect 44692 21292 44698 21304
rect 45005 21301 45017 21304
rect 45051 21301 45063 21335
rect 46658 21332 46664 21344
rect 46619 21304 46664 21332
rect 45005 21295 45063 21301
rect 46658 21292 46664 21304
rect 46716 21292 46722 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 23477 21131 23535 21137
rect 23477 21128 23489 21131
rect 23440 21100 23489 21128
rect 23440 21088 23446 21100
rect 23477 21097 23489 21100
rect 23523 21097 23535 21131
rect 25774 21128 25780 21140
rect 25735 21100 25780 21128
rect 23477 21091 23535 21097
rect 25774 21088 25780 21100
rect 25832 21088 25838 21140
rect 31202 21128 31208 21140
rect 27632 21100 31208 21128
rect 25682 20952 25688 21004
rect 25740 20992 25746 21004
rect 27632 21001 27660 21100
rect 31202 21088 31208 21100
rect 31260 21088 31266 21140
rect 32398 21128 32404 21140
rect 32359 21100 32404 21128
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 32766 21088 32772 21140
rect 32824 21128 32830 21140
rect 35618 21128 35624 21140
rect 32824 21100 35624 21128
rect 32824 21088 32830 21100
rect 35618 21088 35624 21100
rect 35676 21088 35682 21140
rect 36170 21088 36176 21140
rect 36228 21128 36234 21140
rect 36722 21128 36728 21140
rect 36228 21100 36728 21128
rect 36228 21088 36234 21100
rect 36722 21088 36728 21100
rect 36780 21088 36786 21140
rect 36814 21088 36820 21140
rect 36872 21128 36878 21140
rect 37642 21128 37648 21140
rect 36872 21100 37648 21128
rect 36872 21088 36878 21100
rect 37642 21088 37648 21100
rect 37700 21088 37706 21140
rect 37734 21088 37740 21140
rect 37792 21128 37798 21140
rect 38013 21131 38071 21137
rect 38013 21128 38025 21131
rect 37792 21100 38025 21128
rect 37792 21088 37798 21100
rect 38013 21097 38025 21100
rect 38059 21128 38071 21131
rect 38378 21128 38384 21140
rect 38059 21100 38384 21128
rect 38059 21097 38071 21100
rect 38013 21091 38071 21097
rect 38378 21088 38384 21100
rect 38436 21088 38442 21140
rect 40586 21128 40592 21140
rect 38948 21100 40592 21128
rect 27706 21020 27712 21072
rect 27764 21060 27770 21072
rect 28350 21060 28356 21072
rect 27764 21032 28356 21060
rect 27764 21020 27770 21032
rect 28350 21020 28356 21032
rect 28408 21020 28414 21072
rect 38841 21063 38899 21069
rect 38841 21060 38853 21063
rect 30208 21032 38853 21060
rect 30208 21001 30236 21032
rect 38841 21029 38853 21032
rect 38887 21029 38899 21063
rect 38841 21023 38899 21029
rect 27617 20995 27675 21001
rect 25740 20964 25820 20992
rect 25740 20952 25746 20964
rect 23661 20927 23719 20933
rect 23661 20893 23673 20927
rect 23707 20924 23719 20927
rect 23750 20924 23756 20936
rect 23707 20896 23756 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 23842 20884 23848 20936
rect 23900 20924 23906 20936
rect 25792 20933 25820 20964
rect 27617 20961 27629 20995
rect 27663 20961 27675 20995
rect 27617 20955 27675 20961
rect 30193 20995 30251 21001
rect 30193 20961 30205 20995
rect 30239 20961 30251 20995
rect 30193 20955 30251 20961
rect 32585 20995 32643 21001
rect 32585 20961 32597 20995
rect 32631 20992 32643 20995
rect 33226 20992 33232 21004
rect 32631 20964 33232 20992
rect 32631 20961 32643 20964
rect 32585 20955 32643 20961
rect 33226 20952 33232 20964
rect 33284 20952 33290 21004
rect 33597 20995 33655 21001
rect 33597 20992 33609 20995
rect 33336 20964 33609 20992
rect 25133 20927 25191 20933
rect 23900 20896 23945 20924
rect 23900 20884 23906 20896
rect 25133 20893 25145 20927
rect 25179 20893 25191 20927
rect 25133 20887 25191 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 25777 20927 25835 20933
rect 25363 20896 25728 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 25148 20856 25176 20887
rect 25590 20856 25596 20868
rect 25148 20828 25596 20856
rect 25590 20816 25596 20828
rect 25648 20816 25654 20868
rect 25700 20800 25728 20896
rect 25777 20893 25789 20927
rect 25823 20893 25835 20927
rect 25777 20887 25835 20893
rect 25869 20927 25927 20933
rect 25869 20893 25881 20927
rect 25915 20924 25927 20927
rect 25958 20924 25964 20936
rect 25915 20896 25964 20924
rect 25915 20893 25927 20896
rect 25869 20887 25927 20893
rect 25958 20884 25964 20896
rect 26016 20884 26022 20936
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20924 30159 20927
rect 30147 20896 30236 20924
rect 30147 20893 30159 20896
rect 30101 20887 30159 20893
rect 30208 20868 30236 20896
rect 32214 20884 32220 20936
rect 32272 20924 32278 20936
rect 32309 20927 32367 20933
rect 32309 20924 32321 20927
rect 32272 20896 32321 20924
rect 32272 20884 32278 20896
rect 32309 20893 32321 20896
rect 32355 20893 32367 20927
rect 32309 20887 32367 20893
rect 26050 20856 26056 20868
rect 26011 20828 26056 20856
rect 26050 20816 26056 20828
rect 26108 20816 26114 20868
rect 27341 20859 27399 20865
rect 27341 20825 27353 20859
rect 27387 20856 27399 20859
rect 27890 20856 27896 20868
rect 27387 20828 27896 20856
rect 27387 20825 27399 20828
rect 27341 20819 27399 20825
rect 27890 20816 27896 20828
rect 27948 20816 27954 20868
rect 30190 20816 30196 20868
rect 30248 20816 30254 20868
rect 32324 20856 32352 20887
rect 32950 20856 32956 20868
rect 32324 20828 32956 20856
rect 32950 20816 32956 20828
rect 33008 20856 33014 20868
rect 33336 20856 33364 20964
rect 33597 20961 33609 20964
rect 33643 20961 33655 20995
rect 33597 20955 33655 20961
rect 33980 20964 36308 20992
rect 33980 20936 34008 20964
rect 33781 20927 33839 20933
rect 33781 20893 33793 20927
rect 33827 20893 33839 20927
rect 33781 20887 33839 20893
rect 33873 20927 33931 20933
rect 33873 20893 33885 20927
rect 33919 20924 33931 20927
rect 33962 20924 33968 20936
rect 33919 20896 33968 20924
rect 33919 20893 33931 20896
rect 33873 20887 33931 20893
rect 33796 20856 33824 20887
rect 33962 20884 33968 20896
rect 34020 20884 34026 20936
rect 34882 20884 34888 20936
rect 34940 20924 34946 20936
rect 35526 20924 35532 20936
rect 34940 20896 35532 20924
rect 34940 20884 34946 20896
rect 35526 20884 35532 20896
rect 35584 20884 35590 20936
rect 35713 20927 35771 20933
rect 35713 20893 35725 20927
rect 35759 20924 35771 20927
rect 35986 20924 35992 20936
rect 35759 20896 35992 20924
rect 35759 20893 35771 20896
rect 35713 20887 35771 20893
rect 35986 20884 35992 20896
rect 36044 20884 36050 20936
rect 34054 20856 34060 20868
rect 33008 20828 33364 20856
rect 33428 20828 34060 20856
rect 33008 20816 33014 20828
rect 24946 20788 24952 20800
rect 24907 20760 24952 20788
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 25682 20748 25688 20800
rect 25740 20788 25746 20800
rect 26973 20791 27031 20797
rect 26973 20788 26985 20791
rect 25740 20760 26985 20788
rect 25740 20748 25746 20760
rect 26973 20757 26985 20760
rect 27019 20757 27031 20791
rect 26973 20751 27031 20757
rect 27433 20791 27491 20797
rect 27433 20757 27445 20791
rect 27479 20788 27491 20791
rect 27522 20788 27528 20800
rect 27479 20760 27528 20788
rect 27479 20757 27491 20760
rect 27433 20751 27491 20757
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 29730 20788 29736 20800
rect 29691 20760 29736 20788
rect 29730 20748 29736 20760
rect 29788 20748 29794 20800
rect 31846 20788 31852 20800
rect 31807 20760 31852 20788
rect 31846 20748 31852 20760
rect 31904 20748 31910 20800
rect 32398 20748 32404 20800
rect 32456 20788 32462 20800
rect 32585 20791 32643 20797
rect 32585 20788 32597 20791
rect 32456 20760 32597 20788
rect 32456 20748 32462 20760
rect 32585 20757 32597 20760
rect 32631 20757 32643 20791
rect 32585 20751 32643 20757
rect 33137 20791 33195 20797
rect 33137 20757 33149 20791
rect 33183 20788 33195 20791
rect 33428 20788 33456 20828
rect 34054 20816 34060 20828
rect 34112 20816 34118 20868
rect 35544 20856 35572 20884
rect 35802 20856 35808 20868
rect 35544 20828 35808 20856
rect 35802 20816 35808 20828
rect 35860 20816 35866 20868
rect 35897 20859 35955 20865
rect 35897 20825 35909 20859
rect 35943 20856 35955 20859
rect 36078 20856 36084 20868
rect 35943 20828 36084 20856
rect 35943 20825 35955 20828
rect 35897 20819 35955 20825
rect 36078 20816 36084 20828
rect 36136 20816 36142 20868
rect 36280 20856 36308 20964
rect 36354 20952 36360 21004
rect 36412 20992 36418 21004
rect 36909 20995 36967 21001
rect 36909 20992 36921 20995
rect 36412 20964 36921 20992
rect 36412 20952 36418 20964
rect 36909 20961 36921 20964
rect 36955 20992 36967 20995
rect 37182 20992 37188 21004
rect 36955 20964 37188 20992
rect 36955 20961 36967 20964
rect 36909 20955 36967 20961
rect 37182 20952 37188 20964
rect 37240 20952 37246 21004
rect 37642 20952 37648 21004
rect 37700 20992 37706 21004
rect 38948 20992 38976 21100
rect 40586 21088 40592 21100
rect 40644 21088 40650 21140
rect 41049 21131 41107 21137
rect 41049 21097 41061 21131
rect 41095 21128 41107 21131
rect 41230 21128 41236 21140
rect 41095 21100 41236 21128
rect 41095 21097 41107 21100
rect 41049 21091 41107 21097
rect 41230 21088 41236 21100
rect 41288 21128 41294 21140
rect 41877 21131 41935 21137
rect 41877 21128 41889 21131
rect 41288 21100 41889 21128
rect 41288 21088 41294 21100
rect 41877 21097 41889 21100
rect 41923 21097 41935 21131
rect 41877 21091 41935 21097
rect 42702 21088 42708 21140
rect 42760 21128 42766 21140
rect 42760 21100 43116 21128
rect 42760 21088 42766 21100
rect 39206 21020 39212 21072
rect 39264 21060 39270 21072
rect 39850 21060 39856 21072
rect 39264 21032 39856 21060
rect 39264 21020 39270 21032
rect 39850 21020 39856 21032
rect 39908 21020 39914 21072
rect 40494 21020 40500 21072
rect 40552 21060 40558 21072
rect 43088 21060 43116 21100
rect 45094 21088 45100 21140
rect 45152 21128 45158 21140
rect 46201 21131 46259 21137
rect 46201 21128 46213 21131
rect 45152 21100 46213 21128
rect 45152 21088 45158 21100
rect 46201 21097 46213 21100
rect 46247 21097 46259 21131
rect 46201 21091 46259 21097
rect 45112 21060 45140 21088
rect 40552 21032 42932 21060
rect 40552 21020 40558 21032
rect 37700 20964 38976 20992
rect 39025 20995 39083 21001
rect 37700 20952 37706 20964
rect 39025 20961 39037 20995
rect 39071 20992 39083 20995
rect 39390 20992 39396 21004
rect 39071 20964 39396 20992
rect 39071 20961 39083 20964
rect 39025 20955 39083 20961
rect 39390 20952 39396 20964
rect 39448 20952 39454 21004
rect 40129 20995 40187 21001
rect 40129 20961 40141 20995
rect 40175 20992 40187 20995
rect 40175 20964 41736 20992
rect 40175 20961 40187 20964
rect 40129 20955 40187 20961
rect 36446 20884 36452 20936
rect 36504 20924 36510 20936
rect 36541 20927 36599 20933
rect 36541 20924 36553 20927
rect 36504 20896 36553 20924
rect 36504 20884 36510 20896
rect 36541 20893 36553 20896
rect 36587 20893 36599 20927
rect 36541 20887 36599 20893
rect 36630 20884 36636 20936
rect 36688 20924 36694 20936
rect 37001 20927 37059 20933
rect 36688 20896 36733 20924
rect 36688 20884 36694 20896
rect 37001 20893 37013 20927
rect 37047 20924 37059 20927
rect 37274 20924 37280 20936
rect 37047 20896 37280 20924
rect 37047 20893 37059 20896
rect 37001 20887 37059 20893
rect 37274 20884 37280 20896
rect 37332 20924 37338 20936
rect 37734 20924 37740 20936
rect 37332 20896 37740 20924
rect 37332 20884 37338 20896
rect 37734 20884 37740 20896
rect 37792 20884 37798 20936
rect 38197 20927 38255 20933
rect 38197 20893 38209 20927
rect 38243 20924 38255 20927
rect 38838 20924 38844 20936
rect 38243 20896 38844 20924
rect 38243 20893 38255 20896
rect 38197 20887 38255 20893
rect 38838 20884 38844 20896
rect 38896 20884 38902 20936
rect 39114 20884 39120 20936
rect 39172 20924 39178 20936
rect 40144 20924 40172 20955
rect 41708 20933 41736 20964
rect 41966 20952 41972 21004
rect 42024 20992 42030 21004
rect 42904 21001 42932 21032
rect 43088 21032 45140 21060
rect 42889 20995 42947 21001
rect 42024 20964 42656 20992
rect 42024 20952 42030 20964
rect 39172 20896 39217 20924
rect 39316 20896 40172 20924
rect 40313 20927 40371 20933
rect 39172 20884 39178 20896
rect 37458 20856 37464 20868
rect 36280 20828 37320 20856
rect 37419 20828 37464 20856
rect 37292 20800 37320 20828
rect 37458 20816 37464 20828
rect 37516 20816 37522 20868
rect 38381 20859 38439 20865
rect 38381 20825 38393 20859
rect 38427 20856 38439 20859
rect 38562 20856 38568 20868
rect 38427 20828 38568 20856
rect 38427 20825 38439 20828
rect 38381 20819 38439 20825
rect 38562 20816 38568 20828
rect 38620 20856 38626 20868
rect 39206 20856 39212 20868
rect 38620 20828 39212 20856
rect 38620 20816 38626 20828
rect 39206 20816 39212 20828
rect 39264 20856 39270 20868
rect 39316 20856 39344 20896
rect 40313 20893 40325 20927
rect 40359 20893 40371 20927
rect 40313 20887 40371 20893
rect 41693 20927 41751 20933
rect 41693 20893 41705 20927
rect 41739 20924 41751 20927
rect 42518 20924 42524 20936
rect 41739 20896 42524 20924
rect 41739 20893 41751 20896
rect 41693 20887 41751 20893
rect 39264 20828 39344 20856
rect 39393 20859 39451 20865
rect 39264 20816 39270 20828
rect 39393 20825 39405 20859
rect 39439 20825 39451 20859
rect 39393 20819 39451 20825
rect 39485 20859 39543 20865
rect 39485 20825 39497 20859
rect 39531 20856 39543 20859
rect 40034 20856 40040 20868
rect 39531 20828 40040 20856
rect 39531 20825 39543 20828
rect 39485 20819 39543 20825
rect 33594 20788 33600 20800
rect 33183 20760 33456 20788
rect 33555 20760 33600 20788
rect 33183 20757 33195 20760
rect 33137 20751 33195 20757
rect 33594 20748 33600 20760
rect 33652 20748 33658 20800
rect 35526 20788 35532 20800
rect 35487 20760 35532 20788
rect 35526 20748 35532 20760
rect 35584 20748 35590 20800
rect 35986 20748 35992 20800
rect 36044 20788 36050 20800
rect 36357 20791 36415 20797
rect 36357 20788 36369 20791
rect 36044 20760 36369 20788
rect 36044 20748 36050 20760
rect 36357 20757 36369 20760
rect 36403 20757 36415 20791
rect 36814 20788 36820 20800
rect 36775 20760 36820 20788
rect 36357 20751 36415 20757
rect 36814 20748 36820 20760
rect 36872 20748 36878 20800
rect 37274 20788 37280 20800
rect 37187 20760 37280 20788
rect 37274 20748 37280 20760
rect 37332 20788 37338 20800
rect 37550 20788 37556 20800
rect 37332 20760 37556 20788
rect 37332 20748 37338 20760
rect 37550 20748 37556 20760
rect 37608 20748 37614 20800
rect 39114 20748 39120 20800
rect 39172 20788 39178 20800
rect 39408 20788 39436 20819
rect 40034 20816 40040 20828
rect 40092 20816 40098 20868
rect 39172 20760 39436 20788
rect 39172 20748 39178 20760
rect 39942 20748 39948 20800
rect 40000 20788 40006 20800
rect 40328 20788 40356 20887
rect 42518 20884 42524 20896
rect 42576 20884 42582 20936
rect 42628 20933 42656 20964
rect 42889 20961 42901 20995
rect 42935 20961 42947 20995
rect 42889 20955 42947 20961
rect 43088 20933 43116 21032
rect 43530 20952 43536 21004
rect 43588 20992 43594 21004
rect 43588 20964 45692 20992
rect 43588 20952 43594 20964
rect 45664 20936 45692 20964
rect 42613 20927 42671 20933
rect 42613 20893 42625 20927
rect 42659 20893 42671 20927
rect 42613 20887 42671 20893
rect 42705 20927 42763 20933
rect 42705 20893 42717 20927
rect 42751 20893 42763 20927
rect 42705 20887 42763 20893
rect 42797 20927 42855 20933
rect 42797 20893 42809 20927
rect 42843 20924 42855 20927
rect 43073 20927 43131 20933
rect 42843 20896 43008 20924
rect 42843 20893 42855 20896
rect 42797 20887 42855 20893
rect 42720 20856 42748 20887
rect 42536 20828 42748 20856
rect 42980 20856 43008 20896
rect 43073 20893 43085 20927
rect 43119 20893 43131 20927
rect 43073 20887 43131 20893
rect 43717 20927 43775 20933
rect 43717 20893 43729 20927
rect 43763 20924 43775 20927
rect 43806 20924 43812 20936
rect 43763 20896 43812 20924
rect 43763 20893 43775 20896
rect 43717 20887 43775 20893
rect 43806 20884 43812 20896
rect 43864 20884 43870 20936
rect 43901 20927 43959 20933
rect 43901 20893 43913 20927
rect 43947 20924 43959 20927
rect 44174 20924 44180 20936
rect 43947 20896 44180 20924
rect 43947 20893 43959 20896
rect 43901 20887 43959 20893
rect 44174 20884 44180 20896
rect 44232 20924 44238 20936
rect 45186 20924 45192 20936
rect 44232 20896 45192 20924
rect 44232 20884 44238 20896
rect 45186 20884 45192 20896
rect 45244 20924 45250 20936
rect 45281 20927 45339 20933
rect 45281 20924 45293 20927
rect 45244 20896 45293 20924
rect 45244 20884 45250 20896
rect 45281 20893 45293 20896
rect 45327 20893 45339 20927
rect 45281 20887 45339 20893
rect 45646 20884 45652 20936
rect 45704 20924 45710 20936
rect 45741 20927 45799 20933
rect 45741 20924 45753 20927
rect 45704 20896 45753 20924
rect 45704 20884 45710 20896
rect 45741 20893 45753 20896
rect 45787 20893 45799 20927
rect 45741 20887 45799 20893
rect 44450 20856 44456 20868
rect 42980 20828 44456 20856
rect 42536 20800 42564 20828
rect 40494 20788 40500 20800
rect 40000 20760 40356 20788
rect 40455 20760 40500 20788
rect 40000 20748 40006 20760
rect 40494 20748 40500 20760
rect 40552 20748 40558 20800
rect 42150 20748 42156 20800
rect 42208 20788 42214 20800
rect 42429 20791 42487 20797
rect 42429 20788 42441 20791
rect 42208 20760 42441 20788
rect 42208 20748 42214 20760
rect 42429 20757 42441 20760
rect 42475 20757 42487 20791
rect 42429 20751 42487 20757
rect 42518 20748 42524 20800
rect 42576 20748 42582 20800
rect 42794 20748 42800 20800
rect 42852 20788 42858 20800
rect 42980 20788 43008 20828
rect 44450 20816 44456 20828
rect 44508 20856 44514 20868
rect 45373 20859 45431 20865
rect 45373 20856 45385 20859
rect 44508 20828 45385 20856
rect 44508 20816 44514 20828
rect 45373 20825 45385 20828
rect 45419 20825 45431 20859
rect 45373 20819 45431 20825
rect 42852 20760 43008 20788
rect 43533 20791 43591 20797
rect 42852 20748 42858 20760
rect 43533 20757 43545 20791
rect 43579 20788 43591 20791
rect 43714 20788 43720 20800
rect 43579 20760 43720 20788
rect 43579 20757 43591 20760
rect 43533 20751 43591 20757
rect 43714 20748 43720 20760
rect 43772 20748 43778 20800
rect 43990 20748 43996 20800
rect 44048 20788 44054 20800
rect 44361 20791 44419 20797
rect 44361 20788 44373 20791
rect 44048 20760 44373 20788
rect 44048 20748 44054 20760
rect 44361 20757 44373 20760
rect 44407 20757 44419 20791
rect 44361 20751 44419 20757
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 26970 20544 26976 20596
rect 27028 20584 27034 20596
rect 28721 20587 28779 20593
rect 28721 20584 28733 20587
rect 27028 20556 28733 20584
rect 27028 20544 27034 20556
rect 28721 20553 28733 20556
rect 28767 20553 28779 20587
rect 28721 20547 28779 20553
rect 35526 20544 35532 20596
rect 35584 20584 35590 20596
rect 35805 20587 35863 20593
rect 35805 20584 35817 20587
rect 35584 20556 35817 20584
rect 35584 20544 35590 20556
rect 35805 20553 35817 20556
rect 35851 20553 35863 20587
rect 37550 20584 37556 20596
rect 37511 20556 37556 20584
rect 35805 20547 35863 20553
rect 37550 20544 37556 20556
rect 37608 20584 37614 20596
rect 38470 20584 38476 20596
rect 37608 20556 38476 20584
rect 37608 20544 37614 20556
rect 38470 20544 38476 20556
rect 38528 20584 38534 20596
rect 38565 20587 38623 20593
rect 38565 20584 38577 20587
rect 38528 20556 38577 20584
rect 38528 20544 38534 20556
rect 38565 20553 38577 20556
rect 38611 20553 38623 20587
rect 38565 20547 38623 20553
rect 39022 20544 39028 20596
rect 39080 20584 39086 20596
rect 39298 20584 39304 20596
rect 39080 20556 39304 20584
rect 39080 20544 39086 20556
rect 39298 20544 39304 20556
rect 39356 20584 39362 20596
rect 39393 20587 39451 20593
rect 39393 20584 39405 20587
rect 39356 20556 39405 20584
rect 39356 20544 39362 20556
rect 39393 20553 39405 20556
rect 39439 20553 39451 20587
rect 39393 20547 39451 20553
rect 39482 20544 39488 20596
rect 39540 20584 39546 20596
rect 39540 20556 40172 20584
rect 39540 20544 39546 20556
rect 23566 20476 23572 20528
rect 23624 20516 23630 20528
rect 23661 20519 23719 20525
rect 23661 20516 23673 20519
rect 23624 20488 23673 20516
rect 23624 20476 23630 20488
rect 23661 20485 23673 20488
rect 23707 20485 23719 20519
rect 32309 20519 32367 20525
rect 32309 20516 32321 20519
rect 23661 20479 23719 20485
rect 29932 20488 31524 20516
rect 25596 20460 25648 20466
rect 29932 20460 29960 20488
rect 23014 20408 23020 20460
rect 23072 20408 23078 20460
rect 25682 20408 25688 20460
rect 25740 20448 25746 20460
rect 25740 20420 25785 20448
rect 25740 20408 25746 20420
rect 27246 20408 27252 20460
rect 27304 20448 27310 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27304 20420 27537 20448
rect 27304 20408 27310 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 27709 20451 27767 20457
rect 27709 20417 27721 20451
rect 27755 20448 27767 20451
rect 27890 20448 27896 20460
rect 27755 20420 27896 20448
rect 27755 20417 27767 20420
rect 27709 20411 27767 20417
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28997 20451 29055 20457
rect 28997 20417 29009 20451
rect 29043 20448 29055 20451
rect 29914 20448 29920 20460
rect 29043 20420 29920 20448
rect 29043 20417 29055 20420
rect 28997 20411 29055 20417
rect 29914 20408 29920 20420
rect 29972 20408 29978 20460
rect 30190 20448 30196 20460
rect 30151 20420 30196 20448
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 30374 20408 30380 20460
rect 30432 20448 30438 20460
rect 31113 20451 31171 20457
rect 31113 20448 31125 20451
rect 30432 20420 31125 20448
rect 30432 20408 30438 20420
rect 31113 20417 31125 20420
rect 31159 20417 31171 20451
rect 31113 20411 31171 20417
rect 31297 20451 31355 20457
rect 31297 20417 31309 20451
rect 31343 20417 31355 20451
rect 31297 20411 31355 20417
rect 31389 20451 31447 20457
rect 31389 20417 31401 20451
rect 31435 20417 31447 20451
rect 31389 20411 31447 20417
rect 25596 20402 25648 20408
rect 22830 20340 22836 20392
rect 22888 20380 22894 20392
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 22888 20352 24685 20380
rect 22888 20340 22894 20352
rect 24673 20349 24685 20352
rect 24719 20349 24731 20383
rect 28718 20380 28724 20392
rect 28679 20352 28724 20380
rect 24673 20343 24731 20349
rect 28718 20340 28724 20352
rect 28776 20340 28782 20392
rect 28905 20383 28963 20389
rect 28905 20349 28917 20383
rect 28951 20380 28963 20383
rect 29730 20380 29736 20392
rect 28951 20352 29736 20380
rect 28951 20349 28963 20352
rect 28905 20343 28963 20349
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 27522 20312 27528 20324
rect 27483 20284 27528 20312
rect 27522 20272 27528 20284
rect 27580 20272 27586 20324
rect 29730 20244 29736 20256
rect 29691 20216 29736 20244
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 30282 20244 30288 20256
rect 30243 20216 30288 20244
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 31312 20244 31340 20411
rect 31404 20312 31432 20411
rect 31496 20380 31524 20488
rect 31588 20488 32321 20516
rect 31588 20457 31616 20488
rect 32309 20485 32321 20488
rect 32355 20485 32367 20519
rect 32309 20479 32367 20485
rect 32490 20476 32496 20528
rect 32548 20516 32554 20528
rect 35621 20519 35679 20525
rect 32548 20488 32720 20516
rect 32548 20476 32554 20488
rect 32692 20457 32720 20488
rect 35621 20485 35633 20519
rect 35667 20516 35679 20519
rect 35986 20516 35992 20528
rect 35667 20488 35992 20516
rect 35667 20485 35679 20488
rect 35621 20479 35679 20485
rect 35986 20476 35992 20488
rect 36044 20476 36050 20528
rect 36078 20476 36084 20528
rect 36136 20516 36142 20528
rect 40144 20525 40172 20556
rect 40678 20544 40684 20596
rect 40736 20584 40742 20596
rect 41138 20584 41144 20596
rect 40736 20556 41144 20584
rect 40736 20544 40742 20556
rect 41138 20544 41144 20556
rect 41196 20584 41202 20596
rect 41782 20584 41788 20596
rect 41196 20556 41788 20584
rect 41196 20544 41202 20556
rect 41782 20544 41788 20556
rect 41840 20544 41846 20596
rect 41966 20544 41972 20596
rect 42024 20584 42030 20596
rect 42024 20556 42748 20584
rect 42024 20544 42030 20556
rect 38841 20519 38899 20525
rect 36136 20488 36492 20516
rect 36136 20476 36142 20488
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31665 20451 31723 20457
rect 31665 20417 31677 20451
rect 31711 20417 31723 20451
rect 31665 20411 31723 20417
rect 32585 20451 32643 20457
rect 32585 20417 32597 20451
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 32677 20451 32735 20457
rect 32677 20417 32689 20451
rect 32723 20417 32735 20451
rect 32677 20411 32735 20417
rect 31680 20380 31708 20411
rect 31496 20352 31708 20380
rect 31846 20312 31852 20324
rect 31404 20284 31852 20312
rect 31846 20272 31852 20284
rect 31904 20272 31910 20324
rect 32600 20312 32628 20411
rect 32766 20408 32772 20460
rect 32824 20448 32830 20460
rect 32953 20451 33011 20457
rect 32824 20420 32869 20448
rect 32824 20408 32830 20420
rect 32953 20417 32965 20451
rect 32999 20448 33011 20451
rect 33042 20448 33048 20460
rect 32999 20420 33048 20448
rect 32999 20417 33011 20420
rect 32953 20411 33011 20417
rect 33042 20408 33048 20420
rect 33100 20408 33106 20460
rect 33870 20448 33876 20460
rect 33831 20420 33876 20448
rect 33870 20408 33876 20420
rect 33928 20408 33934 20460
rect 34701 20451 34759 20457
rect 34701 20417 34713 20451
rect 34747 20448 34759 20451
rect 34882 20448 34888 20460
rect 34747 20420 34888 20448
rect 34747 20417 34759 20420
rect 34701 20411 34759 20417
rect 34882 20408 34888 20420
rect 34940 20408 34946 20460
rect 35894 20448 35900 20460
rect 35855 20420 35900 20448
rect 35894 20408 35900 20420
rect 35952 20408 35958 20460
rect 36354 20448 36360 20460
rect 36267 20420 36360 20448
rect 36354 20408 36360 20420
rect 36412 20408 36418 20460
rect 34149 20383 34207 20389
rect 34149 20349 34161 20383
rect 34195 20380 34207 20383
rect 34790 20380 34796 20392
rect 34195 20352 34796 20380
rect 34195 20349 34207 20352
rect 34149 20343 34207 20349
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 35710 20340 35716 20392
rect 35768 20380 35774 20392
rect 36372 20380 36400 20408
rect 36464 20389 36492 20488
rect 38841 20485 38853 20519
rect 38887 20516 38899 20519
rect 40129 20519 40187 20525
rect 38887 20488 40080 20516
rect 38887 20485 38899 20488
rect 38841 20479 38899 20485
rect 36541 20451 36599 20457
rect 36541 20417 36553 20451
rect 36587 20448 36599 20451
rect 36630 20448 36636 20460
rect 36587 20420 36636 20448
rect 36587 20417 36599 20420
rect 36541 20411 36599 20417
rect 36630 20408 36636 20420
rect 36688 20408 36694 20460
rect 37458 20448 37464 20460
rect 37419 20420 37464 20448
rect 37458 20408 37464 20420
rect 37516 20408 37522 20460
rect 37737 20451 37795 20457
rect 37737 20417 37749 20451
rect 37783 20448 37795 20451
rect 39298 20448 39304 20460
rect 37783 20420 39304 20448
rect 37783 20417 37795 20420
rect 37737 20411 37795 20417
rect 39298 20408 39304 20420
rect 39356 20408 39362 20460
rect 39393 20451 39451 20457
rect 39393 20417 39405 20451
rect 39439 20417 39451 20451
rect 39393 20411 39451 20417
rect 39577 20451 39635 20457
rect 39577 20417 39589 20451
rect 39623 20448 39635 20451
rect 39942 20448 39948 20460
rect 39623 20420 39948 20448
rect 39623 20417 39635 20420
rect 39577 20411 39635 20417
rect 35768 20352 36400 20380
rect 36449 20383 36507 20389
rect 35768 20340 35774 20352
rect 36449 20349 36461 20383
rect 36495 20380 36507 20383
rect 39408 20380 39436 20411
rect 39942 20408 39948 20420
rect 40000 20408 40006 20460
rect 40052 20448 40080 20488
rect 40129 20485 40141 20519
rect 40175 20485 40187 20519
rect 40129 20479 40187 20485
rect 40218 20476 40224 20528
rect 40276 20516 40282 20528
rect 40329 20519 40387 20525
rect 40329 20516 40341 20519
rect 40276 20488 40341 20516
rect 40276 20476 40282 20488
rect 40329 20485 40341 20488
rect 40375 20485 40387 20519
rect 40329 20479 40387 20485
rect 40494 20476 40500 20528
rect 40552 20516 40558 20528
rect 42613 20519 42671 20525
rect 42613 20516 42625 20519
rect 40552 20488 42625 20516
rect 40552 20476 40558 20488
rect 42613 20485 42625 20488
rect 42659 20485 42671 20519
rect 42613 20479 42671 20485
rect 40862 20448 40868 20460
rect 40052 20420 40868 20448
rect 40862 20408 40868 20420
rect 40920 20448 40926 20460
rect 40957 20451 41015 20457
rect 40957 20448 40969 20451
rect 40920 20420 40969 20448
rect 40920 20408 40926 20420
rect 40957 20417 40969 20420
rect 41003 20417 41015 20451
rect 40957 20411 41015 20417
rect 41046 20408 41052 20460
rect 41104 20448 41110 20460
rect 41141 20451 41199 20457
rect 41141 20448 41153 20451
rect 41104 20420 41153 20448
rect 41104 20408 41110 20420
rect 41141 20417 41153 20420
rect 41187 20417 41199 20451
rect 41141 20411 41199 20417
rect 41785 20451 41843 20457
rect 41785 20417 41797 20451
rect 41831 20448 41843 20451
rect 41874 20448 41880 20460
rect 41831 20420 41880 20448
rect 41831 20417 41843 20420
rect 41785 20411 41843 20417
rect 41874 20408 41880 20420
rect 41932 20408 41938 20460
rect 41969 20451 42027 20457
rect 41969 20417 41981 20451
rect 42015 20448 42027 20451
rect 42242 20448 42248 20460
rect 42015 20420 42248 20448
rect 42015 20417 42027 20420
rect 41969 20411 42027 20417
rect 42242 20408 42248 20420
rect 42300 20448 42306 20460
rect 42426 20448 42432 20460
rect 42300 20420 42432 20448
rect 42300 20408 42306 20420
rect 42426 20408 42432 20420
rect 42484 20408 42490 20460
rect 42720 20457 42748 20556
rect 43438 20544 43444 20596
rect 43496 20584 43502 20596
rect 43806 20584 43812 20596
rect 43496 20556 43812 20584
rect 43496 20544 43502 20556
rect 43806 20544 43812 20556
rect 43864 20584 43870 20596
rect 44519 20587 44577 20593
rect 44519 20584 44531 20587
rect 43864 20556 44531 20584
rect 43864 20544 43870 20556
rect 44519 20553 44531 20556
rect 44565 20553 44577 20587
rect 44519 20547 44577 20553
rect 44729 20519 44787 20525
rect 44729 20485 44741 20519
rect 44775 20485 44787 20519
rect 44729 20479 44787 20485
rect 42705 20451 42763 20457
rect 42705 20417 42717 20451
rect 42751 20417 42763 20451
rect 42886 20448 42892 20460
rect 42847 20420 42892 20448
rect 42705 20411 42763 20417
rect 42886 20408 42892 20420
rect 42944 20408 42950 20460
rect 43346 20408 43352 20460
rect 43404 20448 43410 20460
rect 43625 20451 43683 20457
rect 43625 20448 43637 20451
rect 43404 20420 43637 20448
rect 43404 20408 43410 20420
rect 43625 20417 43637 20420
rect 43671 20417 43683 20451
rect 43625 20411 43683 20417
rect 43714 20408 43720 20460
rect 43772 20448 43778 20460
rect 43809 20451 43867 20457
rect 43809 20448 43821 20451
rect 43772 20420 43821 20448
rect 43772 20408 43778 20420
rect 43809 20417 43821 20420
rect 43855 20417 43867 20451
rect 43809 20411 43867 20417
rect 44174 20408 44180 20460
rect 44232 20448 44238 20460
rect 44744 20448 44772 20479
rect 45094 20476 45100 20528
rect 45152 20516 45158 20528
rect 45465 20519 45523 20525
rect 45465 20516 45477 20519
rect 45152 20488 45477 20516
rect 45152 20476 45158 20488
rect 45465 20485 45477 20488
rect 45511 20485 45523 20519
rect 45465 20479 45523 20485
rect 45186 20448 45192 20460
rect 44232 20420 44772 20448
rect 45147 20420 45192 20448
rect 44232 20408 44238 20420
rect 45186 20408 45192 20420
rect 45244 20408 45250 20460
rect 45646 20448 45652 20460
rect 45607 20420 45652 20448
rect 45646 20408 45652 20420
rect 45704 20408 45710 20460
rect 41230 20380 41236 20392
rect 36495 20352 38654 20380
rect 39408 20352 41236 20380
rect 36495 20349 36507 20352
rect 36449 20343 36507 20349
rect 32600 20284 34284 20312
rect 33410 20244 33416 20256
rect 31312 20216 33416 20244
rect 33410 20204 33416 20216
rect 33468 20204 33474 20256
rect 33686 20244 33692 20256
rect 33647 20216 33692 20244
rect 33686 20204 33692 20216
rect 33744 20204 33750 20256
rect 34054 20244 34060 20256
rect 34015 20216 34060 20244
rect 34054 20204 34060 20216
rect 34112 20204 34118 20256
rect 34256 20244 34284 20284
rect 34330 20272 34336 20324
rect 34388 20312 34394 20324
rect 35621 20315 35679 20321
rect 35621 20312 35633 20315
rect 34388 20284 35633 20312
rect 34388 20272 34394 20284
rect 35621 20281 35633 20284
rect 35667 20281 35679 20315
rect 37734 20312 37740 20324
rect 37695 20284 37740 20312
rect 35621 20275 35679 20281
rect 37734 20272 37740 20284
rect 37792 20272 37798 20324
rect 38626 20312 38654 20352
rect 41230 20340 41236 20352
rect 41288 20380 41294 20392
rect 42058 20380 42064 20392
rect 41288 20352 42064 20380
rect 41288 20340 41294 20352
rect 42058 20340 42064 20352
rect 42116 20340 42122 20392
rect 40218 20312 40224 20324
rect 38626 20284 40224 20312
rect 40218 20272 40224 20284
rect 40276 20272 40282 20324
rect 41046 20312 41052 20324
rect 40328 20284 41052 20312
rect 34885 20247 34943 20253
rect 34885 20244 34897 20247
rect 34256 20216 34897 20244
rect 34885 20213 34897 20216
rect 34931 20244 34943 20247
rect 35434 20244 35440 20256
rect 34931 20216 35440 20244
rect 34931 20213 34943 20216
rect 34885 20207 34943 20213
rect 35434 20204 35440 20216
rect 35492 20244 35498 20256
rect 36354 20244 36360 20256
rect 35492 20216 36360 20244
rect 35492 20204 35498 20216
rect 36354 20204 36360 20216
rect 36412 20244 36418 20256
rect 36630 20244 36636 20256
rect 36412 20216 36636 20244
rect 36412 20204 36418 20216
rect 36630 20204 36636 20216
rect 36688 20204 36694 20256
rect 39298 20204 39304 20256
rect 39356 20244 39362 20256
rect 40126 20244 40132 20256
rect 39356 20216 40132 20244
rect 39356 20204 39362 20216
rect 40126 20204 40132 20216
rect 40184 20204 40190 20256
rect 40328 20253 40356 20284
rect 41046 20272 41052 20284
rect 41104 20272 41110 20324
rect 43622 20312 43628 20324
rect 43583 20284 43628 20312
rect 43622 20272 43628 20284
rect 43680 20272 43686 20324
rect 44266 20272 44272 20324
rect 44324 20312 44330 20324
rect 45922 20312 45928 20324
rect 44324 20284 45928 20312
rect 44324 20272 44330 20284
rect 45922 20272 45928 20284
rect 45980 20272 45986 20324
rect 40313 20247 40371 20253
rect 40313 20213 40325 20247
rect 40359 20213 40371 20247
rect 40313 20207 40371 20213
rect 40497 20247 40555 20253
rect 40497 20213 40509 20247
rect 40543 20244 40555 20247
rect 40586 20244 40592 20256
rect 40543 20216 40592 20244
rect 40543 20213 40555 20216
rect 40497 20207 40555 20213
rect 40586 20204 40592 20216
rect 40644 20204 40650 20256
rect 41138 20244 41144 20256
rect 41099 20216 41144 20244
rect 41138 20204 41144 20216
rect 41196 20204 41202 20256
rect 41690 20204 41696 20256
rect 41748 20244 41754 20256
rect 41785 20247 41843 20253
rect 41785 20244 41797 20247
rect 41748 20216 41797 20244
rect 41748 20204 41754 20216
rect 41785 20213 41797 20216
rect 41831 20213 41843 20247
rect 44358 20244 44364 20256
rect 44319 20216 44364 20244
rect 41785 20207 41843 20213
rect 44358 20204 44364 20216
rect 44416 20204 44422 20256
rect 44542 20244 44548 20256
rect 44503 20216 44548 20244
rect 44542 20204 44548 20216
rect 44600 20204 44606 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 23201 20043 23259 20049
rect 23201 20009 23213 20043
rect 23247 20040 23259 20043
rect 23658 20040 23664 20052
rect 23247 20012 23664 20040
rect 23247 20009 23259 20012
rect 23201 20003 23259 20009
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 23750 20000 23756 20052
rect 23808 20040 23814 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23808 20012 24041 20040
rect 23808 20000 23814 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24029 20003 24087 20009
rect 25777 20043 25835 20049
rect 25777 20009 25789 20043
rect 25823 20040 25835 20043
rect 26050 20040 26056 20052
rect 25823 20012 26056 20040
rect 25823 20009 25835 20012
rect 25777 20003 25835 20009
rect 26050 20000 26056 20012
rect 26108 20000 26114 20052
rect 27246 20040 27252 20052
rect 27207 20012 27252 20040
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 27433 20043 27491 20049
rect 27433 20009 27445 20043
rect 27479 20040 27491 20043
rect 28258 20040 28264 20052
rect 27479 20012 28264 20040
rect 27479 20009 27491 20012
rect 27433 20003 27491 20009
rect 25406 19932 25412 19984
rect 25464 19972 25470 19984
rect 25685 19975 25743 19981
rect 25685 19972 25697 19975
rect 25464 19944 25697 19972
rect 25464 19932 25470 19944
rect 25685 19941 25697 19944
rect 25731 19972 25743 19975
rect 26237 19975 26295 19981
rect 26237 19972 26249 19975
rect 25731 19944 26249 19972
rect 25731 19941 25743 19944
rect 25685 19935 25743 19941
rect 26237 19941 26249 19944
rect 26283 19941 26295 19975
rect 26237 19935 26295 19941
rect 22830 19904 22836 19916
rect 22791 19876 22836 19904
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 26697 19907 26755 19913
rect 26697 19873 26709 19907
rect 26743 19904 26755 19907
rect 27448 19904 27476 20003
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 30742 20040 30748 20052
rect 30703 20012 30748 20040
rect 30742 20000 30748 20012
rect 30800 20000 30806 20052
rect 32033 20043 32091 20049
rect 32033 20009 32045 20043
rect 32079 20040 32091 20043
rect 32490 20040 32496 20052
rect 32079 20012 32496 20040
rect 32079 20009 32091 20012
rect 32033 20003 32091 20009
rect 32490 20000 32496 20012
rect 32548 20000 32554 20052
rect 33134 20000 33140 20052
rect 33192 20040 33198 20052
rect 33321 20043 33379 20049
rect 33321 20040 33333 20043
rect 33192 20012 33333 20040
rect 33192 20000 33198 20012
rect 33321 20009 33333 20012
rect 33367 20009 33379 20043
rect 33321 20003 33379 20009
rect 34054 20000 34060 20052
rect 34112 20040 34118 20052
rect 34333 20043 34391 20049
rect 34333 20040 34345 20043
rect 34112 20012 34345 20040
rect 34112 20000 34118 20012
rect 34333 20009 34345 20012
rect 34379 20040 34391 20043
rect 35618 20040 35624 20052
rect 34379 20012 35624 20040
rect 34379 20009 34391 20012
rect 34333 20003 34391 20009
rect 35618 20000 35624 20012
rect 35676 20000 35682 20052
rect 35802 20000 35808 20052
rect 35860 20040 35866 20052
rect 40770 20040 40776 20052
rect 35860 20012 40776 20040
rect 35860 20000 35866 20012
rect 40770 20000 40776 20012
rect 40828 20040 40834 20052
rect 40828 20012 41276 20040
rect 40828 20000 40834 20012
rect 27801 19975 27859 19981
rect 27801 19941 27813 19975
rect 27847 19972 27859 19975
rect 32858 19972 32864 19984
rect 27847 19944 32864 19972
rect 27847 19941 27859 19944
rect 27801 19935 27859 19941
rect 32858 19932 32864 19944
rect 32916 19932 32922 19984
rect 35894 19972 35900 19984
rect 35855 19944 35900 19972
rect 35894 19932 35900 19944
rect 35952 19932 35958 19984
rect 35986 19932 35992 19984
rect 36044 19972 36050 19984
rect 36446 19972 36452 19984
rect 36044 19944 36452 19972
rect 36044 19932 36050 19944
rect 36446 19932 36452 19944
rect 36504 19972 36510 19984
rect 36998 19972 37004 19984
rect 36504 19944 37004 19972
rect 36504 19932 36510 19944
rect 36998 19932 37004 19944
rect 37056 19972 37062 19984
rect 40678 19972 40684 19984
rect 37056 19944 40684 19972
rect 37056 19932 37062 19944
rect 40678 19932 40684 19944
rect 40736 19932 40742 19984
rect 26743 19876 27476 19904
rect 26743 19873 26755 19876
rect 26697 19867 26755 19873
rect 27890 19864 27896 19916
rect 27948 19904 27954 19916
rect 28721 19907 28779 19913
rect 27948 19876 28580 19904
rect 27948 19864 27954 19876
rect 23014 19836 23020 19848
rect 22927 19808 23020 19836
rect 23014 19796 23020 19808
rect 23072 19796 23078 19848
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23532 19808 23673 19836
rect 23532 19796 23538 19808
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23661 19799 23719 19805
rect 23750 19796 23756 19848
rect 23808 19836 23814 19848
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 23808 19808 23857 19836
rect 23808 19796 23814 19808
rect 23845 19805 23857 19808
rect 23891 19836 23903 19839
rect 24946 19836 24952 19848
rect 23891 19808 24952 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 26602 19836 26608 19848
rect 26563 19808 26608 19836
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 28258 19836 28264 19848
rect 28219 19808 28264 19836
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19805 28503 19839
rect 28552 19836 28580 19876
rect 28721 19873 28733 19907
rect 28767 19904 28779 19907
rect 29086 19904 29092 19916
rect 28767 19876 29092 19904
rect 28767 19873 28779 19876
rect 28721 19867 28779 19873
rect 29086 19864 29092 19876
rect 29144 19864 29150 19916
rect 31757 19907 31815 19913
rect 31757 19873 31769 19907
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 32677 19907 32735 19913
rect 32677 19873 32689 19907
rect 32723 19904 32735 19907
rect 35526 19904 35532 19916
rect 32723 19876 35532 19904
rect 32723 19873 32735 19876
rect 32677 19867 32735 19873
rect 28813 19839 28871 19845
rect 28813 19836 28825 19839
rect 28552 19808 28825 19836
rect 28445 19799 28503 19805
rect 28813 19805 28825 19808
rect 28859 19805 28871 19839
rect 28813 19799 28871 19805
rect 23032 19700 23060 19796
rect 25314 19768 25320 19780
rect 25275 19740 25320 19768
rect 25314 19728 25320 19740
rect 25372 19728 25378 19780
rect 27433 19771 27491 19777
rect 27433 19737 27445 19771
rect 27479 19768 27491 19771
rect 27614 19768 27620 19780
rect 27479 19740 27620 19768
rect 27479 19737 27491 19740
rect 27433 19731 27491 19737
rect 27614 19728 27620 19740
rect 27672 19768 27678 19780
rect 28460 19768 28488 19799
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30282 19845 30288 19848
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 29788 19808 30113 19836
rect 29788 19796 29794 19808
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30280 19836 30288 19845
rect 30243 19808 30288 19836
rect 30101 19799 30159 19805
rect 30280 19799 30288 19808
rect 30282 19796 30288 19799
rect 30340 19796 30346 19848
rect 30558 19845 30564 19848
rect 30515 19839 30564 19845
rect 30396 19833 30454 19839
rect 30396 19830 30408 19833
rect 30392 19814 30408 19830
rect 30379 19799 30408 19814
rect 30442 19799 30454 19833
rect 30515 19805 30527 19839
rect 30561 19805 30564 19839
rect 30515 19799 30564 19805
rect 27672 19740 28488 19768
rect 30379 19793 30454 19799
rect 30558 19796 30564 19799
rect 30616 19796 30622 19848
rect 30379 19786 30420 19793
rect 27672 19728 27678 19740
rect 30379 19712 30407 19786
rect 31772 19768 31800 19867
rect 31835 19839 31893 19845
rect 31835 19805 31847 19839
rect 31881 19836 31893 19839
rect 32692 19836 32720 19867
rect 35526 19864 35532 19876
rect 35584 19864 35590 19916
rect 41138 19904 41144 19916
rect 38856 19876 41144 19904
rect 31881 19808 32720 19836
rect 31881 19805 31893 19808
rect 31835 19799 31893 19805
rect 33042 19796 33048 19848
rect 33100 19836 33106 19848
rect 33502 19836 33508 19848
rect 33100 19808 33508 19836
rect 33100 19796 33106 19808
rect 33502 19796 33508 19808
rect 33560 19796 33566 19848
rect 33778 19836 33784 19848
rect 33739 19808 33784 19836
rect 33778 19796 33784 19808
rect 33836 19796 33842 19848
rect 34238 19796 34244 19848
rect 34296 19836 34302 19848
rect 35342 19836 35348 19848
rect 34296 19808 35348 19836
rect 34296 19796 34302 19808
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 35434 19796 35440 19848
rect 35492 19836 35498 19848
rect 35897 19839 35955 19845
rect 35897 19836 35909 19839
rect 35492 19808 35909 19836
rect 35492 19796 35498 19808
rect 35897 19805 35909 19808
rect 35943 19805 35955 19839
rect 36078 19836 36084 19848
rect 36039 19808 36084 19836
rect 35897 19799 35955 19805
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 36173 19839 36231 19845
rect 36173 19805 36185 19839
rect 36219 19805 36231 19839
rect 36173 19799 36231 19805
rect 33689 19771 33747 19777
rect 33689 19768 33701 19771
rect 31772 19740 33701 19768
rect 33689 19737 33701 19740
rect 33735 19768 33747 19771
rect 33962 19768 33968 19780
rect 33735 19740 33968 19768
rect 33735 19737 33747 19740
rect 33689 19731 33747 19737
rect 33962 19728 33968 19740
rect 34020 19728 34026 19780
rect 34054 19728 34060 19780
rect 34112 19768 34118 19780
rect 35802 19768 35808 19780
rect 34112 19740 35808 19768
rect 34112 19728 34118 19740
rect 35802 19728 35808 19740
rect 35860 19728 35866 19780
rect 36188 19768 36216 19799
rect 36354 19796 36360 19848
rect 36412 19836 36418 19848
rect 37277 19839 37335 19845
rect 37277 19836 37289 19839
rect 36412 19808 37289 19836
rect 36412 19796 36418 19808
rect 37277 19805 37289 19808
rect 37323 19805 37335 19839
rect 37458 19836 37464 19848
rect 37419 19808 37464 19836
rect 37277 19799 37335 19805
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 37826 19796 37832 19848
rect 37884 19836 37890 19848
rect 37921 19839 37979 19845
rect 37921 19836 37933 19839
rect 37884 19808 37933 19836
rect 37884 19796 37890 19808
rect 37921 19805 37933 19808
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 38105 19839 38163 19845
rect 38105 19805 38117 19839
rect 38151 19836 38163 19839
rect 38194 19836 38200 19848
rect 38151 19808 38200 19836
rect 38151 19805 38163 19808
rect 38105 19799 38163 19805
rect 38194 19796 38200 19808
rect 38252 19836 38258 19848
rect 38470 19836 38476 19848
rect 38252 19808 38476 19836
rect 38252 19796 38258 19808
rect 38470 19796 38476 19808
rect 38528 19796 38534 19848
rect 38856 19845 38884 19876
rect 38841 19839 38899 19845
rect 38841 19805 38853 19839
rect 38887 19805 38899 19839
rect 38841 19799 38899 19805
rect 38933 19839 38991 19845
rect 38933 19805 38945 19839
rect 38979 19836 38991 19839
rect 39209 19839 39267 19845
rect 38979 19808 39160 19836
rect 38979 19805 38991 19808
rect 38933 19799 38991 19805
rect 39022 19768 39028 19780
rect 36188 19740 38700 19768
rect 38983 19740 39028 19768
rect 29730 19700 29736 19712
rect 23032 19672 29736 19700
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30374 19660 30380 19712
rect 30432 19660 30438 19712
rect 31846 19660 31852 19712
rect 31904 19700 31910 19712
rect 33318 19700 33324 19712
rect 31904 19672 33324 19700
rect 31904 19660 31910 19672
rect 33318 19660 33324 19672
rect 33376 19700 33382 19712
rect 35434 19700 35440 19712
rect 33376 19672 35440 19700
rect 33376 19660 33382 19672
rect 35434 19660 35440 19672
rect 35492 19660 35498 19712
rect 35526 19660 35532 19712
rect 35584 19700 35590 19712
rect 36446 19700 36452 19712
rect 35584 19672 36452 19700
rect 35584 19660 35590 19672
rect 36446 19660 36452 19672
rect 36504 19700 36510 19712
rect 36633 19703 36691 19709
rect 36633 19700 36645 19703
rect 36504 19672 36645 19700
rect 36504 19660 36510 19672
rect 36633 19669 36645 19672
rect 36679 19669 36691 19703
rect 37366 19700 37372 19712
rect 37327 19672 37372 19700
rect 36633 19663 36691 19669
rect 37366 19660 37372 19672
rect 37424 19660 37430 19712
rect 37458 19660 37464 19712
rect 37516 19700 37522 19712
rect 38672 19709 38700 19740
rect 39022 19728 39028 19740
rect 39080 19728 39086 19780
rect 39132 19768 39160 19808
rect 39209 19805 39221 19839
rect 39255 19836 39267 19839
rect 39482 19836 39488 19848
rect 39255 19808 39488 19836
rect 39255 19805 39267 19808
rect 39209 19799 39267 19805
rect 39482 19796 39488 19808
rect 39540 19796 39546 19848
rect 40034 19836 40040 19848
rect 39995 19808 40040 19836
rect 40034 19796 40040 19808
rect 40092 19796 40098 19848
rect 40218 19836 40224 19848
rect 40179 19808 40224 19836
rect 40218 19796 40224 19808
rect 40276 19796 40282 19848
rect 40328 19845 40356 19876
rect 41138 19864 41144 19876
rect 41196 19864 41202 19916
rect 40313 19839 40371 19845
rect 40313 19805 40325 19839
rect 40359 19805 40371 19839
rect 40494 19836 40500 19848
rect 40455 19808 40500 19836
rect 40313 19799 40371 19805
rect 40494 19796 40500 19808
rect 40552 19796 40558 19848
rect 40586 19796 40592 19848
rect 40644 19836 40650 19848
rect 41248 19836 41276 20012
rect 41966 20000 41972 20052
rect 42024 20040 42030 20052
rect 44818 20040 44824 20052
rect 42024 20012 44824 20040
rect 42024 20000 42030 20012
rect 44818 20000 44824 20012
rect 44876 20000 44882 20052
rect 46014 20000 46020 20052
rect 46072 20040 46078 20052
rect 46201 20043 46259 20049
rect 46201 20040 46213 20043
rect 46072 20012 46213 20040
rect 46072 20000 46078 20012
rect 46201 20009 46213 20012
rect 46247 20009 46259 20043
rect 46201 20003 46259 20009
rect 41690 19972 41696 19984
rect 41651 19944 41696 19972
rect 41690 19932 41696 19944
rect 41748 19932 41754 19984
rect 41874 19932 41880 19984
rect 41932 19972 41938 19984
rect 42334 19972 42340 19984
rect 41932 19944 42340 19972
rect 41932 19932 41938 19944
rect 42334 19932 42340 19944
rect 42392 19972 42398 19984
rect 42429 19975 42487 19981
rect 42429 19972 42441 19975
rect 42392 19944 42441 19972
rect 42392 19932 42398 19944
rect 42429 19941 42441 19944
rect 42475 19941 42487 19975
rect 44637 19975 44695 19981
rect 44637 19972 44649 19975
rect 42429 19935 42487 19941
rect 42996 19944 44649 19972
rect 41601 19907 41659 19913
rect 41601 19873 41613 19907
rect 41647 19904 41659 19907
rect 42996 19904 43024 19944
rect 44637 19941 44649 19944
rect 44683 19941 44695 19975
rect 44637 19935 44695 19941
rect 44082 19904 44088 19916
rect 41647 19876 43024 19904
rect 43088 19876 44088 19904
rect 41647 19873 41659 19876
rect 41601 19867 41659 19873
rect 41506 19836 41512 19848
rect 40644 19808 40689 19836
rect 41248 19808 41512 19836
rect 40644 19796 40650 19808
rect 41506 19796 41512 19808
rect 41564 19796 41570 19848
rect 41782 19836 41788 19848
rect 41743 19808 41788 19836
rect 41782 19796 41788 19808
rect 41840 19796 41846 19848
rect 41966 19836 41972 19848
rect 41927 19808 41972 19836
rect 41966 19796 41972 19808
rect 42024 19796 42030 19848
rect 42610 19796 42616 19848
rect 42668 19836 42674 19848
rect 42705 19839 42763 19845
rect 42705 19836 42717 19839
rect 42668 19808 42717 19836
rect 42668 19796 42674 19808
rect 42705 19805 42717 19808
rect 42751 19836 42763 19839
rect 43088 19836 43116 19876
rect 44082 19864 44088 19876
rect 44140 19864 44146 19916
rect 44266 19904 44272 19916
rect 44227 19876 44272 19904
rect 44266 19864 44272 19876
rect 44324 19864 44330 19916
rect 44450 19904 44456 19916
rect 44411 19876 44456 19904
rect 44450 19864 44456 19876
rect 44508 19864 44514 19916
rect 45186 19904 45192 19916
rect 45147 19876 45192 19904
rect 45186 19864 45192 19876
rect 45244 19864 45250 19916
rect 46658 19904 46664 19916
rect 45480 19876 46664 19904
rect 43438 19836 43444 19848
rect 42751 19808 43116 19836
rect 43180 19808 43444 19836
rect 42751 19805 42763 19808
rect 42705 19799 42763 19805
rect 42429 19771 42487 19777
rect 39132 19740 41736 19768
rect 38013 19703 38071 19709
rect 38013 19700 38025 19703
rect 37516 19672 38025 19700
rect 37516 19660 37522 19672
rect 38013 19669 38025 19672
rect 38059 19669 38071 19703
rect 38013 19663 38071 19669
rect 38657 19703 38715 19709
rect 38657 19669 38669 19703
rect 38703 19669 38715 19703
rect 39040 19700 39068 19728
rect 41708 19712 41736 19740
rect 42429 19737 42441 19771
rect 42475 19768 42487 19771
rect 42886 19768 42892 19780
rect 42475 19740 42892 19768
rect 42475 19737 42487 19740
rect 42429 19731 42487 19737
rect 42886 19728 42892 19740
rect 42944 19728 42950 19780
rect 39482 19700 39488 19712
rect 39040 19672 39488 19700
rect 38657 19663 38715 19669
rect 39482 19660 39488 19672
rect 39540 19660 39546 19712
rect 41322 19700 41328 19712
rect 41283 19672 41328 19700
rect 41322 19660 41328 19672
rect 41380 19660 41386 19712
rect 41690 19660 41696 19712
rect 41748 19700 41754 19712
rect 42613 19703 42671 19709
rect 42613 19700 42625 19703
rect 41748 19672 42625 19700
rect 41748 19660 41754 19672
rect 42613 19669 42625 19672
rect 42659 19700 42671 19703
rect 43180 19700 43208 19808
rect 43438 19796 43444 19808
rect 43496 19796 43502 19848
rect 43809 19839 43867 19845
rect 43809 19805 43821 19839
rect 43855 19836 43867 19839
rect 44174 19836 44180 19848
rect 43855 19808 44180 19836
rect 43855 19805 43867 19808
rect 43809 19799 43867 19805
rect 44174 19796 44180 19808
rect 44232 19796 44238 19848
rect 44361 19839 44419 19845
rect 44361 19805 44373 19839
rect 44407 19805 44419 19839
rect 44468 19836 44496 19864
rect 45480 19848 45508 19876
rect 46658 19864 46664 19876
rect 46716 19864 46722 19916
rect 45373 19839 45431 19845
rect 45373 19836 45385 19839
rect 44468 19808 45385 19836
rect 44361 19799 44419 19805
rect 45373 19805 45385 19808
rect 45419 19805 45431 19839
rect 45373 19799 45431 19805
rect 44082 19728 44088 19780
rect 44140 19768 44146 19780
rect 44376 19768 44404 19799
rect 45462 19796 45468 19848
rect 45520 19836 45526 19848
rect 45649 19839 45707 19845
rect 45520 19808 45613 19836
rect 45520 19796 45526 19808
rect 45649 19805 45661 19839
rect 45695 19805 45707 19839
rect 45649 19799 45707 19805
rect 45741 19839 45799 19845
rect 45741 19805 45753 19839
rect 45787 19836 45799 19839
rect 45922 19836 45928 19848
rect 45787 19808 45928 19836
rect 45787 19805 45799 19808
rect 45741 19799 45799 19805
rect 44140 19740 44404 19768
rect 44140 19728 44146 19740
rect 42659 19672 43208 19700
rect 42659 19669 42671 19672
rect 42613 19663 42671 19669
rect 43346 19660 43352 19712
rect 43404 19700 43410 19712
rect 43625 19703 43683 19709
rect 43625 19700 43637 19703
rect 43404 19672 43637 19700
rect 43404 19660 43410 19672
rect 43625 19669 43637 19672
rect 43671 19669 43683 19703
rect 44376 19700 44404 19740
rect 44637 19771 44695 19777
rect 44637 19737 44649 19771
rect 44683 19768 44695 19771
rect 45094 19768 45100 19780
rect 44683 19740 45100 19768
rect 44683 19737 44695 19740
rect 44637 19731 44695 19737
rect 45094 19728 45100 19740
rect 45152 19768 45158 19780
rect 45664 19768 45692 19799
rect 45152 19740 45692 19768
rect 45152 19728 45158 19740
rect 45462 19700 45468 19712
rect 44376 19672 45468 19700
rect 43625 19663 43683 19669
rect 45462 19660 45468 19672
rect 45520 19660 45526 19712
rect 45554 19660 45560 19712
rect 45612 19700 45618 19712
rect 45756 19700 45784 19799
rect 45922 19796 45928 19808
rect 45980 19796 45986 19848
rect 45612 19672 45784 19700
rect 45612 19660 45618 19672
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 23842 19496 23848 19508
rect 23523 19468 23848 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 27249 19499 27307 19505
rect 27249 19496 27261 19499
rect 26660 19468 27261 19496
rect 26660 19456 26666 19468
rect 27249 19465 27261 19468
rect 27295 19465 27307 19499
rect 27249 19459 27307 19465
rect 30190 19456 30196 19508
rect 30248 19496 30254 19508
rect 37461 19499 37519 19505
rect 37461 19496 37473 19499
rect 30248 19468 30512 19496
rect 30248 19456 30254 19468
rect 27614 19428 27620 19440
rect 27172 19400 27620 19428
rect 23658 19360 23664 19372
rect 23619 19332 23664 19360
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 23750 19320 23756 19372
rect 23808 19360 23814 19372
rect 24210 19360 24216 19372
rect 23808 19332 23853 19360
rect 24171 19332 24216 19360
rect 23808 19320 23814 19332
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 24394 19360 24400 19372
rect 24355 19332 24400 19360
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 25314 19360 25320 19372
rect 25227 19332 25320 19360
rect 25314 19320 25320 19332
rect 25372 19360 25378 19372
rect 25682 19360 25688 19372
rect 25372 19332 25688 19360
rect 25372 19320 25378 19332
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 27172 19369 27200 19400
rect 27614 19388 27620 19400
rect 27672 19388 27678 19440
rect 29472 19400 30328 19428
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 27890 19360 27896 19372
rect 27387 19332 27896 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 29472 19369 29500 19400
rect 28629 19363 28687 19369
rect 28629 19329 28641 19363
rect 28675 19360 28687 19363
rect 29273 19363 29331 19369
rect 29273 19360 29285 19363
rect 28675 19332 29285 19360
rect 28675 19329 28687 19332
rect 28629 19323 28687 19329
rect 29273 19329 29285 19332
rect 29319 19329 29331 19363
rect 29273 19323 29331 19329
rect 29457 19363 29515 19369
rect 29457 19329 29469 19363
rect 29503 19329 29515 19363
rect 29457 19323 29515 19329
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 29733 19363 29791 19369
rect 29595 19332 29684 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 23474 19292 23480 19304
rect 23435 19264 23480 19292
rect 23474 19252 23480 19264
rect 23532 19252 23538 19304
rect 25406 19292 25412 19304
rect 25367 19264 25412 19292
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 28718 19252 28724 19304
rect 28776 19292 28782 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28776 19264 28825 19292
rect 28776 19252 28782 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 24302 19156 24308 19168
rect 24263 19128 24308 19156
rect 24302 19116 24308 19128
rect 24360 19116 24366 19168
rect 25685 19159 25743 19165
rect 25685 19125 25697 19159
rect 25731 19156 25743 19159
rect 25774 19156 25780 19168
rect 25731 19128 25780 19156
rect 25731 19125 25743 19128
rect 25685 19119 25743 19125
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 28442 19156 28448 19168
rect 28403 19128 28448 19156
rect 28442 19116 28448 19128
rect 28500 19116 28506 19168
rect 29656 19156 29684 19332
rect 29733 19329 29745 19363
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19360 29883 19363
rect 29914 19360 29920 19372
rect 29871 19332 29920 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 29748 19292 29776 19323
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 30300 19369 30328 19400
rect 30484 19369 30512 19468
rect 32600 19468 37473 19496
rect 30285 19363 30343 19369
rect 30285 19329 30297 19363
rect 30331 19360 30343 19363
rect 30469 19363 30527 19369
rect 30331 19332 30420 19360
rect 30331 19329 30343 19332
rect 30285 19323 30343 19329
rect 30392 19292 30420 19332
rect 30469 19329 30481 19363
rect 30515 19360 30527 19363
rect 31846 19360 31852 19372
rect 30515 19332 31852 19360
rect 30515 19329 30527 19332
rect 30469 19323 30527 19329
rect 31846 19320 31852 19332
rect 31904 19320 31910 19372
rect 32600 19369 32628 19468
rect 37461 19465 37473 19468
rect 37507 19465 37519 19499
rect 37461 19459 37519 19465
rect 37734 19456 37740 19508
rect 37792 19496 37798 19508
rect 38102 19496 38108 19508
rect 37792 19468 38108 19496
rect 37792 19456 37798 19468
rect 38102 19456 38108 19468
rect 38160 19456 38166 19508
rect 38654 19456 38660 19508
rect 38712 19496 38718 19508
rect 39758 19496 39764 19508
rect 38712 19468 39764 19496
rect 38712 19456 38718 19468
rect 39758 19456 39764 19468
rect 39816 19456 39822 19508
rect 40494 19496 40500 19508
rect 40455 19468 40500 19496
rect 40494 19456 40500 19468
rect 40552 19456 40558 19508
rect 40678 19456 40684 19508
rect 40736 19496 40742 19508
rect 43070 19496 43076 19508
rect 40736 19468 43076 19496
rect 40736 19456 40742 19468
rect 43070 19456 43076 19468
rect 43128 19456 43134 19508
rect 43254 19456 43260 19508
rect 43312 19496 43318 19508
rect 44085 19499 44143 19505
rect 44085 19496 44097 19499
rect 43312 19468 44097 19496
rect 43312 19456 43318 19468
rect 44085 19465 44097 19468
rect 44131 19465 44143 19499
rect 44085 19459 44143 19465
rect 44269 19499 44327 19505
rect 44269 19465 44281 19499
rect 44315 19496 44327 19499
rect 45097 19499 45155 19505
rect 45097 19496 45109 19499
rect 44315 19468 45109 19496
rect 44315 19465 44327 19468
rect 44269 19459 44327 19465
rect 45097 19465 45109 19468
rect 45143 19465 45155 19499
rect 46014 19496 46020 19508
rect 45975 19468 46020 19496
rect 45097 19459 45155 19465
rect 46014 19456 46020 19468
rect 46072 19456 46078 19508
rect 33226 19428 33232 19440
rect 32692 19400 33232 19428
rect 32692 19369 32720 19400
rect 33226 19388 33232 19400
rect 33284 19388 33290 19440
rect 35986 19428 35992 19440
rect 34348 19400 35992 19428
rect 32585 19363 32643 19369
rect 32585 19329 32597 19363
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 32677 19363 32735 19369
rect 32677 19329 32689 19363
rect 32723 19329 32735 19363
rect 32677 19323 32735 19329
rect 32953 19363 33011 19369
rect 32953 19329 32965 19363
rect 32999 19360 33011 19363
rect 33318 19360 33324 19372
rect 32999 19332 33324 19360
rect 32999 19329 33011 19332
rect 32953 19323 33011 19329
rect 33318 19320 33324 19332
rect 33376 19320 33382 19372
rect 34348 19369 34376 19400
rect 35986 19388 35992 19400
rect 36044 19388 36050 19440
rect 36078 19388 36084 19440
rect 36136 19428 36142 19440
rect 36817 19431 36875 19437
rect 36817 19428 36829 19431
rect 36136 19400 36829 19428
rect 36136 19388 36142 19400
rect 36817 19397 36829 19400
rect 36863 19397 36875 19431
rect 36817 19391 36875 19397
rect 37366 19388 37372 19440
rect 37424 19428 37430 19440
rect 40218 19428 40224 19440
rect 37424 19400 40224 19428
rect 37424 19388 37430 19400
rect 34333 19363 34391 19369
rect 34333 19329 34345 19363
rect 34379 19329 34391 19363
rect 34333 19323 34391 19329
rect 34422 19320 34428 19372
rect 34480 19360 34486 19372
rect 34609 19363 34667 19369
rect 34480 19332 34525 19360
rect 34609 19338 34621 19363
rect 34655 19338 34667 19363
rect 35342 19360 35348 19372
rect 34480 19320 34486 19332
rect 32401 19295 32459 19301
rect 32401 19292 32413 19295
rect 29748 19264 30328 19292
rect 30392 19264 32413 19292
rect 30300 19233 30328 19264
rect 32401 19261 32413 19264
rect 32447 19261 32459 19295
rect 34514 19292 34520 19304
rect 34475 19264 34520 19292
rect 32401 19255 32459 19261
rect 34514 19252 34520 19264
rect 34572 19252 34578 19304
rect 34606 19286 34612 19338
rect 34664 19334 34670 19338
rect 34664 19306 34723 19334
rect 35303 19332 35348 19360
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 35434 19320 35440 19372
rect 35492 19360 35498 19372
rect 35492 19332 35537 19360
rect 35492 19320 35498 19332
rect 35802 19320 35808 19372
rect 35860 19360 35866 19372
rect 36354 19360 36360 19372
rect 35860 19332 36216 19360
rect 36315 19332 36360 19360
rect 35860 19320 35866 19332
rect 34664 19286 34670 19306
rect 35529 19295 35587 19301
rect 35529 19292 35541 19295
rect 35360 19264 35541 19292
rect 30285 19227 30343 19233
rect 30285 19193 30297 19227
rect 30331 19193 30343 19227
rect 30285 19187 30343 19193
rect 31386 19184 31392 19236
rect 31444 19224 31450 19236
rect 31481 19227 31539 19233
rect 31481 19224 31493 19227
rect 31444 19196 31493 19224
rect 31444 19184 31450 19196
rect 31481 19193 31493 19196
rect 31527 19193 31539 19227
rect 32858 19224 32864 19236
rect 32819 19196 32864 19224
rect 31481 19187 31539 19193
rect 32858 19184 32864 19196
rect 32916 19184 32922 19236
rect 30558 19156 30564 19168
rect 29656 19128 30564 19156
rect 30558 19116 30564 19128
rect 30616 19116 30622 19168
rect 33318 19116 33324 19168
rect 33376 19156 33382 19168
rect 33413 19159 33471 19165
rect 33413 19156 33425 19159
rect 33376 19128 33425 19156
rect 33376 19116 33382 19128
rect 33413 19125 33425 19128
rect 33459 19125 33471 19159
rect 33413 19119 33471 19125
rect 34149 19159 34207 19165
rect 34149 19125 34161 19159
rect 34195 19156 34207 19159
rect 34330 19156 34336 19168
rect 34195 19128 34336 19156
rect 34195 19125 34207 19128
rect 34149 19119 34207 19125
rect 34330 19116 34336 19128
rect 34388 19116 34394 19168
rect 35161 19159 35219 19165
rect 35161 19125 35173 19159
rect 35207 19156 35219 19159
rect 35250 19156 35256 19168
rect 35207 19128 35256 19156
rect 35207 19125 35219 19128
rect 35161 19119 35219 19125
rect 35250 19116 35256 19128
rect 35308 19116 35314 19168
rect 35360 19156 35388 19264
rect 35529 19261 35541 19264
rect 35575 19261 35587 19295
rect 35529 19255 35587 19261
rect 35621 19295 35679 19301
rect 35621 19261 35633 19295
rect 35667 19292 35679 19295
rect 35986 19292 35992 19304
rect 35667 19264 35992 19292
rect 35667 19261 35679 19264
rect 35621 19255 35679 19261
rect 35986 19252 35992 19264
rect 36044 19252 36050 19304
rect 36188 19233 36216 19332
rect 36354 19320 36360 19332
rect 36412 19320 36418 19372
rect 36541 19363 36599 19369
rect 36541 19329 36553 19363
rect 36587 19360 36599 19363
rect 36630 19360 36636 19372
rect 36587 19332 36636 19360
rect 36587 19329 36599 19332
rect 36541 19323 36599 19329
rect 36630 19320 36636 19332
rect 36688 19320 36694 19372
rect 37734 19360 37740 19372
rect 37384 19332 37740 19360
rect 37384 19304 37412 19332
rect 37734 19320 37740 19332
rect 37792 19320 37798 19372
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 37366 19252 37372 19304
rect 37424 19252 37430 19304
rect 37844 19292 37872 19323
rect 37918 19320 37924 19372
rect 37976 19360 37982 19372
rect 38120 19369 38148 19400
rect 40218 19388 40224 19400
rect 40276 19388 40282 19440
rect 41509 19431 41567 19437
rect 41509 19428 41521 19431
rect 40604 19400 41521 19428
rect 38105 19363 38163 19369
rect 37976 19332 38021 19360
rect 37976 19320 37982 19332
rect 38105 19329 38117 19363
rect 38151 19329 38163 19363
rect 38105 19323 38163 19329
rect 38930 19320 38936 19372
rect 38988 19360 38994 19372
rect 39117 19363 39175 19369
rect 39117 19360 39129 19363
rect 38988 19332 39129 19360
rect 38988 19320 38994 19332
rect 39117 19329 39129 19332
rect 39163 19329 39175 19363
rect 39117 19323 39175 19329
rect 39209 19363 39267 19369
rect 39209 19329 39221 19363
rect 39255 19329 39267 19363
rect 39209 19323 39267 19329
rect 38194 19292 38200 19304
rect 37844 19264 38200 19292
rect 38194 19252 38200 19264
rect 38252 19292 38258 19304
rect 39224 19292 39252 19323
rect 39298 19320 39304 19372
rect 39356 19360 39362 19372
rect 39356 19332 39401 19360
rect 39356 19320 39362 19332
rect 39482 19320 39488 19372
rect 39540 19360 39546 19372
rect 39540 19332 39585 19360
rect 39540 19320 39546 19332
rect 40310 19320 40316 19372
rect 40368 19360 40374 19372
rect 40604 19369 40632 19400
rect 41509 19397 41521 19400
rect 41555 19397 41567 19431
rect 42058 19428 42064 19440
rect 42019 19400 42064 19428
rect 41509 19391 41567 19397
rect 42058 19388 42064 19400
rect 42116 19388 42122 19440
rect 43162 19428 43168 19440
rect 43075 19400 43168 19428
rect 40405 19363 40463 19369
rect 40405 19360 40417 19363
rect 40368 19332 40417 19360
rect 40368 19320 40374 19332
rect 40405 19329 40417 19332
rect 40451 19329 40463 19363
rect 40405 19323 40463 19329
rect 40589 19363 40647 19369
rect 40589 19329 40601 19363
rect 40635 19329 40647 19363
rect 40589 19323 40647 19329
rect 40862 19320 40868 19372
rect 40920 19360 40926 19372
rect 41233 19363 41291 19369
rect 41233 19360 41245 19363
rect 40920 19332 41245 19360
rect 40920 19320 40926 19332
rect 41233 19329 41245 19332
rect 41279 19329 41291 19363
rect 41233 19323 41291 19329
rect 41874 19320 41880 19372
rect 41932 19360 41938 19372
rect 42426 19360 42432 19372
rect 41932 19332 42432 19360
rect 41932 19320 41938 19332
rect 42426 19320 42432 19332
rect 42484 19360 42490 19372
rect 42702 19360 42708 19372
rect 42484 19332 42708 19360
rect 42484 19320 42490 19332
rect 42702 19320 42708 19332
rect 42760 19320 42766 19372
rect 43088 19369 43116 19400
rect 43162 19388 43168 19400
rect 43220 19428 43226 19440
rect 43346 19428 43352 19440
rect 43220 19400 43352 19428
rect 43220 19388 43226 19400
rect 43346 19388 43352 19400
rect 43404 19388 43410 19440
rect 43438 19388 43444 19440
rect 43496 19428 43502 19440
rect 46032 19428 46060 19456
rect 43496 19400 44220 19428
rect 43496 19388 43502 19400
rect 43073 19363 43131 19369
rect 43073 19329 43085 19363
rect 43119 19329 43131 19363
rect 43254 19360 43260 19372
rect 43215 19332 43260 19360
rect 43073 19323 43131 19329
rect 43254 19320 43260 19332
rect 43312 19320 43318 19372
rect 43898 19360 43904 19372
rect 43859 19332 43904 19360
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 44192 19360 44220 19400
rect 45388 19400 46060 19428
rect 45388 19360 45416 19400
rect 44192 19332 45416 19360
rect 41414 19292 41420 19304
rect 38252 19264 41420 19292
rect 38252 19252 38258 19264
rect 41414 19252 41420 19264
rect 41472 19252 41478 19304
rect 41506 19252 41512 19304
rect 41564 19292 41570 19304
rect 41564 19264 41609 19292
rect 41564 19252 41570 19264
rect 41782 19252 41788 19304
rect 41840 19292 41846 19304
rect 43993 19295 44051 19301
rect 41840 19264 43944 19292
rect 41840 19252 41846 19264
rect 36173 19227 36231 19233
rect 36173 19193 36185 19227
rect 36219 19193 36231 19227
rect 36173 19187 36231 19193
rect 36630 19184 36636 19236
rect 36688 19224 36694 19236
rect 36688 19196 41000 19224
rect 36688 19184 36694 19196
rect 36446 19156 36452 19168
rect 35360 19128 36452 19156
rect 36446 19116 36452 19128
rect 36504 19116 36510 19168
rect 36725 19159 36783 19165
rect 36725 19125 36737 19159
rect 36771 19156 36783 19159
rect 37550 19156 37556 19168
rect 36771 19128 37556 19156
rect 36771 19125 36783 19128
rect 36725 19119 36783 19125
rect 37550 19116 37556 19128
rect 37608 19116 37614 19168
rect 37918 19116 37924 19168
rect 37976 19156 37982 19168
rect 38378 19156 38384 19168
rect 37976 19128 38384 19156
rect 37976 19116 37982 19128
rect 38378 19116 38384 19128
rect 38436 19116 38442 19168
rect 38838 19156 38844 19168
rect 38799 19128 38844 19156
rect 38838 19116 38844 19128
rect 38896 19116 38902 19168
rect 40972 19156 41000 19196
rect 41046 19184 41052 19236
rect 41104 19224 41110 19236
rect 43717 19227 43775 19233
rect 43717 19224 43729 19227
rect 41104 19196 43729 19224
rect 41104 19184 41110 19196
rect 43717 19193 43729 19196
rect 43763 19193 43775 19227
rect 43916 19224 43944 19264
rect 43993 19261 44005 19295
rect 44039 19292 44051 19295
rect 44192 19292 44220 19332
rect 45388 19304 45416 19332
rect 45557 19363 45615 19369
rect 45557 19329 45569 19363
rect 45603 19360 45615 19363
rect 45830 19360 45836 19372
rect 45603 19332 45836 19360
rect 45603 19329 45615 19332
rect 45557 19323 45615 19329
rect 45830 19320 45836 19332
rect 45888 19320 45894 19372
rect 44039 19264 44220 19292
rect 44361 19295 44419 19301
rect 44039 19261 44051 19264
rect 43993 19255 44051 19261
rect 44361 19261 44373 19295
rect 44407 19261 44419 19295
rect 44361 19255 44419 19261
rect 44266 19224 44272 19236
rect 43916 19196 44272 19224
rect 43717 19187 43775 19193
rect 44266 19184 44272 19196
rect 44324 19224 44330 19236
rect 44376 19224 44404 19255
rect 45370 19252 45376 19304
rect 45428 19252 45434 19304
rect 44324 19196 44404 19224
rect 44324 19184 44330 19196
rect 41325 19159 41383 19165
rect 41325 19156 41337 19159
rect 40972 19128 41337 19156
rect 41325 19125 41337 19128
rect 41371 19156 41383 19159
rect 41782 19156 41788 19168
rect 41371 19128 41788 19156
rect 41371 19125 41383 19128
rect 41325 19119 41383 19125
rect 41782 19116 41788 19128
rect 41840 19116 41846 19168
rect 43070 19156 43076 19168
rect 43031 19128 43076 19156
rect 43070 19116 43076 19128
rect 43128 19156 43134 19168
rect 44082 19156 44088 19168
rect 43128 19128 44088 19156
rect 43128 19116 43134 19128
rect 44082 19116 44088 19128
rect 44140 19116 44146 19168
rect 44910 19116 44916 19168
rect 44968 19156 44974 19168
rect 45278 19156 45284 19168
rect 44968 19128 45284 19156
rect 44968 19116 44974 19128
rect 45278 19116 45284 19128
rect 45336 19116 45342 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 23569 18955 23627 18961
rect 23569 18952 23581 18955
rect 23532 18924 23581 18952
rect 23532 18912 23538 18924
rect 23569 18921 23581 18924
rect 23615 18921 23627 18955
rect 25958 18952 25964 18964
rect 25919 18924 25964 18952
rect 23569 18915 23627 18921
rect 25958 18912 25964 18924
rect 26016 18912 26022 18964
rect 27614 18952 27620 18964
rect 27575 18924 27620 18952
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 27816 18924 31754 18952
rect 27816 18896 27844 18924
rect 27798 18884 27804 18896
rect 27711 18856 27804 18884
rect 27798 18844 27804 18856
rect 27856 18844 27862 18896
rect 31726 18884 31754 18924
rect 33042 18912 33048 18964
rect 33100 18952 33106 18964
rect 35437 18955 35495 18961
rect 35437 18952 35449 18955
rect 33100 18924 35449 18952
rect 33100 18912 33106 18924
rect 35437 18921 35449 18924
rect 35483 18921 35495 18955
rect 35437 18915 35495 18921
rect 36078 18912 36084 18964
rect 36136 18952 36142 18964
rect 36173 18955 36231 18961
rect 36173 18952 36185 18955
rect 36136 18924 36185 18952
rect 36136 18912 36142 18924
rect 36173 18921 36185 18924
rect 36219 18921 36231 18955
rect 39022 18952 39028 18964
rect 36173 18915 36231 18921
rect 36280 18924 39028 18952
rect 34885 18887 34943 18893
rect 34885 18884 34897 18887
rect 31726 18856 34897 18884
rect 34885 18853 34897 18856
rect 34931 18853 34943 18887
rect 34885 18847 34943 18853
rect 35526 18844 35532 18896
rect 35584 18884 35590 18896
rect 36280 18884 36308 18924
rect 39022 18912 39028 18924
rect 39080 18912 39086 18964
rect 39298 18912 39304 18964
rect 39356 18952 39362 18964
rect 39485 18955 39543 18961
rect 39485 18952 39497 18955
rect 39356 18924 39497 18952
rect 39356 18912 39362 18924
rect 39485 18921 39497 18924
rect 39531 18921 39543 18955
rect 39485 18915 39543 18921
rect 41064 18924 41460 18952
rect 35584 18856 36308 18884
rect 35584 18844 35590 18856
rect 36354 18844 36360 18896
rect 36412 18884 36418 18896
rect 36630 18884 36636 18896
rect 36412 18856 36636 18884
rect 36412 18844 36418 18856
rect 36630 18844 36636 18856
rect 36688 18844 36694 18896
rect 37458 18884 37464 18896
rect 37419 18856 37464 18884
rect 37458 18844 37464 18856
rect 37516 18844 37522 18896
rect 37553 18887 37611 18893
rect 37553 18853 37565 18887
rect 37599 18884 37611 18887
rect 38194 18884 38200 18896
rect 37599 18856 38200 18884
rect 37599 18853 37611 18856
rect 37553 18847 37611 18853
rect 38194 18844 38200 18856
rect 38252 18844 38258 18896
rect 38930 18844 38936 18896
rect 38988 18884 38994 18896
rect 41064 18884 41092 18924
rect 38988 18856 41092 18884
rect 38988 18844 38994 18856
rect 41138 18844 41144 18896
rect 41196 18844 41202 18896
rect 41432 18884 41460 18924
rect 41506 18912 41512 18964
rect 41564 18952 41570 18964
rect 42426 18952 42432 18964
rect 41564 18924 42432 18952
rect 41564 18912 41570 18924
rect 42426 18912 42432 18924
rect 42484 18952 42490 18964
rect 42705 18955 42763 18961
rect 42705 18952 42717 18955
rect 42484 18924 42717 18952
rect 42484 18912 42490 18924
rect 42705 18921 42717 18924
rect 42751 18921 42763 18955
rect 42705 18915 42763 18921
rect 44174 18912 44180 18964
rect 44232 18952 44238 18964
rect 44361 18955 44419 18961
rect 44361 18952 44373 18955
rect 44232 18924 44373 18952
rect 44232 18912 44238 18924
rect 44361 18921 44373 18924
rect 44407 18921 44419 18955
rect 44361 18915 44419 18921
rect 46106 18912 46112 18964
rect 46164 18952 46170 18964
rect 46201 18955 46259 18961
rect 46201 18952 46213 18955
rect 46164 18924 46213 18952
rect 46164 18912 46170 18924
rect 46201 18921 46213 18924
rect 46247 18921 46259 18955
rect 46201 18915 46259 18921
rect 43438 18884 43444 18896
rect 41432 18856 42104 18884
rect 43399 18856 43444 18884
rect 23385 18819 23443 18825
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 23566 18816 23572 18828
rect 23431 18788 23572 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 23566 18776 23572 18788
rect 23624 18816 23630 18828
rect 28442 18816 28448 18828
rect 23624 18788 28448 18816
rect 23624 18776 23630 18788
rect 28442 18776 28448 18788
rect 28500 18776 28506 18828
rect 31754 18816 31760 18828
rect 31036 18788 31760 18816
rect 31036 18760 31064 18788
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 33965 18819 34023 18825
rect 33965 18816 33977 18819
rect 32232 18788 33977 18816
rect 32232 18760 32260 18788
rect 33965 18785 33977 18788
rect 34011 18785 34023 18819
rect 37185 18819 37243 18825
rect 37185 18816 37197 18819
rect 33965 18779 34023 18785
rect 34164 18788 37197 18816
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18748 23351 18751
rect 24302 18748 24308 18760
rect 23339 18720 24308 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24636 18720 24777 18748
rect 24636 18708 24642 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18748 25007 18751
rect 25038 18748 25044 18760
rect 24995 18720 25044 18748
rect 24995 18717 25007 18720
rect 24949 18711 25007 18717
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 25774 18748 25780 18760
rect 25735 18720 25780 18748
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 25958 18748 25964 18760
rect 25919 18720 25964 18748
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 31018 18748 31024 18760
rect 30979 18720 31024 18748
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 31113 18751 31171 18757
rect 31113 18717 31125 18751
rect 31159 18717 31171 18751
rect 31113 18711 31171 18717
rect 31205 18751 31263 18757
rect 31205 18717 31217 18751
rect 31251 18717 31263 18751
rect 31386 18748 31392 18760
rect 31347 18720 31392 18748
rect 31205 18711 31263 18717
rect 28074 18680 28080 18692
rect 28035 18652 28080 18680
rect 28074 18640 28080 18652
rect 28132 18680 28138 18692
rect 28537 18683 28595 18689
rect 28537 18680 28549 18683
rect 28132 18652 28549 18680
rect 28132 18640 28138 18652
rect 28537 18649 28549 18652
rect 28583 18649 28595 18683
rect 28537 18643 28595 18649
rect 31128 18624 31156 18711
rect 31220 18680 31248 18711
rect 31386 18708 31392 18720
rect 31444 18708 31450 18760
rect 32214 18748 32220 18760
rect 32127 18720 32220 18748
rect 32214 18708 32220 18720
rect 32272 18708 32278 18760
rect 33042 18748 33048 18760
rect 33003 18720 33048 18748
rect 33042 18708 33048 18720
rect 33100 18708 33106 18760
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18748 33195 18751
rect 33594 18748 33600 18760
rect 33183 18720 33600 18748
rect 33183 18717 33195 18720
rect 33137 18711 33195 18717
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 34164 18757 34192 18788
rect 37185 18785 37197 18788
rect 37231 18785 37243 18819
rect 37185 18779 37243 18785
rect 37918 18776 37924 18828
rect 37976 18816 37982 18828
rect 38838 18816 38844 18828
rect 37976 18788 38844 18816
rect 37976 18776 37982 18788
rect 38838 18776 38844 18788
rect 38896 18776 38902 18828
rect 39482 18776 39488 18828
rect 39540 18816 39546 18828
rect 41156 18816 41184 18844
rect 41233 18819 41291 18825
rect 41233 18816 41245 18819
rect 39540 18788 41245 18816
rect 39540 18776 39546 18788
rect 41233 18785 41245 18788
rect 41279 18785 41291 18819
rect 41874 18816 41880 18828
rect 41835 18788 41880 18816
rect 41233 18779 41291 18785
rect 41874 18776 41880 18788
rect 41932 18776 41938 18828
rect 34149 18751 34207 18757
rect 34149 18717 34161 18751
rect 34195 18717 34207 18751
rect 34330 18748 34336 18760
rect 34291 18720 34336 18748
rect 34149 18711 34207 18717
rect 34330 18708 34336 18720
rect 34388 18708 34394 18760
rect 34606 18708 34612 18760
rect 34664 18748 34670 18760
rect 35010 18751 35068 18757
rect 35010 18748 35022 18751
rect 34664 18720 35022 18748
rect 34664 18708 34670 18720
rect 35010 18717 35022 18720
rect 35056 18717 35068 18751
rect 35526 18748 35532 18760
rect 35487 18720 35532 18748
rect 35010 18711 35068 18717
rect 35526 18708 35532 18720
rect 35584 18708 35590 18760
rect 37375 18705 37381 18757
rect 37433 18742 37439 18757
rect 37642 18748 37648 18760
rect 37433 18714 37475 18742
rect 37603 18720 37648 18748
rect 37433 18705 37439 18714
rect 37642 18708 37648 18720
rect 37700 18708 37706 18760
rect 37734 18708 37740 18760
rect 37792 18748 37798 18760
rect 40770 18757 40776 18760
rect 37829 18751 37887 18757
rect 37829 18748 37841 18751
rect 37792 18720 37841 18748
rect 37792 18708 37798 18720
rect 37829 18717 37841 18720
rect 37875 18717 37887 18751
rect 40742 18751 40776 18757
rect 40742 18748 40754 18751
rect 37829 18711 37887 18717
rect 37936 18720 40264 18748
rect 31849 18683 31907 18689
rect 31849 18680 31861 18683
rect 31220 18652 31861 18680
rect 31849 18649 31861 18652
rect 31895 18649 31907 18683
rect 32030 18680 32036 18692
rect 31991 18652 32036 18680
rect 31849 18643 31907 18649
rect 32030 18640 32036 18652
rect 32088 18640 32094 18692
rect 33318 18640 33324 18692
rect 33376 18680 33382 18692
rect 33413 18683 33471 18689
rect 33413 18680 33425 18683
rect 33376 18652 33425 18680
rect 33376 18640 33382 18652
rect 33413 18649 33425 18652
rect 33459 18649 33471 18683
rect 33413 18643 33471 18649
rect 33505 18683 33563 18689
rect 33505 18649 33517 18683
rect 33551 18680 33563 18683
rect 36357 18683 36415 18689
rect 33551 18652 36308 18680
rect 33551 18649 33563 18652
rect 33505 18643 33563 18649
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24210 18612 24216 18624
rect 23900 18584 24216 18612
rect 23900 18572 23906 18584
rect 24210 18572 24216 18584
rect 24268 18612 24274 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 24268 18584 24593 18612
rect 24268 18572 24274 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 30745 18615 30803 18621
rect 30745 18612 30757 18615
rect 25648 18584 30757 18612
rect 25648 18572 25654 18584
rect 30745 18581 30757 18584
rect 30791 18581 30803 18615
rect 30745 18575 30803 18581
rect 31110 18572 31116 18624
rect 31168 18572 31174 18624
rect 32674 18572 32680 18624
rect 32732 18612 32738 18624
rect 32861 18615 32919 18621
rect 32861 18612 32873 18615
rect 32732 18584 32873 18612
rect 32732 18572 32738 18584
rect 32861 18581 32873 18584
rect 32907 18581 32919 18615
rect 32861 18575 32919 18581
rect 35069 18615 35127 18621
rect 35069 18581 35081 18615
rect 35115 18612 35127 18615
rect 35342 18612 35348 18624
rect 35115 18584 35348 18612
rect 35115 18581 35127 18584
rect 35069 18575 35127 18581
rect 35342 18572 35348 18584
rect 35400 18572 35406 18624
rect 36280 18612 36308 18652
rect 36357 18649 36369 18683
rect 36403 18680 36415 18683
rect 36446 18680 36452 18692
rect 36403 18652 36452 18680
rect 36403 18649 36415 18652
rect 36357 18643 36415 18649
rect 36446 18640 36452 18652
rect 36504 18640 36510 18692
rect 36541 18683 36599 18689
rect 36541 18649 36553 18683
rect 36587 18680 36599 18683
rect 36630 18680 36636 18692
rect 36587 18652 36636 18680
rect 36587 18649 36599 18652
rect 36541 18643 36599 18649
rect 36630 18640 36636 18652
rect 36688 18640 36694 18692
rect 37936 18612 37964 18720
rect 38378 18640 38384 18692
rect 38436 18680 38442 18692
rect 39117 18683 39175 18689
rect 39117 18680 39129 18683
rect 38436 18652 39129 18680
rect 38436 18640 38442 18652
rect 39117 18649 39129 18652
rect 39163 18649 39175 18683
rect 39117 18643 39175 18649
rect 39206 18640 39212 18692
rect 39264 18680 39270 18692
rect 39301 18683 39359 18689
rect 39301 18680 39313 18683
rect 39264 18652 39313 18680
rect 39264 18640 39270 18652
rect 39301 18649 39313 18652
rect 39347 18649 39359 18683
rect 39301 18643 39359 18649
rect 36280 18584 37964 18612
rect 38194 18572 38200 18624
rect 38252 18612 38258 18624
rect 38562 18612 38568 18624
rect 38252 18584 38568 18612
rect 38252 18572 38258 18584
rect 38562 18572 38568 18584
rect 38620 18612 38626 18624
rect 38657 18615 38715 18621
rect 38657 18612 38669 18615
rect 38620 18584 38669 18612
rect 38620 18572 38626 18584
rect 38657 18581 38669 18584
rect 38703 18581 38715 18615
rect 38657 18575 38715 18581
rect 39022 18572 39028 18624
rect 39080 18612 39086 18624
rect 40037 18615 40095 18621
rect 40037 18612 40049 18615
rect 39080 18584 40049 18612
rect 39080 18572 39086 18584
rect 40037 18581 40049 18584
rect 40083 18581 40095 18615
rect 40236 18612 40264 18720
rect 40684 18720 40754 18748
rect 40494 18640 40500 18692
rect 40552 18680 40558 18692
rect 40684 18680 40712 18720
rect 40742 18717 40754 18720
rect 40828 18748 40834 18760
rect 40828 18720 40890 18748
rect 40742 18711 40776 18717
rect 40770 18708 40776 18711
rect 40828 18708 40834 18720
rect 41046 18708 41052 18760
rect 41104 18748 41110 18760
rect 41141 18751 41199 18757
rect 41141 18748 41153 18751
rect 41104 18720 41153 18748
rect 41104 18708 41110 18720
rect 41141 18717 41153 18720
rect 41187 18717 41199 18751
rect 42076 18748 42104 18856
rect 43438 18844 43444 18856
rect 43496 18844 43502 18896
rect 44266 18844 44272 18896
rect 44324 18884 44330 18896
rect 45281 18887 45339 18893
rect 45281 18884 45293 18887
rect 44324 18856 45293 18884
rect 44324 18844 44330 18856
rect 45281 18853 45293 18856
rect 45327 18853 45339 18887
rect 45281 18847 45339 18853
rect 42794 18816 42800 18828
rect 42352 18788 42800 18816
rect 42352 18757 42380 18788
rect 42794 18776 42800 18788
rect 42852 18776 42858 18828
rect 43165 18819 43223 18825
rect 43165 18785 43177 18819
rect 43211 18785 43223 18819
rect 43714 18816 43720 18828
rect 43165 18779 43223 18785
rect 43364 18788 43720 18816
rect 42337 18751 42395 18757
rect 42337 18748 42349 18751
rect 41141 18711 41199 18717
rect 41616 18720 42012 18748
rect 42076 18720 42349 18748
rect 41616 18680 41644 18720
rect 40552 18652 40712 18680
rect 41386 18652 41644 18680
rect 41984 18680 42012 18720
rect 42337 18717 42349 18720
rect 42383 18717 42395 18751
rect 43180 18748 43208 18779
rect 43364 18757 43392 18788
rect 43714 18776 43720 18788
rect 43772 18776 43778 18828
rect 46124 18816 46152 18912
rect 44468 18788 46152 18816
rect 42337 18711 42395 18717
rect 42444 18720 43208 18748
rect 43349 18751 43407 18757
rect 42444 18680 42472 18720
rect 43349 18717 43361 18751
rect 43395 18717 43407 18751
rect 43349 18711 43407 18717
rect 43533 18751 43591 18757
rect 43533 18717 43545 18751
rect 43579 18717 43591 18751
rect 43533 18711 43591 18717
rect 41984 18652 42472 18680
rect 40552 18640 40558 18652
rect 40589 18615 40647 18621
rect 40589 18612 40601 18615
rect 40236 18584 40601 18612
rect 40037 18575 40095 18581
rect 40589 18581 40601 18584
rect 40635 18581 40647 18615
rect 40589 18575 40647 18581
rect 40773 18615 40831 18621
rect 40773 18581 40785 18615
rect 40819 18612 40831 18615
rect 41386 18612 41414 18652
rect 42518 18640 42524 18692
rect 42576 18680 42582 18692
rect 42576 18652 42621 18680
rect 42576 18640 42582 18652
rect 43548 18624 43576 18711
rect 43622 18708 43628 18760
rect 43680 18748 43686 18760
rect 43680 18720 43725 18748
rect 43680 18708 43686 18720
rect 43806 18708 43812 18760
rect 43864 18748 43870 18760
rect 44468 18757 44496 18788
rect 44453 18751 44511 18757
rect 43864 18720 43909 18748
rect 43864 18708 43870 18720
rect 44453 18717 44465 18751
rect 44499 18717 44511 18751
rect 44453 18711 44511 18717
rect 44910 18708 44916 18760
rect 44968 18748 44974 18760
rect 45189 18751 45247 18757
rect 45189 18748 45201 18751
rect 44968 18720 45201 18748
rect 44968 18708 44974 18720
rect 45189 18717 45201 18720
rect 45235 18717 45247 18751
rect 45189 18711 45247 18717
rect 45649 18751 45707 18757
rect 45649 18717 45661 18751
rect 45695 18748 45707 18751
rect 45830 18748 45836 18760
rect 45695 18720 45836 18748
rect 45695 18717 45707 18720
rect 45649 18711 45707 18717
rect 45830 18708 45836 18720
rect 45888 18708 45894 18760
rect 40819 18584 41414 18612
rect 40819 18581 40831 18584
rect 40773 18575 40831 18581
rect 41506 18572 41512 18624
rect 41564 18612 41570 18624
rect 43530 18612 43536 18624
rect 41564 18584 43536 18612
rect 41564 18572 41570 18584
rect 43530 18572 43536 18584
rect 43588 18572 43594 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 30361 18411 30419 18417
rect 30361 18377 30373 18411
rect 30407 18408 30419 18411
rect 32122 18408 32128 18420
rect 30407 18380 32128 18408
rect 30407 18377 30419 18380
rect 30361 18371 30419 18377
rect 32122 18368 32128 18380
rect 32180 18368 32186 18420
rect 33226 18408 33232 18420
rect 33187 18380 33232 18408
rect 33226 18368 33232 18380
rect 33284 18368 33290 18420
rect 34698 18368 34704 18420
rect 34756 18408 34762 18420
rect 37826 18408 37832 18420
rect 34756 18380 34928 18408
rect 34756 18368 34762 18380
rect 30558 18340 30564 18352
rect 30519 18312 30564 18340
rect 30558 18300 30564 18312
rect 30616 18300 30622 18352
rect 31110 18340 31116 18352
rect 31071 18312 31116 18340
rect 31110 18300 31116 18312
rect 31168 18300 31174 18352
rect 34054 18340 34060 18352
rect 32784 18312 34060 18340
rect 23566 18272 23572 18284
rect 23527 18244 23572 18272
rect 23566 18232 23572 18244
rect 23624 18232 23630 18284
rect 23842 18272 23848 18284
rect 23803 18244 23848 18272
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 24394 18232 24400 18284
rect 24452 18272 24458 18284
rect 24581 18275 24639 18281
rect 24581 18272 24593 18275
rect 24452 18244 24593 18272
rect 24452 18232 24458 18244
rect 24581 18241 24593 18244
rect 24627 18241 24639 18275
rect 24581 18235 24639 18241
rect 25685 18275 25743 18281
rect 25685 18241 25697 18275
rect 25731 18272 25743 18275
rect 25774 18272 25780 18284
rect 25731 18244 25780 18272
rect 25731 18241 25743 18244
rect 25685 18235 25743 18241
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 27522 18272 27528 18284
rect 27483 18244 27528 18272
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 28997 18275 29055 18281
rect 28997 18241 29009 18275
rect 29043 18272 29055 18275
rect 29914 18272 29920 18284
rect 29043 18244 29920 18272
rect 29043 18241 29055 18244
rect 28997 18235 29055 18241
rect 29914 18232 29920 18244
rect 29972 18232 29978 18284
rect 31389 18275 31447 18281
rect 31389 18241 31401 18275
rect 31435 18272 31447 18275
rect 32030 18272 32036 18284
rect 31435 18244 32036 18272
rect 31435 18241 31447 18244
rect 31389 18235 31447 18241
rect 32030 18232 32036 18244
rect 32088 18272 32094 18284
rect 32490 18272 32496 18284
rect 32088 18244 32496 18272
rect 32088 18232 32094 18244
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 32784 18281 32812 18312
rect 34054 18300 34060 18312
rect 34112 18300 34118 18352
rect 32769 18275 32827 18281
rect 32769 18241 32781 18275
rect 32815 18241 32827 18275
rect 32769 18235 32827 18241
rect 33229 18275 33287 18281
rect 33229 18241 33241 18275
rect 33275 18272 33287 18275
rect 33318 18272 33324 18284
rect 33275 18244 33324 18272
rect 33275 18241 33287 18244
rect 33229 18235 33287 18241
rect 25593 18207 25651 18213
rect 25593 18173 25605 18207
rect 25639 18173 25651 18207
rect 25593 18167 25651 18173
rect 27617 18207 27675 18213
rect 27617 18173 27629 18207
rect 27663 18204 27675 18207
rect 27798 18204 27804 18216
rect 27663 18176 27804 18204
rect 27663 18173 27675 18176
rect 27617 18167 27675 18173
rect 24302 18136 24308 18148
rect 24263 18108 24308 18136
rect 24302 18096 24308 18108
rect 24360 18096 24366 18148
rect 25608 18136 25636 18167
rect 27798 18164 27804 18176
rect 27856 18164 27862 18216
rect 28718 18204 28724 18216
rect 28679 18176 28724 18204
rect 28718 18164 28724 18176
rect 28776 18164 28782 18216
rect 31113 18207 31171 18213
rect 31113 18173 31125 18207
rect 31159 18204 31171 18207
rect 32214 18204 32220 18216
rect 31159 18176 32220 18204
rect 31159 18173 31171 18176
rect 31113 18167 31171 18173
rect 32214 18164 32220 18176
rect 32272 18164 32278 18216
rect 25958 18136 25964 18148
rect 25608 18108 25964 18136
rect 25958 18096 25964 18108
rect 26016 18136 26022 18148
rect 28813 18139 28871 18145
rect 28813 18136 28825 18139
rect 26016 18108 28825 18136
rect 26016 18096 26022 18108
rect 28813 18105 28825 18108
rect 28859 18105 28871 18139
rect 31938 18136 31944 18148
rect 28813 18099 28871 18105
rect 30392 18108 31944 18136
rect 25317 18071 25375 18077
rect 25317 18037 25329 18071
rect 25363 18068 25375 18071
rect 25498 18068 25504 18080
rect 25363 18040 25504 18068
rect 25363 18037 25375 18040
rect 25317 18031 25375 18037
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 27246 18068 27252 18080
rect 27207 18040 27252 18068
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 28905 18071 28963 18077
rect 28905 18037 28917 18071
rect 28951 18068 28963 18071
rect 30006 18068 30012 18080
rect 28951 18040 30012 18068
rect 28951 18037 28963 18040
rect 28905 18031 28963 18037
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 30190 18068 30196 18080
rect 30151 18040 30196 18068
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 30392 18077 30420 18108
rect 31938 18096 31944 18108
rect 31996 18096 32002 18148
rect 32950 18096 32956 18148
rect 33008 18136 33014 18148
rect 33244 18136 33272 18235
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 33413 18275 33471 18281
rect 33413 18241 33425 18275
rect 33459 18241 33471 18275
rect 33413 18235 33471 18241
rect 33428 18204 33456 18235
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 34900 18281 34928 18380
rect 35912 18380 37832 18408
rect 34701 18275 34759 18281
rect 34701 18272 34713 18275
rect 34480 18244 34713 18272
rect 34480 18232 34486 18244
rect 34701 18241 34713 18244
rect 34747 18241 34759 18275
rect 34701 18235 34759 18241
rect 34885 18275 34943 18281
rect 34885 18241 34897 18275
rect 34931 18241 34943 18275
rect 34885 18235 34943 18241
rect 33428 18176 34652 18204
rect 33008 18108 33916 18136
rect 33008 18096 33014 18108
rect 33888 18080 33916 18108
rect 30377 18071 30435 18077
rect 30377 18037 30389 18071
rect 30423 18037 30435 18071
rect 30377 18031 30435 18037
rect 31297 18071 31355 18077
rect 31297 18037 31309 18071
rect 31343 18068 31355 18071
rect 31386 18068 31392 18080
rect 31343 18040 31392 18068
rect 31343 18037 31355 18040
rect 31297 18031 31355 18037
rect 31386 18028 31392 18040
rect 31444 18068 31450 18080
rect 32309 18071 32367 18077
rect 32309 18068 32321 18071
rect 31444 18040 32321 18068
rect 31444 18028 31450 18040
rect 32309 18037 32321 18040
rect 32355 18037 32367 18071
rect 32582 18068 32588 18080
rect 32543 18040 32588 18068
rect 32309 18031 32367 18037
rect 32582 18028 32588 18040
rect 32640 18028 32646 18080
rect 33870 18068 33876 18080
rect 33831 18040 33876 18068
rect 33870 18028 33876 18040
rect 33928 18028 33934 18080
rect 34624 18068 34652 18176
rect 34716 18136 34744 18235
rect 34900 18204 34928 18235
rect 35434 18232 35440 18284
rect 35492 18272 35498 18284
rect 35802 18272 35808 18284
rect 35492 18244 35808 18272
rect 35492 18232 35498 18244
rect 35802 18232 35808 18244
rect 35860 18232 35866 18284
rect 35912 18281 35940 18380
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 38378 18408 38384 18420
rect 38304 18380 38384 18408
rect 36906 18340 36912 18352
rect 36004 18312 36912 18340
rect 36004 18281 36032 18312
rect 36906 18300 36912 18312
rect 36964 18300 36970 18352
rect 35897 18275 35955 18281
rect 35897 18241 35909 18275
rect 35943 18241 35955 18275
rect 35897 18235 35955 18241
rect 35989 18275 36047 18281
rect 35989 18241 36001 18275
rect 36035 18241 36047 18275
rect 36170 18272 36176 18284
rect 36131 18244 36176 18272
rect 35989 18235 36047 18241
rect 36170 18232 36176 18244
rect 36228 18232 36234 18284
rect 36265 18275 36323 18281
rect 36265 18241 36277 18275
rect 36311 18272 36323 18275
rect 36538 18272 36544 18284
rect 36311 18244 36544 18272
rect 36311 18241 36323 18244
rect 36265 18235 36323 18241
rect 36538 18232 36544 18244
rect 36596 18232 36602 18284
rect 37366 18232 37372 18284
rect 37424 18272 37430 18284
rect 37826 18272 37832 18284
rect 37424 18244 37832 18272
rect 37424 18232 37430 18244
rect 37826 18232 37832 18244
rect 37884 18232 37890 18284
rect 38304 18281 38332 18380
rect 38378 18368 38384 18380
rect 38436 18368 38442 18420
rect 39298 18368 39304 18420
rect 39356 18408 39362 18420
rect 39669 18411 39727 18417
rect 39669 18408 39681 18411
rect 39356 18380 39681 18408
rect 39356 18368 39362 18380
rect 39669 18377 39681 18380
rect 39715 18377 39727 18411
rect 39669 18371 39727 18377
rect 39758 18368 39764 18420
rect 39816 18408 39822 18420
rect 40402 18408 40408 18420
rect 39816 18380 40408 18408
rect 39816 18368 39822 18380
rect 40402 18368 40408 18380
rect 40460 18368 40466 18420
rect 40586 18368 40592 18420
rect 40644 18408 40650 18420
rect 41049 18411 41107 18417
rect 41049 18408 41061 18411
rect 40644 18380 41061 18408
rect 40644 18368 40650 18380
rect 41049 18377 41061 18380
rect 41095 18377 41107 18411
rect 42794 18408 42800 18420
rect 42755 18380 42800 18408
rect 41049 18371 41107 18377
rect 42794 18368 42800 18380
rect 42852 18368 42858 18420
rect 43530 18368 43536 18420
rect 43588 18408 43594 18420
rect 43809 18411 43867 18417
rect 43809 18408 43821 18411
rect 43588 18380 43821 18408
rect 43588 18368 43594 18380
rect 43809 18377 43821 18380
rect 43855 18377 43867 18411
rect 43809 18371 43867 18377
rect 42978 18300 42984 18352
rect 43036 18340 43042 18352
rect 43349 18343 43407 18349
rect 43349 18340 43361 18343
rect 43036 18312 43361 18340
rect 43036 18300 43042 18312
rect 43349 18309 43361 18312
rect 43395 18340 43407 18343
rect 43438 18340 43444 18352
rect 43395 18312 43444 18340
rect 43395 18309 43407 18312
rect 43349 18303 43407 18309
rect 43438 18300 43444 18312
rect 43496 18340 43502 18352
rect 43496 18312 45416 18340
rect 43496 18300 43502 18312
rect 38289 18275 38347 18281
rect 38289 18241 38301 18275
rect 38335 18241 38347 18275
rect 38289 18235 38347 18241
rect 38378 18232 38384 18284
rect 38436 18272 38442 18284
rect 38473 18275 38531 18281
rect 38473 18272 38485 18275
rect 38436 18244 38485 18272
rect 38436 18232 38442 18244
rect 38473 18241 38485 18244
rect 38519 18241 38531 18275
rect 38473 18235 38531 18241
rect 38654 18232 38660 18284
rect 38712 18272 38718 18284
rect 38749 18275 38807 18281
rect 38749 18272 38761 18275
rect 38712 18244 38761 18272
rect 38712 18232 38718 18244
rect 38749 18241 38761 18244
rect 38795 18241 38807 18275
rect 39482 18272 39488 18284
rect 39443 18244 39488 18272
rect 38749 18235 38807 18241
rect 39482 18232 39488 18244
rect 39540 18232 39546 18284
rect 39574 18232 39580 18284
rect 39632 18272 39638 18284
rect 39853 18275 39911 18281
rect 39853 18272 39865 18275
rect 39632 18244 39865 18272
rect 39632 18232 39638 18244
rect 39853 18241 39865 18244
rect 39899 18241 39911 18275
rect 39853 18235 39911 18241
rect 40865 18275 40923 18281
rect 40865 18241 40877 18275
rect 40911 18272 40923 18275
rect 41322 18272 41328 18284
rect 40911 18244 41328 18272
rect 40911 18241 40923 18244
rect 40865 18235 40923 18241
rect 41322 18232 41328 18244
rect 41380 18232 41386 18284
rect 42797 18275 42855 18281
rect 42797 18241 42809 18275
rect 42843 18272 42855 18275
rect 42886 18272 42892 18284
rect 42843 18244 42892 18272
rect 42843 18241 42855 18244
rect 42797 18235 42855 18241
rect 42886 18232 42892 18244
rect 42944 18232 42950 18284
rect 43254 18232 43260 18284
rect 43312 18272 43318 18284
rect 43806 18272 43812 18284
rect 43312 18244 43812 18272
rect 43312 18232 43318 18244
rect 43806 18232 43812 18244
rect 43864 18232 43870 18284
rect 43993 18275 44051 18281
rect 43993 18241 44005 18275
rect 44039 18272 44051 18275
rect 44266 18272 44272 18284
rect 44039 18244 44272 18272
rect 44039 18241 44051 18244
rect 43993 18235 44051 18241
rect 44266 18232 44272 18244
rect 44324 18232 44330 18284
rect 44910 18232 44916 18284
rect 44968 18272 44974 18284
rect 45388 18281 45416 18312
rect 45097 18275 45155 18281
rect 45097 18272 45109 18275
rect 44968 18244 45109 18272
rect 44968 18232 44974 18244
rect 45097 18241 45109 18244
rect 45143 18241 45155 18275
rect 45097 18235 45155 18241
rect 45373 18275 45431 18281
rect 45373 18241 45385 18275
rect 45419 18241 45431 18275
rect 45373 18235 45431 18241
rect 37734 18204 37740 18216
rect 34900 18176 37740 18204
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 38566 18207 38624 18213
rect 38566 18173 38578 18207
rect 38612 18204 38624 18207
rect 38838 18204 38844 18216
rect 38612 18176 38844 18204
rect 38612 18173 38624 18176
rect 38566 18167 38624 18173
rect 38838 18164 38844 18176
rect 38896 18164 38902 18216
rect 39393 18207 39451 18213
rect 39393 18173 39405 18207
rect 39439 18204 39451 18207
rect 40310 18204 40316 18216
rect 39439 18176 40316 18204
rect 39439 18173 39451 18176
rect 39393 18167 39451 18173
rect 40310 18164 40316 18176
rect 40368 18164 40374 18216
rect 41233 18207 41291 18213
rect 41233 18173 41245 18207
rect 41279 18204 41291 18207
rect 41506 18204 41512 18216
rect 41279 18176 41512 18204
rect 41279 18173 41291 18176
rect 41233 18167 41291 18173
rect 41506 18164 41512 18176
rect 41564 18164 41570 18216
rect 42518 18164 42524 18216
rect 42576 18204 42582 18216
rect 42705 18207 42763 18213
rect 42705 18204 42717 18207
rect 42576 18176 42717 18204
rect 42576 18164 42582 18176
rect 42705 18173 42717 18176
rect 42751 18204 42763 18207
rect 44542 18204 44548 18216
rect 42751 18176 44548 18204
rect 42751 18173 42763 18176
rect 42705 18167 42763 18173
rect 44542 18164 44548 18176
rect 44600 18204 44606 18216
rect 45186 18204 45192 18216
rect 44600 18176 45192 18204
rect 44600 18164 44606 18176
rect 45186 18164 45192 18176
rect 45244 18164 45250 18216
rect 35618 18136 35624 18148
rect 34716 18108 35624 18136
rect 35618 18096 35624 18108
rect 35676 18096 35682 18148
rect 38654 18136 38660 18148
rect 38488 18108 38660 18136
rect 38488 18080 38516 18108
rect 38654 18096 38660 18108
rect 38712 18136 38718 18148
rect 46474 18136 46480 18148
rect 38712 18108 38757 18136
rect 39040 18108 46480 18136
rect 38712 18096 38718 18108
rect 39040 18080 39068 18108
rect 46474 18096 46480 18108
rect 46532 18096 46538 18148
rect 35069 18071 35127 18077
rect 35069 18068 35081 18071
rect 34624 18040 35081 18068
rect 35069 18037 35081 18040
rect 35115 18068 35127 18071
rect 35434 18068 35440 18080
rect 35115 18040 35440 18068
rect 35115 18037 35127 18040
rect 35069 18031 35127 18037
rect 35434 18028 35440 18040
rect 35492 18028 35498 18080
rect 35713 18071 35771 18077
rect 35713 18037 35725 18071
rect 35759 18068 35771 18071
rect 35894 18068 35900 18080
rect 35759 18040 35900 18068
rect 35759 18037 35771 18040
rect 35713 18031 35771 18037
rect 35894 18028 35900 18040
rect 35952 18028 35958 18080
rect 36446 18028 36452 18080
rect 36504 18068 36510 18080
rect 36817 18071 36875 18077
rect 36817 18068 36829 18071
rect 36504 18040 36829 18068
rect 36504 18028 36510 18040
rect 36817 18037 36829 18040
rect 36863 18068 36875 18071
rect 38194 18068 38200 18080
rect 36863 18040 38200 18068
rect 36863 18037 36875 18040
rect 36817 18031 36875 18037
rect 38194 18028 38200 18040
rect 38252 18028 38258 18080
rect 38470 18028 38476 18080
rect 38528 18028 38534 18080
rect 38930 18068 38936 18080
rect 38891 18040 38936 18068
rect 38930 18028 38936 18040
rect 38988 18028 38994 18080
rect 39022 18028 39028 18080
rect 39080 18028 39086 18080
rect 40129 18071 40187 18077
rect 40129 18037 40141 18071
rect 40175 18068 40187 18071
rect 40681 18071 40739 18077
rect 40681 18068 40693 18071
rect 40175 18040 40693 18068
rect 40175 18037 40187 18040
rect 40129 18031 40187 18037
rect 40681 18037 40693 18040
rect 40727 18037 40739 18071
rect 40681 18031 40739 18037
rect 43162 18028 43168 18080
rect 43220 18068 43226 18080
rect 44453 18071 44511 18077
rect 44453 18068 44465 18071
rect 43220 18040 44465 18068
rect 43220 18028 43226 18040
rect 44453 18037 44465 18040
rect 44499 18037 44511 18071
rect 44453 18031 44511 18037
rect 45465 18071 45523 18077
rect 45465 18037 45477 18071
rect 45511 18068 45523 18071
rect 45738 18068 45744 18080
rect 45511 18040 45744 18068
rect 45511 18037 45523 18040
rect 45465 18031 45523 18037
rect 45738 18028 45744 18040
rect 45796 18028 45802 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 24394 17824 24400 17876
rect 24452 17864 24458 17876
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 24452 17836 24685 17864
rect 24452 17824 24458 17836
rect 24673 17833 24685 17836
rect 24719 17833 24731 17867
rect 24673 17827 24731 17833
rect 27157 17867 27215 17873
rect 27157 17833 27169 17867
rect 27203 17864 27215 17867
rect 27522 17864 27528 17876
rect 27203 17836 27528 17864
rect 27203 17833 27215 17836
rect 27157 17827 27215 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 29730 17864 29736 17876
rect 29691 17836 29736 17864
rect 29730 17824 29736 17836
rect 29788 17824 29794 17876
rect 32950 17864 32956 17876
rect 32911 17836 32956 17864
rect 32950 17824 32956 17836
rect 33008 17824 33014 17876
rect 33410 17864 33416 17876
rect 33371 17836 33416 17864
rect 33410 17824 33416 17836
rect 33468 17824 33474 17876
rect 36170 17824 36176 17876
rect 36228 17864 36234 17876
rect 37366 17864 37372 17876
rect 36228 17836 37372 17864
rect 36228 17824 36234 17836
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 38194 17864 38200 17876
rect 38155 17836 38200 17864
rect 38194 17824 38200 17836
rect 38252 17824 38258 17876
rect 38378 17824 38384 17876
rect 38436 17864 38442 17876
rect 40678 17864 40684 17876
rect 38436 17836 40684 17864
rect 38436 17824 38442 17836
rect 40678 17824 40684 17836
rect 40736 17824 40742 17876
rect 41506 17864 41512 17876
rect 41467 17836 41512 17864
rect 41506 17824 41512 17836
rect 41564 17824 41570 17876
rect 42058 17824 42064 17876
rect 42116 17864 42122 17876
rect 42518 17864 42524 17876
rect 42116 17836 42524 17864
rect 42116 17824 42122 17836
rect 42518 17824 42524 17836
rect 42576 17824 42582 17876
rect 43438 17824 43444 17876
rect 43496 17864 43502 17876
rect 43533 17867 43591 17873
rect 43533 17864 43545 17867
rect 43496 17836 43545 17864
rect 43496 17824 43502 17836
rect 43533 17833 43545 17836
rect 43579 17833 43591 17867
rect 43533 17827 43591 17833
rect 25406 17756 25412 17808
rect 25464 17796 25470 17808
rect 25501 17799 25559 17805
rect 25501 17796 25513 17799
rect 25464 17768 25513 17796
rect 25464 17756 25470 17768
rect 25501 17765 25513 17768
rect 25547 17796 25559 17799
rect 27341 17799 27399 17805
rect 25547 17768 26464 17796
rect 25547 17765 25559 17768
rect 25501 17759 25559 17765
rect 24578 17660 24584 17672
rect 24539 17632 24584 17660
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 25038 17660 25044 17672
rect 24811 17632 25044 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 25498 17620 25504 17672
rect 25556 17660 25562 17672
rect 25685 17663 25743 17669
rect 25685 17660 25697 17663
rect 25556 17632 25697 17660
rect 25556 17620 25562 17632
rect 25685 17629 25697 17632
rect 25731 17629 25743 17663
rect 25866 17660 25872 17672
rect 25827 17632 25872 17660
rect 25685 17623 25743 17629
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 25958 17620 25964 17672
rect 26016 17660 26022 17672
rect 26436 17669 26464 17768
rect 27341 17765 27353 17799
rect 27387 17796 27399 17799
rect 28074 17796 28080 17808
rect 27387 17768 28080 17796
rect 27387 17765 27399 17768
rect 27341 17759 27399 17765
rect 28074 17756 28080 17768
rect 28132 17796 28138 17808
rect 30101 17799 30159 17805
rect 28132 17768 28212 17796
rect 28132 17756 28138 17768
rect 26421 17663 26479 17669
rect 26016 17632 26061 17660
rect 26016 17620 26022 17632
rect 26421 17629 26433 17663
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 26510 17620 26516 17672
rect 26568 17660 26574 17672
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 26568 17632 26617 17660
rect 26568 17620 26574 17632
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 26605 17623 26663 17629
rect 27617 17595 27675 17601
rect 27617 17561 27629 17595
rect 27663 17592 27675 17595
rect 27798 17592 27804 17604
rect 27663 17564 27804 17592
rect 27663 17561 27675 17564
rect 27617 17555 27675 17561
rect 27798 17552 27804 17564
rect 27856 17552 27862 17604
rect 26050 17484 26056 17536
rect 26108 17524 26114 17536
rect 28184 17533 28212 17768
rect 30101 17765 30113 17799
rect 30147 17796 30159 17799
rect 30190 17796 30196 17808
rect 30147 17768 30196 17796
rect 30147 17765 30159 17768
rect 30101 17759 30159 17765
rect 30190 17756 30196 17768
rect 30248 17756 30254 17808
rect 31849 17799 31907 17805
rect 31849 17796 31861 17799
rect 30852 17768 31861 17796
rect 30009 17731 30067 17737
rect 30009 17697 30021 17731
rect 30055 17728 30067 17731
rect 30852 17728 30880 17768
rect 31849 17765 31861 17768
rect 31895 17765 31907 17799
rect 31849 17759 31907 17765
rect 35529 17799 35587 17805
rect 35529 17765 35541 17799
rect 35575 17796 35587 17799
rect 36814 17796 36820 17808
rect 35575 17768 36820 17796
rect 35575 17765 35587 17768
rect 35529 17759 35587 17765
rect 36814 17756 36820 17768
rect 36872 17756 36878 17808
rect 38841 17799 38899 17805
rect 38841 17796 38853 17799
rect 37200 17768 38853 17796
rect 30055 17700 30880 17728
rect 30929 17731 30987 17737
rect 30055 17697 30067 17700
rect 30009 17691 30067 17697
rect 30929 17697 30941 17731
rect 30975 17728 30987 17731
rect 30975 17700 31754 17728
rect 30975 17697 30987 17700
rect 30929 17691 30987 17697
rect 29914 17660 29920 17672
rect 29875 17632 29920 17660
rect 29914 17620 29920 17632
rect 29972 17620 29978 17672
rect 30193 17663 30251 17669
rect 30193 17629 30205 17663
rect 30239 17629 30251 17663
rect 31386 17660 31392 17672
rect 31347 17632 31392 17660
rect 30193 17623 30251 17629
rect 28718 17552 28724 17604
rect 28776 17592 28782 17604
rect 29454 17592 29460 17604
rect 28776 17564 29460 17592
rect 28776 17552 28782 17564
rect 29454 17552 29460 17564
rect 29512 17592 29518 17604
rect 30208 17592 30236 17623
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 31726 17660 31754 17700
rect 31938 17688 31944 17740
rect 31996 17728 32002 17740
rect 34057 17731 34115 17737
rect 31996 17700 32076 17728
rect 31996 17688 32002 17700
rect 32048 17669 32076 17700
rect 34057 17697 34069 17731
rect 34103 17728 34115 17731
rect 34698 17728 34704 17740
rect 34103 17700 34704 17728
rect 34103 17697 34115 17700
rect 34057 17691 34115 17697
rect 34698 17688 34704 17700
rect 34756 17688 34762 17740
rect 35434 17728 35440 17740
rect 35395 17700 35440 17728
rect 35434 17688 35440 17700
rect 35492 17688 35498 17740
rect 36262 17728 36268 17740
rect 35535 17700 36268 17728
rect 32033 17663 32091 17669
rect 31726 17632 31984 17660
rect 31846 17592 31852 17604
rect 29512 17564 30236 17592
rect 31807 17564 31852 17592
rect 29512 17552 29518 17564
rect 31846 17552 31852 17564
rect 31904 17552 31910 17604
rect 31956 17592 31984 17632
rect 32033 17629 32045 17663
rect 32079 17629 32091 17663
rect 32033 17623 32091 17629
rect 32122 17620 32128 17672
rect 32180 17660 32186 17672
rect 32180 17632 32225 17660
rect 32180 17620 32186 17632
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 34422 17660 34428 17672
rect 33468 17632 34428 17660
rect 33468 17620 33474 17632
rect 34422 17620 34428 17632
rect 34480 17660 34486 17672
rect 35535 17660 35563 17700
rect 36262 17688 36268 17700
rect 36320 17728 36326 17740
rect 36320 17700 36952 17728
rect 36320 17688 36326 17700
rect 34480 17632 35563 17660
rect 35956 17663 36014 17669
rect 34480 17620 34486 17632
rect 35956 17629 35968 17663
rect 36002 17660 36014 17663
rect 36002 17632 36676 17660
rect 36002 17629 36014 17632
rect 35956 17623 36014 17629
rect 36648 17592 36676 17632
rect 36722 17620 36728 17672
rect 36780 17660 36786 17672
rect 36924 17669 36952 17700
rect 36817 17663 36875 17669
rect 36817 17660 36829 17663
rect 36780 17632 36829 17660
rect 36780 17620 36786 17632
rect 36817 17629 36829 17632
rect 36863 17629 36875 17663
rect 36817 17623 36875 17629
rect 36910 17663 36968 17669
rect 36910 17629 36922 17663
rect 36956 17629 36968 17663
rect 36910 17623 36968 17629
rect 37093 17663 37151 17669
rect 37093 17629 37105 17663
rect 37139 17660 37151 17663
rect 37200 17660 37228 17768
rect 38841 17765 38853 17768
rect 38887 17765 38899 17799
rect 41690 17796 41696 17808
rect 38841 17759 38899 17765
rect 40972 17768 41696 17796
rect 37550 17688 37556 17740
rect 37608 17728 37614 17740
rect 37734 17728 37740 17740
rect 37608 17700 37740 17728
rect 37608 17688 37614 17700
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 37921 17731 37979 17737
rect 37921 17697 37933 17731
rect 37967 17697 37979 17731
rect 37921 17691 37979 17697
rect 37139 17632 37228 17660
rect 37323 17663 37381 17669
rect 37139 17629 37151 17632
rect 37093 17623 37151 17629
rect 37323 17629 37335 17663
rect 37369 17660 37381 17663
rect 37936 17660 37964 17691
rect 38102 17688 38108 17740
rect 38160 17728 38166 17740
rect 40494 17728 40500 17740
rect 38160 17700 40500 17728
rect 38160 17688 38166 17700
rect 40494 17688 40500 17700
rect 40552 17688 40558 17740
rect 40972 17679 41000 17768
rect 41690 17756 41696 17768
rect 41748 17756 41754 17808
rect 42794 17796 42800 17808
rect 42260 17768 42800 17796
rect 41414 17728 41420 17740
rect 41064 17700 41420 17728
rect 40957 17673 41015 17679
rect 37369 17632 37964 17660
rect 38381 17663 38439 17669
rect 37369 17629 37381 17632
rect 37323 17623 37381 17629
rect 38381 17629 38393 17663
rect 38427 17629 38439 17663
rect 38838 17660 38844 17672
rect 38799 17632 38844 17660
rect 38381 17623 38439 17629
rect 37182 17592 37188 17604
rect 31956 17564 36216 17592
rect 36648 17564 37188 17592
rect 26513 17527 26571 17533
rect 26513 17524 26525 17527
rect 26108 17496 26525 17524
rect 26108 17484 26114 17496
rect 26513 17493 26525 17496
rect 26559 17493 26571 17527
rect 26513 17487 26571 17493
rect 28169 17527 28227 17533
rect 28169 17493 28181 17527
rect 28215 17524 28227 17527
rect 28442 17524 28448 17536
rect 28215 17496 28448 17524
rect 28215 17493 28227 17496
rect 28169 17487 28227 17493
rect 28442 17484 28448 17496
rect 28500 17484 28506 17536
rect 31110 17484 31116 17536
rect 31168 17524 31174 17536
rect 31205 17527 31263 17533
rect 31205 17524 31217 17527
rect 31168 17496 31217 17524
rect 31168 17484 31174 17496
rect 31205 17493 31217 17496
rect 31251 17493 31263 17527
rect 31205 17487 31263 17493
rect 31297 17527 31355 17533
rect 31297 17493 31309 17527
rect 31343 17524 31355 17527
rect 31386 17524 31392 17536
rect 31343 17496 31392 17524
rect 31343 17493 31355 17496
rect 31297 17487 31355 17493
rect 31386 17484 31392 17496
rect 31444 17484 31450 17536
rect 33778 17524 33784 17536
rect 33739 17496 33784 17524
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 33873 17527 33931 17533
rect 33873 17493 33885 17527
rect 33919 17524 33931 17527
rect 34054 17524 34060 17536
rect 33919 17496 34060 17524
rect 33919 17493 33931 17496
rect 33873 17487 33931 17493
rect 34054 17484 34060 17496
rect 34112 17484 34118 17536
rect 35894 17524 35900 17536
rect 35855 17496 35900 17524
rect 35894 17484 35900 17496
rect 35952 17484 35958 17536
rect 36078 17524 36084 17536
rect 36039 17496 36084 17524
rect 36078 17484 36084 17496
rect 36136 17484 36142 17536
rect 36188 17524 36216 17564
rect 37182 17552 37188 17564
rect 37240 17552 37246 17604
rect 37642 17552 37648 17604
rect 37700 17592 37706 17604
rect 38396 17592 38424 17623
rect 38838 17620 38844 17632
rect 38896 17620 38902 17672
rect 39114 17660 39120 17672
rect 39027 17632 39120 17660
rect 39114 17620 39120 17632
rect 39172 17660 39178 17672
rect 39942 17660 39948 17672
rect 39172 17632 39948 17660
rect 39172 17620 39178 17632
rect 39942 17620 39948 17632
rect 40000 17620 40006 17672
rect 40126 17660 40132 17672
rect 40087 17632 40132 17660
rect 40126 17620 40132 17632
rect 40184 17620 40190 17672
rect 40405 17663 40463 17669
rect 40405 17629 40417 17663
rect 40451 17629 40463 17663
rect 40957 17639 40969 17673
rect 41003 17639 41015 17673
rect 41064 17669 41092 17700
rect 41414 17688 41420 17700
rect 41472 17688 41478 17740
rect 41506 17688 41512 17740
rect 41564 17728 41570 17740
rect 42260 17737 42288 17768
rect 42794 17756 42800 17768
rect 42852 17756 42858 17808
rect 42886 17756 42892 17808
rect 42944 17796 42950 17808
rect 44177 17799 44235 17805
rect 44177 17796 44189 17799
rect 42944 17768 44189 17796
rect 42944 17756 42950 17768
rect 44177 17765 44189 17768
rect 44223 17765 44235 17799
rect 45189 17799 45247 17805
rect 45189 17796 45201 17799
rect 44177 17759 44235 17765
rect 44468 17768 45201 17796
rect 42245 17731 42303 17737
rect 42245 17728 42257 17731
rect 41564 17700 42257 17728
rect 41564 17688 41570 17700
rect 42245 17697 42257 17700
rect 42291 17697 42303 17731
rect 44468 17728 44496 17768
rect 45189 17765 45201 17768
rect 45235 17765 45247 17799
rect 45189 17759 45247 17765
rect 42245 17691 42303 17697
rect 42352 17700 44496 17728
rect 40957 17633 41015 17639
rect 41049 17663 41107 17669
rect 40405 17623 40463 17629
rect 41049 17629 41061 17663
rect 41095 17629 41107 17663
rect 41230 17660 41236 17672
rect 41191 17632 41236 17660
rect 41049 17623 41107 17629
rect 38470 17592 38476 17604
rect 37700 17564 38476 17592
rect 37700 17552 37706 17564
rect 38470 17552 38476 17564
rect 38528 17552 38534 17604
rect 40218 17592 40224 17604
rect 39224 17564 40224 17592
rect 39224 17536 39252 17564
rect 40218 17552 40224 17564
rect 40276 17552 40282 17604
rect 37461 17527 37519 17533
rect 37461 17524 37473 17527
rect 36188 17496 37473 17524
rect 37461 17493 37473 17496
rect 37507 17493 37519 17527
rect 37461 17487 37519 17493
rect 39025 17527 39083 17533
rect 39025 17493 39037 17527
rect 39071 17524 39083 17527
rect 39206 17524 39212 17536
rect 39071 17496 39212 17524
rect 39071 17493 39083 17496
rect 39025 17487 39083 17493
rect 39206 17484 39212 17496
rect 39264 17484 39270 17536
rect 40310 17524 40316 17536
rect 40271 17496 40316 17524
rect 40310 17484 40316 17496
rect 40368 17484 40374 17536
rect 40420 17524 40448 17623
rect 41215 17620 41236 17632
rect 41288 17620 41294 17672
rect 41322 17663 41380 17669
rect 41322 17629 41334 17663
rect 41368 17660 41380 17663
rect 42352 17660 42380 17700
rect 42426 17660 42432 17672
rect 41368 17654 41460 17660
rect 41524 17654 42380 17660
rect 41368 17632 42380 17654
rect 41368 17629 41380 17632
rect 41322 17623 41380 17629
rect 41432 17626 41552 17632
rect 42418 17620 42432 17660
rect 42484 17620 42490 17672
rect 42702 17620 42708 17672
rect 42760 17660 42766 17672
rect 43162 17660 43168 17672
rect 42760 17632 43168 17660
rect 42760 17620 42766 17632
rect 43162 17620 43168 17632
rect 43220 17620 43226 17672
rect 44468 17669 44496 17700
rect 44910 17688 44916 17740
rect 44968 17728 44974 17740
rect 44968 17700 46060 17728
rect 44968 17688 44974 17700
rect 44453 17663 44511 17669
rect 44453 17629 44465 17663
rect 44499 17629 44511 17663
rect 44453 17623 44511 17629
rect 45094 17620 45100 17672
rect 45152 17660 45158 17672
rect 45189 17663 45247 17669
rect 45189 17660 45201 17663
rect 45152 17632 45201 17660
rect 45152 17620 45158 17632
rect 45189 17629 45201 17632
rect 45235 17629 45247 17663
rect 45189 17623 45247 17629
rect 45373 17663 45431 17669
rect 45373 17629 45385 17663
rect 45419 17660 45431 17663
rect 45462 17660 45468 17672
rect 45419 17632 45468 17660
rect 45419 17629 45431 17632
rect 45373 17623 45431 17629
rect 45462 17620 45468 17632
rect 45520 17620 45526 17672
rect 45830 17660 45836 17672
rect 45791 17632 45836 17660
rect 45830 17620 45836 17632
rect 45888 17620 45894 17672
rect 46032 17669 46060 17700
rect 46017 17663 46075 17669
rect 46017 17629 46029 17663
rect 46063 17629 46075 17663
rect 46017 17623 46075 17629
rect 41215 17592 41243 17620
rect 42418 17601 42446 17620
rect 42383 17595 42446 17601
rect 41215 17564 42288 17592
rect 41966 17524 41972 17536
rect 40420 17496 41972 17524
rect 41966 17484 41972 17496
rect 42024 17484 42030 17536
rect 42260 17524 42288 17564
rect 42383 17561 42395 17595
rect 42429 17564 42446 17595
rect 42518 17592 42524 17604
rect 42479 17564 42524 17592
rect 42429 17561 42441 17564
rect 42383 17555 42441 17561
rect 42518 17552 42524 17564
rect 42576 17552 42582 17604
rect 42610 17552 42616 17604
rect 42668 17592 42674 17604
rect 43530 17601 43536 17604
rect 43517 17595 43536 17601
rect 42668 17564 42761 17592
rect 42668 17552 42674 17564
rect 43517 17561 43529 17595
rect 43517 17555 43536 17561
rect 43530 17552 43536 17555
rect 43588 17552 43594 17604
rect 43717 17595 43775 17601
rect 43717 17561 43729 17595
rect 43763 17592 43775 17595
rect 43990 17592 43996 17604
rect 43763 17564 43996 17592
rect 43763 17561 43775 17564
rect 43717 17555 43775 17561
rect 43990 17552 43996 17564
rect 44048 17552 44054 17604
rect 44174 17592 44180 17604
rect 44135 17564 44180 17592
rect 44174 17552 44180 17564
rect 44232 17552 44238 17604
rect 42628 17524 42656 17552
rect 42260 17496 42656 17524
rect 42794 17484 42800 17536
rect 42852 17524 42858 17536
rect 42889 17527 42947 17533
rect 42889 17524 42901 17527
rect 42852 17496 42901 17524
rect 42852 17484 42858 17496
rect 42889 17493 42901 17496
rect 42935 17493 42947 17527
rect 42889 17487 42947 17493
rect 43254 17484 43260 17536
rect 43312 17524 43318 17536
rect 43349 17527 43407 17533
rect 43349 17524 43361 17527
rect 43312 17496 43361 17524
rect 43312 17484 43318 17496
rect 43349 17493 43361 17496
rect 43395 17493 43407 17527
rect 43349 17487 43407 17493
rect 44361 17527 44419 17533
rect 44361 17493 44373 17527
rect 44407 17524 44419 17527
rect 44542 17524 44548 17536
rect 44407 17496 44548 17524
rect 44407 17493 44419 17496
rect 44361 17487 44419 17493
rect 44542 17484 44548 17496
rect 44600 17524 44606 17536
rect 45833 17527 45891 17533
rect 45833 17524 45845 17527
rect 44600 17496 45845 17524
rect 44600 17484 44606 17496
rect 45833 17493 45845 17496
rect 45879 17493 45891 17527
rect 45833 17487 45891 17493
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 31938 17280 31944 17332
rect 31996 17320 32002 17332
rect 32309 17323 32367 17329
rect 32309 17320 32321 17323
rect 31996 17292 32321 17320
rect 31996 17280 32002 17292
rect 32309 17289 32321 17292
rect 32355 17289 32367 17323
rect 33410 17320 33416 17332
rect 33371 17292 33416 17320
rect 32309 17283 32367 17289
rect 33410 17280 33416 17292
rect 33468 17280 33474 17332
rect 34054 17320 34060 17332
rect 34015 17292 34060 17320
rect 34054 17280 34060 17292
rect 34112 17280 34118 17332
rect 34238 17280 34244 17332
rect 34296 17280 34302 17332
rect 36538 17320 36544 17332
rect 34348 17292 35480 17320
rect 2498 17212 2504 17264
rect 2556 17252 2562 17264
rect 25225 17255 25283 17261
rect 25225 17252 25237 17255
rect 2556 17224 25237 17252
rect 2556 17212 2562 17224
rect 25225 17221 25237 17224
rect 25271 17221 25283 17255
rect 25225 17215 25283 17221
rect 31386 17212 31392 17264
rect 31444 17252 31450 17264
rect 33226 17252 33232 17264
rect 31444 17224 33232 17252
rect 31444 17212 31450 17224
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 1903 17156 2421 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 2409 17153 2421 17156
rect 2455 17184 2467 17187
rect 16850 17184 16856 17196
rect 2455 17156 16856 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 23658 17184 23664 17196
rect 23571 17156 23664 17184
rect 23658 17144 23664 17156
rect 23716 17184 23722 17196
rect 23934 17184 23940 17196
rect 23716 17156 23940 17184
rect 23716 17144 23722 17156
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 24210 17184 24216 17196
rect 24171 17156 24216 17184
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 25038 17144 25044 17196
rect 25096 17184 25102 17196
rect 25593 17187 25651 17193
rect 25593 17184 25605 17187
rect 25096 17156 25605 17184
rect 25096 17144 25102 17156
rect 25593 17153 25605 17156
rect 25639 17153 25651 17187
rect 26050 17184 26056 17196
rect 26011 17156 26056 17184
rect 25593 17147 25651 17153
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 29178 17184 29184 17196
rect 29139 17156 29184 17184
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 30098 17184 30104 17196
rect 30059 17156 30104 17184
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 27614 17116 27620 17128
rect 27575 17088 27620 17116
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 32324 17125 32352 17224
rect 33226 17212 33232 17224
rect 33284 17212 33290 17264
rect 32582 17184 32588 17196
rect 32543 17156 32588 17184
rect 32582 17144 32588 17156
rect 32640 17184 32646 17196
rect 32950 17184 32956 17196
rect 32640 17156 32956 17184
rect 32640 17144 32646 17156
rect 32950 17144 32956 17156
rect 33008 17144 33014 17196
rect 34256 17193 34284 17280
rect 34348 17196 34376 17292
rect 34425 17255 34483 17261
rect 34425 17221 34437 17255
rect 34471 17252 34483 17255
rect 35237 17255 35295 17261
rect 35237 17252 35249 17255
rect 34471 17224 35249 17252
rect 34471 17221 34483 17224
rect 34425 17215 34483 17221
rect 35237 17221 35249 17224
rect 35283 17252 35295 17255
rect 35342 17252 35348 17264
rect 35283 17224 35348 17252
rect 35283 17221 35295 17224
rect 35237 17215 35295 17221
rect 35342 17212 35348 17224
rect 35400 17212 35406 17264
rect 35452 17261 35480 17292
rect 35912 17292 36544 17320
rect 35437 17255 35495 17261
rect 35437 17221 35449 17255
rect 35483 17221 35495 17255
rect 35437 17215 35495 17221
rect 33505 17187 33563 17193
rect 33505 17153 33517 17187
rect 33551 17184 33563 17187
rect 34241 17187 34299 17193
rect 33551 17156 34100 17184
rect 33551 17153 33563 17156
rect 33505 17147 33563 17153
rect 32309 17119 32367 17125
rect 32309 17085 32321 17119
rect 32355 17085 32367 17119
rect 32309 17079 32367 17085
rect 32493 17119 32551 17125
rect 32493 17085 32505 17119
rect 32539 17116 32551 17119
rect 33962 17116 33968 17128
rect 32539 17088 33968 17116
rect 32539 17085 32551 17088
rect 32493 17079 32551 17085
rect 33962 17076 33968 17088
rect 34020 17076 34026 17128
rect 34072 17116 34100 17156
rect 34241 17153 34253 17187
rect 34287 17153 34299 17187
rect 34241 17147 34299 17153
rect 34330 17144 34336 17196
rect 34388 17184 34394 17196
rect 34388 17156 34433 17184
rect 34388 17144 34394 17156
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 35912 17193 35940 17292
rect 36538 17280 36544 17292
rect 36596 17280 36602 17332
rect 36814 17280 36820 17332
rect 36872 17320 36878 17332
rect 37550 17320 37556 17332
rect 36872 17292 37556 17320
rect 36872 17280 36878 17292
rect 37550 17280 37556 17292
rect 37608 17280 37614 17332
rect 37645 17323 37703 17329
rect 37645 17289 37657 17323
rect 37691 17320 37703 17323
rect 37918 17320 37924 17332
rect 37691 17292 37924 17320
rect 37691 17289 37703 17292
rect 37645 17283 37703 17289
rect 37918 17280 37924 17292
rect 37976 17280 37982 17332
rect 38102 17280 38108 17332
rect 38160 17320 38166 17332
rect 39390 17320 39396 17332
rect 38160 17292 39396 17320
rect 38160 17280 38166 17292
rect 39390 17280 39396 17292
rect 39448 17280 39454 17332
rect 39482 17280 39488 17332
rect 39540 17280 39546 17332
rect 40770 17320 40776 17332
rect 40683 17292 40776 17320
rect 40770 17280 40776 17292
rect 40828 17320 40834 17332
rect 41506 17320 41512 17332
rect 40828 17292 41512 17320
rect 40828 17280 40834 17292
rect 41506 17280 41512 17292
rect 41564 17280 41570 17332
rect 42058 17320 42064 17332
rect 42019 17292 42064 17320
rect 42058 17280 42064 17292
rect 42116 17280 42122 17332
rect 39022 17252 39028 17264
rect 36004 17224 39028 17252
rect 34609 17187 34667 17193
rect 34609 17184 34621 17187
rect 34572 17156 34621 17184
rect 34572 17144 34578 17156
rect 34609 17153 34621 17156
rect 34655 17153 34667 17187
rect 34609 17147 34667 17153
rect 35897 17187 35955 17193
rect 35897 17153 35909 17187
rect 35943 17153 35955 17187
rect 35897 17147 35955 17153
rect 34532 17116 34560 17144
rect 34072 17088 34560 17116
rect 1670 17048 1676 17060
rect 1631 17020 1676 17048
rect 1670 17008 1676 17020
rect 1728 17008 1734 17060
rect 27246 17048 27252 17060
rect 27207 17020 27252 17048
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 30653 17051 30711 17057
rect 30653 17017 30665 17051
rect 30699 17048 30711 17051
rect 36004 17048 36032 17224
rect 39022 17212 39028 17224
rect 39080 17212 39086 17264
rect 36081 17187 36139 17193
rect 36081 17153 36093 17187
rect 36127 17184 36139 17187
rect 36541 17187 36599 17193
rect 36541 17184 36553 17187
rect 36127 17156 36553 17184
rect 36127 17153 36139 17156
rect 36081 17147 36139 17153
rect 36541 17153 36553 17156
rect 36587 17153 36599 17187
rect 36541 17147 36599 17153
rect 36556 17116 36584 17147
rect 36630 17144 36636 17196
rect 36688 17184 36694 17196
rect 36725 17187 36783 17193
rect 36725 17184 36737 17187
rect 36688 17156 36737 17184
rect 36688 17144 36694 17156
rect 36725 17153 36737 17156
rect 36771 17153 36783 17187
rect 36725 17147 36783 17153
rect 37461 17187 37519 17193
rect 37461 17153 37473 17187
rect 37507 17184 37519 17187
rect 37550 17184 37556 17196
rect 37507 17156 37556 17184
rect 37507 17153 37519 17156
rect 37461 17147 37519 17153
rect 37550 17144 37556 17156
rect 37608 17144 37614 17196
rect 37734 17184 37740 17196
rect 37695 17156 37740 17184
rect 37734 17144 37740 17156
rect 37792 17184 37798 17196
rect 37792 17156 38516 17184
rect 37792 17144 37798 17156
rect 38378 17116 38384 17128
rect 36556 17088 38384 17116
rect 38378 17076 38384 17088
rect 38436 17076 38442 17128
rect 38488 17116 38516 17156
rect 38654 17144 38660 17196
rect 38712 17184 38718 17196
rect 39209 17187 39267 17193
rect 39209 17184 39221 17187
rect 38712 17156 39221 17184
rect 38712 17144 38718 17156
rect 39209 17153 39221 17156
rect 39255 17184 39267 17187
rect 39298 17184 39304 17196
rect 39255 17156 39304 17184
rect 39255 17153 39267 17156
rect 39209 17147 39267 17153
rect 39298 17144 39304 17156
rect 39356 17144 39362 17196
rect 39393 17187 39451 17193
rect 39393 17153 39405 17187
rect 39439 17184 39451 17187
rect 39500 17184 39528 17280
rect 40494 17212 40500 17264
rect 40552 17252 40558 17264
rect 43257 17255 43315 17261
rect 43257 17252 43269 17255
rect 40552 17224 43269 17252
rect 40552 17212 40558 17224
rect 43257 17221 43269 17224
rect 43303 17221 43315 17255
rect 45002 17252 45008 17264
rect 43257 17215 43315 17221
rect 44314 17224 45008 17252
rect 39439 17156 39528 17184
rect 39439 17153 39451 17156
rect 39393 17147 39451 17153
rect 39574 17144 39580 17196
rect 39632 17184 39638 17196
rect 39853 17187 39911 17193
rect 39853 17184 39865 17187
rect 39632 17156 39865 17184
rect 39632 17144 39638 17156
rect 39853 17153 39865 17156
rect 39899 17153 39911 17187
rect 40678 17184 40684 17196
rect 40639 17156 40684 17184
rect 39853 17147 39911 17153
rect 40678 17144 40684 17156
rect 40736 17144 40742 17196
rect 40954 17184 40960 17196
rect 40915 17156 40960 17184
rect 40954 17144 40960 17156
rect 41012 17144 41018 17196
rect 41322 17144 41328 17196
rect 41380 17184 41386 17196
rect 41417 17187 41475 17193
rect 41417 17184 41429 17187
rect 41380 17156 41429 17184
rect 41380 17144 41386 17156
rect 41417 17153 41429 17156
rect 41463 17153 41475 17187
rect 42610 17184 42616 17196
rect 42571 17156 42616 17184
rect 41417 17147 41475 17153
rect 42610 17144 42616 17156
rect 42668 17144 42674 17196
rect 42794 17184 42800 17196
rect 42755 17156 42800 17184
rect 42794 17144 42800 17156
rect 42852 17144 42858 17196
rect 42886 17144 42892 17196
rect 42944 17184 42950 17196
rect 43070 17193 43076 17196
rect 43027 17187 43076 17193
rect 42944 17156 42989 17184
rect 42944 17144 42950 17156
rect 43027 17153 43039 17187
rect 43073 17153 43076 17187
rect 43027 17147 43076 17153
rect 43070 17144 43076 17147
rect 43128 17144 43134 17196
rect 43530 17144 43536 17196
rect 43588 17184 43594 17196
rect 44314 17193 44342 17224
rect 45002 17212 45008 17224
rect 45060 17252 45066 17264
rect 45060 17224 45416 17252
rect 45060 17212 45066 17224
rect 44299 17187 44357 17193
rect 44299 17184 44311 17187
rect 43588 17156 44311 17184
rect 43588 17144 43594 17156
rect 44299 17153 44311 17156
rect 44345 17153 44357 17187
rect 44299 17147 44357 17153
rect 44453 17187 44511 17193
rect 44453 17153 44465 17187
rect 44499 17184 44511 17187
rect 44910 17184 44916 17196
rect 44499 17156 44916 17184
rect 44499 17153 44511 17156
rect 44453 17147 44511 17153
rect 44910 17144 44916 17156
rect 44968 17144 44974 17196
rect 45388 17193 45416 17224
rect 45373 17187 45431 17193
rect 45373 17153 45385 17187
rect 45419 17153 45431 17187
rect 58069 17187 58127 17193
rect 58069 17184 58081 17187
rect 45373 17147 45431 17153
rect 57440 17156 58081 17184
rect 57440 17128 57468 17156
rect 58069 17153 58081 17156
rect 58115 17153 58127 17187
rect 58069 17147 58127 17153
rect 39114 17116 39120 17128
rect 38488 17088 39120 17116
rect 39114 17076 39120 17088
rect 39172 17076 39178 17128
rect 39945 17119 40003 17125
rect 39945 17116 39957 17119
rect 39316 17088 39957 17116
rect 30699 17020 36032 17048
rect 30699 17017 30711 17020
rect 30653 17011 30711 17017
rect 36630 17008 36636 17060
rect 36688 17048 36694 17060
rect 36906 17048 36912 17060
rect 36688 17020 36912 17048
rect 36688 17008 36694 17020
rect 36906 17008 36912 17020
rect 36964 17008 36970 17060
rect 37182 17008 37188 17060
rect 37240 17048 37246 17060
rect 37461 17051 37519 17057
rect 37461 17048 37473 17051
rect 37240 17020 37473 17048
rect 37240 17008 37246 17020
rect 37461 17017 37473 17020
rect 37507 17017 37519 17051
rect 37461 17011 37519 17017
rect 37642 17008 37648 17060
rect 37700 17008 37706 17060
rect 37918 17008 37924 17060
rect 37976 17048 37982 17060
rect 38562 17048 38568 17060
rect 37976 17020 38568 17048
rect 37976 17008 37982 17020
rect 38562 17008 38568 17020
rect 38620 17048 38626 17060
rect 39316 17048 39344 17088
rect 39945 17085 39957 17088
rect 39991 17085 40003 17119
rect 45005 17119 45063 17125
rect 45005 17116 45017 17119
rect 39945 17079 40003 17085
rect 41432 17088 45017 17116
rect 41432 17060 41460 17088
rect 45005 17085 45017 17088
rect 45051 17085 45063 17119
rect 57422 17116 57428 17128
rect 57383 17088 57428 17116
rect 45005 17079 45063 17085
rect 57422 17076 57428 17088
rect 57480 17076 57486 17128
rect 38620 17020 39344 17048
rect 39393 17051 39451 17057
rect 38620 17008 38626 17020
rect 39393 17017 39405 17051
rect 39439 17048 39451 17051
rect 40126 17048 40132 17060
rect 39439 17020 40132 17048
rect 39439 17017 39451 17020
rect 39393 17011 39451 17017
rect 40126 17008 40132 17020
rect 40184 17008 40190 17060
rect 41414 17008 41420 17060
rect 41472 17008 41478 17060
rect 41966 17008 41972 17060
rect 42024 17048 42030 17060
rect 43530 17048 43536 17060
rect 42024 17020 43536 17048
rect 42024 17008 42030 17020
rect 43530 17008 43536 17020
rect 43588 17008 43594 17060
rect 43990 17008 43996 17060
rect 44048 17048 44054 17060
rect 44085 17051 44143 17057
rect 44085 17048 44097 17051
rect 44048 17020 44097 17048
rect 44048 17008 44054 17020
rect 44085 17017 44097 17020
rect 44131 17017 44143 17051
rect 58250 17048 58256 17060
rect 58211 17020 58256 17048
rect 44085 17011 44143 17017
rect 58250 17008 58256 17020
rect 58308 17008 58314 17060
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 2372 16952 22845 16980
rect 2372 16940 2378 16952
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 25958 16940 25964 16992
rect 26016 16980 26022 16992
rect 27157 16983 27215 16989
rect 27157 16980 27169 16983
rect 26016 16952 27169 16980
rect 26016 16940 26022 16952
rect 27157 16949 27169 16952
rect 27203 16949 27215 16983
rect 27157 16943 27215 16949
rect 33229 16983 33287 16989
rect 33229 16949 33241 16983
rect 33275 16980 33287 16983
rect 33318 16980 33324 16992
rect 33275 16952 33324 16980
rect 33275 16949 33287 16952
rect 33229 16943 33287 16949
rect 33318 16940 33324 16952
rect 33376 16940 33382 16992
rect 33962 16940 33968 16992
rect 34020 16980 34026 16992
rect 35069 16983 35127 16989
rect 35069 16980 35081 16983
rect 34020 16952 35081 16980
rect 34020 16940 34026 16952
rect 35069 16949 35081 16952
rect 35115 16949 35127 16983
rect 35069 16943 35127 16949
rect 35253 16983 35311 16989
rect 35253 16949 35265 16983
rect 35299 16980 35311 16983
rect 35989 16983 36047 16989
rect 35989 16980 36001 16983
rect 35299 16952 36001 16980
rect 35299 16949 35311 16952
rect 35253 16943 35311 16949
rect 35989 16949 36001 16952
rect 36035 16980 36047 16983
rect 36262 16980 36268 16992
rect 36035 16952 36268 16980
rect 36035 16949 36047 16952
rect 35989 16943 36047 16949
rect 36262 16940 36268 16952
rect 36320 16940 36326 16992
rect 36538 16980 36544 16992
rect 36499 16952 36544 16980
rect 36538 16940 36544 16952
rect 36596 16940 36602 16992
rect 36722 16940 36728 16992
rect 36780 16980 36786 16992
rect 37660 16980 37688 17008
rect 36780 16952 37688 16980
rect 36780 16940 36786 16952
rect 37734 16940 37740 16992
rect 37792 16980 37798 16992
rect 38010 16980 38016 16992
rect 37792 16952 38016 16980
rect 37792 16940 37798 16952
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 38102 16940 38108 16992
rect 38160 16980 38166 16992
rect 38473 16983 38531 16989
rect 38473 16980 38485 16983
rect 38160 16952 38485 16980
rect 38160 16940 38166 16952
rect 38473 16949 38485 16952
rect 38519 16949 38531 16983
rect 38473 16943 38531 16949
rect 39945 16983 40003 16989
rect 39945 16949 39957 16983
rect 39991 16980 40003 16983
rect 40034 16980 40040 16992
rect 39991 16952 40040 16980
rect 39991 16949 40003 16952
rect 39945 16943 40003 16949
rect 40034 16940 40040 16952
rect 40092 16940 40098 16992
rect 40221 16983 40279 16989
rect 40221 16949 40233 16983
rect 40267 16980 40279 16983
rect 40402 16980 40408 16992
rect 40267 16952 40408 16980
rect 40267 16949 40279 16952
rect 40221 16943 40279 16949
rect 40402 16940 40408 16952
rect 40460 16940 40466 16992
rect 40954 16980 40960 16992
rect 40915 16952 40960 16980
rect 40954 16940 40960 16952
rect 41012 16940 41018 16992
rect 41322 16940 41328 16992
rect 41380 16980 41386 16992
rect 43162 16980 43168 16992
rect 41380 16952 43168 16980
rect 41380 16940 41386 16952
rect 43162 16940 43168 16952
rect 43220 16980 43226 16992
rect 43898 16980 43904 16992
rect 43220 16952 43904 16980
rect 43220 16940 43226 16952
rect 43898 16940 43904 16952
rect 43956 16940 43962 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 25041 16779 25099 16785
rect 25041 16745 25053 16779
rect 25087 16776 25099 16779
rect 25130 16776 25136 16788
rect 25087 16748 25136 16776
rect 25087 16745 25099 16748
rect 25041 16739 25099 16745
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 25240 16748 27752 16776
rect 24578 16668 24584 16720
rect 24636 16708 24642 16720
rect 25240 16708 25268 16748
rect 24636 16680 25268 16708
rect 24636 16668 24642 16680
rect 25866 16668 25872 16720
rect 25924 16708 25930 16720
rect 27617 16711 27675 16717
rect 27617 16708 27629 16711
rect 25924 16680 27629 16708
rect 25924 16668 25930 16680
rect 27617 16677 27629 16680
rect 27663 16677 27675 16711
rect 27724 16708 27752 16748
rect 28350 16736 28356 16788
rect 28408 16776 28414 16788
rect 28629 16779 28687 16785
rect 28629 16776 28641 16779
rect 28408 16748 28641 16776
rect 28408 16736 28414 16748
rect 28629 16745 28641 16748
rect 28675 16745 28687 16779
rect 28629 16739 28687 16745
rect 28997 16779 29055 16785
rect 28997 16745 29009 16779
rect 29043 16776 29055 16779
rect 29178 16776 29184 16788
rect 29043 16748 29184 16776
rect 29043 16745 29055 16748
rect 28997 16739 29055 16745
rect 29178 16736 29184 16748
rect 29236 16736 29242 16788
rect 33778 16736 33784 16788
rect 33836 16776 33842 16788
rect 33965 16779 34023 16785
rect 33965 16776 33977 16779
rect 33836 16748 33977 16776
rect 33836 16736 33842 16748
rect 33965 16745 33977 16748
rect 34011 16745 34023 16779
rect 33965 16739 34023 16745
rect 34330 16736 34336 16788
rect 34388 16776 34394 16788
rect 37274 16776 37280 16788
rect 34388 16748 37280 16776
rect 34388 16736 34394 16748
rect 37274 16736 37280 16748
rect 37332 16736 37338 16788
rect 37366 16736 37372 16788
rect 37424 16776 37430 16788
rect 38010 16776 38016 16788
rect 37424 16748 38016 16776
rect 37424 16736 37430 16748
rect 38010 16736 38016 16748
rect 38068 16776 38074 16788
rect 38068 16748 38792 16776
rect 38068 16736 38074 16748
rect 31665 16711 31723 16717
rect 31665 16708 31677 16711
rect 27724 16680 31677 16708
rect 27617 16671 27675 16677
rect 31665 16677 31677 16680
rect 31711 16677 31723 16711
rect 33318 16708 33324 16720
rect 31665 16671 31723 16677
rect 32600 16680 33324 16708
rect 26881 16643 26939 16649
rect 26881 16609 26893 16643
rect 26927 16640 26939 16643
rect 27246 16640 27252 16652
rect 26927 16612 27252 16640
rect 26927 16609 26939 16612
rect 26881 16603 26939 16609
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27488 16612 27997 16640
rect 27488 16600 27494 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 25225 16575 25283 16581
rect 25225 16572 25237 16575
rect 25004 16544 25237 16572
rect 25004 16532 25010 16544
rect 25225 16541 25237 16544
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 25332 16448 25360 16535
rect 25406 16532 25412 16584
rect 25464 16572 25470 16584
rect 25501 16575 25559 16581
rect 25501 16572 25513 16575
rect 25464 16544 25513 16572
rect 25464 16532 25470 16544
rect 25501 16541 25513 16544
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 25593 16575 25651 16581
rect 25593 16541 25605 16575
rect 25639 16541 25651 16575
rect 25593 16535 25651 16541
rect 26789 16575 26847 16581
rect 26789 16541 26801 16575
rect 26835 16572 26847 16575
rect 27614 16572 27620 16584
rect 26835 16544 27620 16572
rect 26835 16541 26847 16544
rect 26789 16535 26847 16541
rect 25608 16504 25636 16535
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16572 27859 16575
rect 27890 16572 27896 16584
rect 27847 16544 27896 16572
rect 27847 16541 27859 16544
rect 27801 16535 27859 16541
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 28534 16572 28540 16584
rect 28495 16544 28540 16572
rect 28534 16532 28540 16544
rect 28592 16532 28598 16584
rect 31570 16572 31576 16584
rect 31531 16544 31576 16572
rect 31570 16532 31576 16544
rect 31628 16532 31634 16584
rect 31941 16575 31999 16581
rect 31941 16541 31953 16575
rect 31987 16541 31999 16575
rect 32214 16572 32220 16584
rect 32175 16544 32220 16572
rect 31941 16535 31999 16541
rect 28350 16504 28356 16516
rect 25608 16476 28356 16504
rect 25314 16396 25320 16448
rect 25372 16396 25378 16448
rect 25406 16396 25412 16448
rect 25464 16436 25470 16448
rect 25608 16436 25636 16476
rect 28350 16464 28356 16476
rect 28408 16464 28414 16516
rect 25464 16408 25636 16436
rect 27157 16439 27215 16445
rect 25464 16396 25470 16408
rect 27157 16405 27169 16439
rect 27203 16436 27215 16439
rect 27430 16436 27436 16448
rect 27203 16408 27436 16436
rect 27203 16405 27215 16408
rect 27157 16399 27215 16405
rect 27430 16396 27436 16408
rect 27488 16396 27494 16448
rect 31956 16436 31984 16535
rect 32214 16532 32220 16544
rect 32272 16532 32278 16584
rect 32398 16572 32404 16584
rect 32359 16544 32404 16572
rect 32398 16532 32404 16544
rect 32456 16532 32462 16584
rect 32600 16581 32628 16680
rect 33318 16668 33324 16680
rect 33376 16668 33382 16720
rect 35526 16668 35532 16720
rect 35584 16708 35590 16720
rect 37921 16711 37979 16717
rect 37921 16708 37933 16711
rect 35584 16680 37933 16708
rect 35584 16668 35590 16680
rect 37921 16677 37933 16680
rect 37967 16677 37979 16711
rect 38194 16708 38200 16720
rect 38155 16680 38200 16708
rect 37921 16671 37979 16677
rect 38194 16668 38200 16680
rect 38252 16668 38258 16720
rect 38289 16711 38347 16717
rect 38289 16677 38301 16711
rect 38335 16708 38347 16711
rect 38378 16708 38384 16720
rect 38335 16680 38384 16708
rect 38335 16677 38347 16680
rect 38289 16671 38347 16677
rect 38378 16668 38384 16680
rect 38436 16668 38442 16720
rect 36265 16643 36323 16649
rect 36265 16609 36277 16643
rect 36311 16640 36323 16643
rect 36630 16640 36636 16652
rect 36311 16612 36636 16640
rect 36311 16609 36323 16612
rect 36265 16603 36323 16609
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 37001 16643 37059 16649
rect 37001 16609 37013 16643
rect 37047 16640 37059 16643
rect 37642 16640 37648 16652
rect 37047 16612 37648 16640
rect 37047 16609 37059 16612
rect 37001 16603 37059 16609
rect 37642 16600 37648 16612
rect 37700 16600 37706 16652
rect 38764 16640 38792 16748
rect 38930 16736 38936 16788
rect 38988 16776 38994 16788
rect 39209 16779 39267 16785
rect 39209 16776 39221 16779
rect 38988 16748 39221 16776
rect 38988 16736 38994 16748
rect 39209 16745 39221 16748
rect 39255 16745 39267 16779
rect 39209 16739 39267 16745
rect 39298 16736 39304 16788
rect 39356 16776 39362 16788
rect 41322 16776 41328 16788
rect 39356 16748 41328 16776
rect 39356 16736 39362 16748
rect 41322 16736 41328 16748
rect 41380 16736 41386 16788
rect 42337 16779 42395 16785
rect 42337 16745 42349 16779
rect 42383 16776 42395 16779
rect 43622 16776 43628 16788
rect 42383 16748 43628 16776
rect 42383 16745 42395 16748
rect 42337 16739 42395 16745
rect 43622 16736 43628 16748
rect 43680 16776 43686 16788
rect 44082 16776 44088 16788
rect 43680 16748 44088 16776
rect 43680 16736 43686 16748
rect 44082 16736 44088 16748
rect 44140 16736 44146 16788
rect 38838 16668 38844 16720
rect 38896 16708 38902 16720
rect 41049 16711 41107 16717
rect 41049 16708 41061 16711
rect 38896 16680 41061 16708
rect 38896 16668 38902 16680
rect 41049 16677 41061 16680
rect 41095 16677 41107 16711
rect 41049 16671 41107 16677
rect 39025 16643 39083 16649
rect 39025 16640 39037 16643
rect 38488 16612 38700 16640
rect 38764 16612 39037 16640
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16541 32643 16575
rect 32585 16535 32643 16541
rect 33042 16532 33048 16584
rect 33100 16572 33106 16584
rect 33318 16572 33324 16584
rect 33100 16544 33145 16572
rect 33279 16544 33324 16572
rect 33100 16532 33106 16544
rect 33318 16532 33324 16544
rect 33376 16532 33382 16584
rect 33962 16572 33968 16584
rect 33923 16544 33968 16572
rect 33962 16532 33968 16544
rect 34020 16532 34026 16584
rect 34241 16575 34299 16581
rect 34241 16541 34253 16575
rect 34287 16572 34299 16575
rect 35621 16575 35679 16581
rect 34287 16544 35572 16572
rect 34287 16541 34299 16544
rect 34241 16535 34299 16541
rect 32416 16504 32444 16532
rect 33229 16507 33287 16513
rect 33229 16504 33241 16507
rect 32416 16476 33241 16504
rect 33229 16473 33241 16476
rect 33275 16473 33287 16507
rect 33229 16467 33287 16473
rect 34149 16507 34207 16513
rect 34149 16473 34161 16507
rect 34195 16504 34207 16507
rect 35250 16504 35256 16516
rect 34195 16476 35256 16504
rect 34195 16473 34207 16476
rect 34149 16467 34207 16473
rect 35250 16464 35256 16476
rect 35308 16464 35314 16516
rect 35544 16504 35572 16544
rect 35621 16541 35633 16575
rect 35667 16572 35679 16575
rect 36078 16572 36084 16584
rect 35667 16544 36084 16572
rect 35667 16541 35679 16544
rect 35621 16535 35679 16541
rect 36078 16532 36084 16544
rect 36136 16532 36142 16584
rect 36357 16575 36415 16581
rect 36357 16541 36369 16575
rect 36403 16572 36415 16575
rect 36446 16572 36452 16584
rect 36403 16544 36452 16572
rect 36403 16541 36415 16544
rect 36357 16535 36415 16541
rect 36446 16532 36452 16544
rect 36504 16532 36510 16584
rect 36909 16575 36967 16581
rect 36909 16541 36921 16575
rect 36955 16572 36967 16575
rect 37274 16572 37280 16584
rect 36955 16544 37280 16572
rect 36955 16541 36967 16544
rect 36909 16535 36967 16541
rect 37274 16532 37280 16544
rect 37332 16572 37338 16584
rect 38105 16575 38163 16581
rect 38105 16572 38117 16575
rect 37332 16544 38117 16572
rect 37332 16532 37338 16544
rect 38105 16541 38117 16544
rect 38151 16541 38163 16575
rect 38105 16535 38163 16541
rect 38381 16575 38439 16581
rect 38381 16541 38393 16575
rect 38427 16572 38439 16575
rect 38488 16572 38516 16612
rect 38427 16544 38516 16572
rect 38565 16575 38623 16581
rect 38427 16541 38439 16544
rect 38381 16535 38439 16541
rect 38565 16541 38577 16575
rect 38611 16541 38623 16575
rect 38672 16572 38700 16612
rect 39025 16609 39037 16612
rect 39071 16609 39083 16643
rect 39025 16603 39083 16609
rect 39482 16600 39488 16652
rect 39540 16640 39546 16652
rect 40037 16643 40095 16649
rect 40037 16640 40049 16643
rect 39540 16612 40049 16640
rect 39540 16600 39546 16612
rect 40037 16609 40049 16612
rect 40083 16609 40095 16643
rect 40310 16640 40316 16652
rect 40223 16612 40316 16640
rect 40037 16603 40095 16609
rect 40310 16600 40316 16612
rect 40368 16600 40374 16652
rect 40405 16643 40463 16649
rect 40405 16609 40417 16643
rect 40451 16640 40463 16643
rect 40770 16640 40776 16652
rect 40451 16612 40776 16640
rect 40451 16609 40463 16612
rect 40405 16603 40463 16609
rect 40770 16600 40776 16612
rect 40828 16600 40834 16652
rect 41524 16612 42472 16640
rect 38838 16572 38844 16584
rect 38672 16544 38844 16572
rect 38565 16535 38623 16541
rect 37826 16504 37832 16516
rect 35544 16476 37832 16504
rect 37826 16464 37832 16476
rect 37884 16464 37890 16516
rect 38580 16504 38608 16535
rect 38838 16532 38844 16544
rect 38896 16532 38902 16584
rect 38930 16532 38936 16584
rect 38988 16572 38994 16584
rect 39301 16575 39359 16581
rect 39301 16572 39313 16575
rect 38988 16544 39313 16572
rect 38988 16532 38994 16544
rect 39301 16541 39313 16544
rect 39347 16541 39359 16575
rect 39301 16535 39359 16541
rect 40126 16532 40132 16584
rect 40184 16572 40190 16584
rect 40221 16575 40279 16581
rect 40221 16572 40233 16575
rect 40184 16544 40233 16572
rect 40184 16532 40190 16544
rect 40221 16541 40233 16544
rect 40267 16541 40279 16575
rect 40221 16535 40279 16541
rect 39025 16507 39083 16513
rect 39025 16504 39037 16507
rect 38580 16476 39037 16504
rect 39025 16473 39037 16476
rect 39071 16473 39083 16507
rect 39025 16467 39083 16473
rect 33143 16439 33201 16445
rect 33143 16436 33155 16439
rect 31956 16408 33155 16436
rect 33143 16405 33155 16408
rect 33189 16405 33201 16439
rect 33143 16399 33201 16405
rect 34514 16396 34520 16448
rect 34572 16436 34578 16448
rect 35529 16439 35587 16445
rect 35529 16436 35541 16439
rect 34572 16408 35541 16436
rect 34572 16396 34578 16408
rect 35529 16405 35541 16408
rect 35575 16405 35587 16439
rect 35529 16399 35587 16405
rect 37642 16396 37648 16448
rect 37700 16436 37706 16448
rect 40328 16436 40356 16600
rect 40494 16572 40500 16584
rect 40455 16544 40500 16572
rect 40494 16532 40500 16544
rect 40552 16532 40558 16584
rect 41230 16572 41236 16584
rect 41191 16544 41236 16572
rect 41230 16532 41236 16544
rect 41288 16532 41294 16584
rect 41524 16581 41552 16612
rect 41325 16575 41383 16581
rect 41325 16541 41337 16575
rect 41371 16541 41383 16575
rect 41325 16535 41383 16541
rect 41509 16575 41567 16581
rect 41509 16541 41521 16575
rect 41555 16541 41567 16575
rect 41509 16535 41567 16541
rect 41601 16575 41659 16581
rect 41601 16541 41613 16575
rect 41647 16572 41659 16575
rect 41690 16572 41696 16584
rect 41647 16544 41696 16572
rect 41647 16541 41659 16544
rect 41601 16535 41659 16541
rect 37700 16408 40356 16436
rect 41340 16436 41368 16535
rect 41690 16532 41696 16544
rect 41748 16532 41754 16584
rect 42153 16575 42211 16581
rect 42153 16541 42165 16575
rect 42199 16541 42211 16575
rect 42153 16535 42211 16541
rect 41414 16464 41420 16516
rect 41472 16504 41478 16516
rect 42168 16504 42196 16535
rect 42242 16532 42248 16584
rect 42300 16572 42306 16584
rect 42444 16572 42472 16612
rect 43162 16600 43168 16652
rect 43220 16640 43226 16652
rect 45189 16643 45247 16649
rect 45189 16640 45201 16643
rect 43220 16612 45201 16640
rect 43220 16600 43226 16612
rect 43346 16572 43352 16584
rect 42300 16544 42345 16572
rect 42444 16544 43352 16572
rect 42300 16532 42306 16544
rect 43346 16532 43352 16544
rect 43404 16532 43410 16584
rect 43438 16532 43444 16584
rect 43496 16572 43502 16584
rect 43622 16572 43628 16584
rect 43496 16544 43541 16572
rect 43583 16544 43628 16572
rect 43496 16532 43502 16544
rect 43622 16532 43628 16544
rect 43680 16532 43686 16584
rect 43714 16532 43720 16584
rect 43772 16572 43778 16584
rect 44376 16581 44404 16612
rect 45189 16609 45201 16612
rect 45235 16609 45247 16643
rect 45189 16603 45247 16609
rect 44361 16575 44419 16581
rect 43772 16544 43817 16572
rect 43772 16532 43778 16544
rect 44361 16541 44373 16575
rect 44407 16541 44419 16575
rect 44542 16572 44548 16584
rect 44503 16544 44548 16572
rect 44361 16535 44419 16541
rect 44542 16532 44548 16544
rect 44600 16532 44606 16584
rect 42334 16504 42340 16516
rect 41472 16476 42340 16504
rect 41472 16464 41478 16476
rect 42334 16464 42340 16476
rect 42392 16464 42398 16516
rect 42444 16476 42932 16504
rect 42444 16436 42472 16476
rect 41340 16408 42472 16436
rect 42521 16439 42579 16445
rect 37700 16396 37706 16408
rect 42521 16405 42533 16439
rect 42567 16436 42579 16439
rect 42794 16436 42800 16448
rect 42567 16408 42800 16436
rect 42567 16405 42579 16408
rect 42521 16399 42579 16405
rect 42794 16396 42800 16408
rect 42852 16396 42858 16448
rect 42904 16436 42932 16476
rect 43622 16436 43628 16448
rect 42904 16408 43628 16436
rect 43622 16396 43628 16408
rect 43680 16396 43686 16448
rect 43898 16436 43904 16448
rect 43859 16408 43904 16436
rect 43898 16396 43904 16408
rect 43956 16396 43962 16448
rect 44082 16396 44088 16448
rect 44140 16436 44146 16448
rect 44361 16439 44419 16445
rect 44361 16436 44373 16439
rect 44140 16408 44373 16436
rect 44140 16396 44146 16408
rect 44361 16405 44373 16408
rect 44407 16405 44419 16439
rect 44361 16399 44419 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 24857 16235 24915 16241
rect 24857 16201 24869 16235
rect 24903 16232 24915 16235
rect 25314 16232 25320 16244
rect 24903 16204 25320 16232
rect 24903 16201 24915 16204
rect 24857 16195 24915 16201
rect 25314 16192 25320 16204
rect 25372 16232 25378 16244
rect 28350 16232 28356 16244
rect 25372 16204 26096 16232
rect 28311 16204 28356 16232
rect 25372 16192 25378 16204
rect 25041 16167 25099 16173
rect 25041 16133 25053 16167
rect 25087 16164 25099 16167
rect 25406 16164 25412 16176
rect 25087 16136 25412 16164
rect 25087 16133 25099 16136
rect 25041 16127 25099 16133
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 25777 16167 25835 16173
rect 25777 16133 25789 16167
rect 25823 16164 25835 16167
rect 25958 16164 25964 16176
rect 25823 16136 25964 16164
rect 25823 16133 25835 16136
rect 25777 16127 25835 16133
rect 25958 16124 25964 16136
rect 26016 16124 26022 16176
rect 26068 16164 26096 16204
rect 28350 16192 28356 16204
rect 28408 16192 28414 16244
rect 28534 16192 28540 16244
rect 28592 16192 28598 16244
rect 33321 16235 33379 16241
rect 33321 16201 33333 16235
rect 33367 16232 33379 16235
rect 33594 16232 33600 16244
rect 33367 16204 33600 16232
rect 33367 16201 33379 16204
rect 33321 16195 33379 16201
rect 33594 16192 33600 16204
rect 33652 16192 33658 16244
rect 34606 16232 34612 16244
rect 34567 16204 34612 16232
rect 34606 16192 34612 16204
rect 34664 16192 34670 16244
rect 35342 16192 35348 16244
rect 35400 16232 35406 16244
rect 35437 16235 35495 16241
rect 35437 16232 35449 16235
rect 35400 16204 35449 16232
rect 35400 16192 35406 16204
rect 35437 16201 35449 16204
rect 35483 16201 35495 16235
rect 35437 16195 35495 16201
rect 37826 16192 37832 16244
rect 37884 16232 37890 16244
rect 40494 16232 40500 16244
rect 37884 16204 40500 16232
rect 37884 16192 37890 16204
rect 40494 16192 40500 16204
rect 40552 16232 40558 16244
rect 40770 16232 40776 16244
rect 40552 16204 40776 16232
rect 40552 16192 40558 16204
rect 40770 16192 40776 16204
rect 40828 16192 40834 16244
rect 41506 16232 41512 16244
rect 41467 16204 41512 16232
rect 41506 16192 41512 16204
rect 41564 16192 41570 16244
rect 43622 16192 43628 16244
rect 43680 16232 43686 16244
rect 45462 16232 45468 16244
rect 43680 16204 45468 16232
rect 43680 16192 43686 16204
rect 45462 16192 45468 16204
rect 45520 16192 45526 16244
rect 28552 16164 28580 16192
rect 26068 16136 28580 16164
rect 28626 16124 28632 16176
rect 28684 16164 28690 16176
rect 30098 16164 30104 16176
rect 28684 16136 30104 16164
rect 28684 16124 28690 16136
rect 30098 16124 30104 16136
rect 30156 16124 30162 16176
rect 30561 16167 30619 16173
rect 30561 16133 30573 16167
rect 30607 16164 30619 16167
rect 36449 16167 36507 16173
rect 36449 16164 36461 16167
rect 30607 16136 31340 16164
rect 30607 16133 30619 16136
rect 30561 16127 30619 16133
rect 24765 16099 24823 16105
rect 24765 16065 24777 16099
rect 24811 16065 24823 16099
rect 25498 16096 25504 16108
rect 25459 16068 25504 16096
rect 24765 16059 24823 16065
rect 24780 16028 24808 16059
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16096 25651 16099
rect 25866 16096 25872 16108
rect 25639 16068 25872 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 25866 16056 25872 16068
rect 25924 16056 25930 16108
rect 27430 16096 27436 16108
rect 27391 16068 27436 16096
rect 27430 16056 27436 16068
rect 27488 16056 27494 16108
rect 28537 16099 28595 16105
rect 28537 16096 28549 16099
rect 27816 16068 28549 16096
rect 24946 16028 24952 16040
rect 24780 16000 24952 16028
rect 24946 15988 24952 16000
rect 25004 16028 25010 16040
rect 27816 16037 27844 16068
rect 28537 16065 28549 16068
rect 28583 16096 28595 16099
rect 29086 16096 29092 16108
rect 28583 16068 29092 16096
rect 28583 16065 28595 16068
rect 28537 16059 28595 16065
rect 29086 16056 29092 16068
rect 29144 16056 29150 16108
rect 29454 16096 29460 16108
rect 29415 16068 29460 16096
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 29914 16056 29920 16108
rect 29972 16096 29978 16108
rect 30374 16096 30380 16108
rect 29972 16068 30380 16096
rect 29972 16056 29978 16068
rect 30374 16056 30380 16068
rect 30432 16056 30438 16108
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16096 30711 16099
rect 31110 16096 31116 16108
rect 30699 16068 31116 16096
rect 30699 16065 30711 16068
rect 30653 16059 30711 16065
rect 31110 16056 31116 16068
rect 31168 16056 31174 16108
rect 31312 16105 31340 16136
rect 35544 16136 36461 16164
rect 31297 16099 31355 16105
rect 31297 16065 31309 16099
rect 31343 16096 31355 16099
rect 31386 16096 31392 16108
rect 31343 16068 31392 16096
rect 31343 16065 31355 16068
rect 31297 16059 31355 16065
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 32490 16096 32496 16108
rect 32451 16068 32496 16096
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16096 32735 16099
rect 33134 16096 33140 16108
rect 32723 16068 33140 16096
rect 32723 16065 32735 16068
rect 32677 16059 32735 16065
rect 33134 16056 33140 16068
rect 33192 16056 33198 16108
rect 33318 16099 33376 16105
rect 33318 16065 33330 16099
rect 33364 16065 33376 16099
rect 33318 16059 33376 16065
rect 27525 16031 27583 16037
rect 25004 16000 26648 16028
rect 25004 15988 25010 16000
rect 25038 15960 25044 15972
rect 24999 15932 25044 15960
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 25685 15895 25743 15901
rect 25685 15861 25697 15895
rect 25731 15892 25743 15895
rect 26510 15892 26516 15904
rect 25731 15864 26516 15892
rect 25731 15861 25743 15864
rect 25685 15855 25743 15861
rect 26510 15852 26516 15864
rect 26568 15852 26574 15904
rect 26620 15892 26648 16000
rect 27525 15997 27537 16031
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 27801 16031 27859 16037
rect 27801 15997 27813 16031
rect 27847 15997 27859 16031
rect 28810 16028 28816 16040
rect 28771 16000 28816 16028
rect 27801 15991 27859 15997
rect 27540 15960 27568 15991
rect 28810 15988 28816 16000
rect 28868 15988 28874 16040
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 31205 16031 31263 16037
rect 31205 16028 31217 16031
rect 29779 16000 31217 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 31205 15997 31217 16000
rect 31251 15997 31263 16031
rect 31205 15991 31263 15997
rect 27890 15960 27896 15972
rect 27540 15932 27896 15960
rect 27890 15920 27896 15932
rect 27948 15960 27954 15972
rect 29273 15963 29331 15969
rect 29273 15960 29285 15963
rect 27948 15932 29285 15960
rect 27948 15920 27954 15932
rect 29273 15929 29285 15932
rect 29319 15929 29331 15963
rect 29273 15923 29331 15929
rect 29362 15920 29368 15972
rect 29420 15960 29426 15972
rect 33137 15963 33195 15969
rect 33137 15960 33149 15963
rect 29420 15932 33149 15960
rect 29420 15920 29426 15932
rect 33137 15929 33149 15932
rect 33183 15929 33195 15963
rect 33333 15960 33361 16059
rect 33686 16056 33692 16108
rect 33744 16096 33750 16108
rect 33781 16099 33839 16105
rect 33781 16096 33793 16099
rect 33744 16068 33793 16096
rect 33744 16056 33750 16068
rect 33781 16065 33793 16068
rect 33827 16065 33839 16099
rect 33781 16059 33839 16065
rect 34885 16099 34943 16105
rect 34885 16065 34897 16099
rect 34931 16065 34943 16099
rect 34885 16059 34943 16065
rect 34422 15988 34428 16040
rect 34480 16028 34486 16040
rect 34609 16031 34667 16037
rect 34609 16028 34621 16031
rect 34480 16000 34621 16028
rect 34480 15988 34486 16000
rect 34609 15997 34621 16000
rect 34655 15997 34667 16031
rect 34900 16028 34928 16059
rect 35434 16056 35440 16108
rect 35492 16096 35498 16108
rect 35544 16105 35572 16136
rect 36449 16133 36461 16136
rect 36495 16164 36507 16167
rect 36538 16164 36544 16176
rect 36495 16136 36544 16164
rect 36495 16133 36507 16136
rect 36449 16127 36507 16133
rect 36538 16124 36544 16136
rect 36596 16124 36602 16176
rect 40310 16124 40316 16176
rect 40368 16164 40374 16176
rect 40862 16164 40868 16176
rect 40368 16136 40868 16164
rect 40368 16124 40374 16136
rect 40862 16124 40868 16136
rect 40920 16164 40926 16176
rect 43806 16164 43812 16176
rect 40920 16136 41552 16164
rect 40920 16124 40926 16136
rect 35529 16099 35587 16105
rect 35529 16096 35541 16099
rect 35492 16068 35541 16096
rect 35492 16056 35498 16068
rect 35529 16065 35541 16068
rect 35575 16065 35587 16099
rect 35529 16059 35587 16065
rect 36725 16099 36783 16105
rect 36725 16065 36737 16099
rect 36771 16096 36783 16099
rect 36998 16096 37004 16108
rect 36771 16068 37004 16096
rect 36771 16065 36783 16068
rect 36725 16059 36783 16065
rect 36998 16056 37004 16068
rect 37056 16056 37062 16108
rect 37550 16056 37556 16108
rect 37608 16096 37614 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 37608 16068 37657 16096
rect 37608 16056 37614 16068
rect 37645 16065 37657 16068
rect 37691 16065 37703 16099
rect 37918 16096 37924 16108
rect 37879 16068 37924 16096
rect 37645 16059 37703 16065
rect 37918 16056 37924 16068
rect 37976 16056 37982 16108
rect 39298 16096 39304 16108
rect 39259 16068 39304 16096
rect 39298 16056 39304 16068
rect 39356 16056 39362 16108
rect 39482 16096 39488 16108
rect 39443 16068 39488 16096
rect 39482 16056 39488 16068
rect 39540 16056 39546 16108
rect 39761 16099 39819 16105
rect 39761 16065 39773 16099
rect 39807 16096 39819 16099
rect 40221 16099 40279 16105
rect 40221 16096 40233 16099
rect 39807 16068 40233 16096
rect 39807 16065 39819 16068
rect 39761 16059 39819 16065
rect 40221 16065 40233 16068
rect 40267 16065 40279 16099
rect 40402 16096 40408 16108
rect 40363 16068 40408 16096
rect 40221 16059 40279 16065
rect 40402 16056 40408 16068
rect 40460 16056 40466 16108
rect 41325 16099 41383 16105
rect 41325 16065 41337 16099
rect 41371 16096 41383 16099
rect 41414 16096 41420 16108
rect 41371 16068 41420 16096
rect 41371 16065 41383 16068
rect 41325 16059 41383 16065
rect 41414 16056 41420 16068
rect 41472 16056 41478 16108
rect 41524 16105 41552 16136
rect 41800 16136 43812 16164
rect 41509 16099 41567 16105
rect 41509 16065 41521 16099
rect 41555 16065 41567 16099
rect 41509 16059 41567 16065
rect 35802 16028 35808 16040
rect 34900 16000 35808 16028
rect 34609 15991 34667 15997
rect 35802 15988 35808 16000
rect 35860 15988 35866 16040
rect 36538 16028 36544 16040
rect 36499 16000 36544 16028
rect 36538 15988 36544 16000
rect 36596 15988 36602 16040
rect 39574 16028 39580 16040
rect 39535 16000 39580 16028
rect 39574 15988 39580 16000
rect 39632 15988 39638 16040
rect 40681 16031 40739 16037
rect 40681 15997 40693 16031
rect 40727 16028 40739 16031
rect 40862 16028 40868 16040
rect 40727 16000 40868 16028
rect 40727 15997 40739 16000
rect 40681 15991 40739 15997
rect 40862 15988 40868 16000
rect 40920 16028 40926 16040
rect 41800 16028 41828 16136
rect 43806 16124 43812 16136
rect 43864 16164 43870 16176
rect 44177 16167 44235 16173
rect 43864 16136 44036 16164
rect 43864 16124 43870 16136
rect 41874 16056 41880 16108
rect 41932 16096 41938 16108
rect 43438 16096 43444 16108
rect 41932 16068 43444 16096
rect 41932 16056 41938 16068
rect 43438 16056 43444 16068
rect 43496 16056 43502 16108
rect 43714 16056 43720 16108
rect 43772 16096 43778 16108
rect 43901 16099 43959 16105
rect 43901 16096 43913 16099
rect 43772 16068 43913 16096
rect 43772 16056 43778 16068
rect 43901 16065 43913 16068
rect 43947 16065 43959 16099
rect 44008 16096 44036 16136
rect 44177 16133 44189 16167
rect 44223 16164 44235 16167
rect 44266 16164 44272 16176
rect 44223 16136 44272 16164
rect 44223 16133 44235 16136
rect 44177 16127 44235 16133
rect 44266 16124 44272 16136
rect 44324 16124 44330 16176
rect 44913 16099 44971 16105
rect 44913 16096 44925 16099
rect 44008 16068 44925 16096
rect 43901 16059 43959 16065
rect 44913 16065 44925 16068
rect 44959 16065 44971 16099
rect 45186 16096 45192 16108
rect 45147 16068 45192 16096
rect 44913 16059 44971 16065
rect 45186 16056 45192 16068
rect 45244 16056 45250 16108
rect 40920 16000 41828 16028
rect 40920 15988 40926 16000
rect 43070 15988 43076 16040
rect 43128 16028 43134 16040
rect 43809 16031 43867 16037
rect 43809 16028 43821 16031
rect 43128 16000 43821 16028
rect 43128 15988 43134 16000
rect 43809 15997 43821 16000
rect 43855 15997 43867 16031
rect 43809 15991 43867 15997
rect 44269 16031 44327 16037
rect 44269 15997 44281 16031
rect 44315 16028 44327 16031
rect 44450 16028 44456 16040
rect 44315 16000 44456 16028
rect 44315 15997 44327 16000
rect 44269 15991 44327 15997
rect 33333 15932 35572 15960
rect 33137 15923 33195 15929
rect 28626 15892 28632 15904
rect 26620 15864 28632 15892
rect 28626 15852 28632 15864
rect 28684 15852 28690 15904
rect 28721 15895 28779 15901
rect 28721 15861 28733 15895
rect 28767 15892 28779 15895
rect 29178 15892 29184 15904
rect 28767 15864 29184 15892
rect 28767 15861 28779 15864
rect 28721 15855 28779 15861
rect 29178 15852 29184 15864
rect 29236 15852 29242 15904
rect 29641 15895 29699 15901
rect 29641 15861 29653 15895
rect 29687 15892 29699 15895
rect 30193 15895 30251 15901
rect 30193 15892 30205 15895
rect 29687 15864 30205 15892
rect 29687 15861 29699 15864
rect 29641 15855 29699 15861
rect 30193 15861 30205 15864
rect 30239 15861 30251 15895
rect 30193 15855 30251 15861
rect 31938 15852 31944 15904
rect 31996 15892 32002 15904
rect 32309 15895 32367 15901
rect 32309 15892 32321 15895
rect 31996 15864 32321 15892
rect 31996 15852 32002 15864
rect 32309 15861 32321 15864
rect 32355 15861 32367 15895
rect 32582 15892 32588 15904
rect 32543 15864 32588 15892
rect 32309 15855 32367 15861
rect 32582 15852 32588 15864
rect 32640 15852 32646 15904
rect 33689 15895 33747 15901
rect 33689 15861 33701 15895
rect 33735 15892 33747 15895
rect 33870 15892 33876 15904
rect 33735 15864 33876 15892
rect 33735 15861 33747 15864
rect 33689 15855 33747 15861
rect 33870 15852 33876 15864
rect 33928 15892 33934 15904
rect 34330 15892 34336 15904
rect 33928 15864 34336 15892
rect 33928 15852 33934 15864
rect 34330 15852 34336 15864
rect 34388 15852 34394 15904
rect 34790 15852 34796 15904
rect 34848 15892 34854 15904
rect 35544 15892 35572 15932
rect 36170 15920 36176 15972
rect 36228 15960 36234 15972
rect 37829 15963 37887 15969
rect 37829 15960 37841 15963
rect 36228 15932 37841 15960
rect 36228 15920 36234 15932
rect 37829 15929 37841 15932
rect 37875 15960 37887 15963
rect 39393 15963 39451 15969
rect 37875 15932 39344 15960
rect 37875 15929 37887 15932
rect 37829 15923 37887 15929
rect 35618 15892 35624 15904
rect 34848 15864 34893 15892
rect 35544 15864 35624 15892
rect 34848 15852 34854 15864
rect 35618 15852 35624 15864
rect 35676 15852 35682 15904
rect 36722 15892 36728 15904
rect 36683 15864 36728 15892
rect 36722 15852 36728 15864
rect 36780 15852 36786 15904
rect 36906 15892 36912 15904
rect 36867 15864 36912 15892
rect 36906 15852 36912 15864
rect 36964 15852 36970 15904
rect 37366 15852 37372 15904
rect 37424 15892 37430 15904
rect 37461 15895 37519 15901
rect 37461 15892 37473 15895
rect 37424 15864 37473 15892
rect 37424 15852 37430 15864
rect 37461 15861 37473 15864
rect 37507 15861 37519 15895
rect 37461 15855 37519 15861
rect 37918 15852 37924 15904
rect 37976 15892 37982 15904
rect 38102 15892 38108 15904
rect 37976 15864 38108 15892
rect 37976 15852 37982 15864
rect 38102 15852 38108 15864
rect 38160 15852 38166 15904
rect 39114 15892 39120 15904
rect 39075 15864 39120 15892
rect 39114 15852 39120 15864
rect 39172 15852 39178 15904
rect 39316 15892 39344 15932
rect 39393 15929 39405 15963
rect 39439 15960 39451 15963
rect 40954 15960 40960 15972
rect 39439 15932 40960 15960
rect 39439 15929 39451 15932
rect 39393 15923 39451 15929
rect 40954 15920 40960 15932
rect 41012 15920 41018 15972
rect 43824 15960 43852 15991
rect 44450 15988 44456 16000
rect 44508 16028 44514 16040
rect 44729 16031 44787 16037
rect 44729 16028 44741 16031
rect 44508 16000 44741 16028
rect 44508 15988 44514 16000
rect 44729 15997 44741 16000
rect 44775 15997 44787 16031
rect 44729 15991 44787 15997
rect 43824 15932 45692 15960
rect 45664 15904 45692 15932
rect 39758 15892 39764 15904
rect 39316 15864 39764 15892
rect 39758 15852 39764 15864
rect 39816 15852 39822 15904
rect 40589 15895 40647 15901
rect 40589 15861 40601 15895
rect 40635 15892 40647 15895
rect 40770 15892 40776 15904
rect 40635 15864 40776 15892
rect 40635 15861 40647 15864
rect 40589 15855 40647 15861
rect 40770 15852 40776 15864
rect 40828 15852 40834 15904
rect 43622 15892 43628 15904
rect 43583 15864 43628 15892
rect 43622 15852 43628 15864
rect 43680 15852 43686 15904
rect 45094 15892 45100 15904
rect 45055 15864 45100 15892
rect 45094 15852 45100 15864
rect 45152 15852 45158 15904
rect 45646 15892 45652 15904
rect 45607 15864 45652 15892
rect 45646 15852 45652 15864
rect 45704 15852 45710 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 28721 15691 28779 15697
rect 28721 15688 28733 15691
rect 28592 15660 28733 15688
rect 28592 15648 28598 15660
rect 28721 15657 28733 15660
rect 28767 15657 28779 15691
rect 28721 15651 28779 15657
rect 29089 15691 29147 15697
rect 29089 15657 29101 15691
rect 29135 15688 29147 15691
rect 29270 15688 29276 15700
rect 29135 15660 29276 15688
rect 29135 15657 29147 15660
rect 29089 15651 29147 15657
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 31570 15688 31576 15700
rect 31531 15660 31576 15688
rect 31570 15648 31576 15660
rect 31628 15688 31634 15700
rect 33226 15688 33232 15700
rect 31628 15660 33232 15688
rect 31628 15648 31634 15660
rect 33226 15648 33232 15660
rect 33284 15648 33290 15700
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 34885 15691 34943 15697
rect 34885 15688 34897 15691
rect 34848 15660 34897 15688
rect 34848 15648 34854 15660
rect 34885 15657 34897 15660
rect 34931 15657 34943 15691
rect 34885 15651 34943 15657
rect 35069 15691 35127 15697
rect 35069 15657 35081 15691
rect 35115 15688 35127 15691
rect 35342 15688 35348 15700
rect 35115 15660 35348 15688
rect 35115 15657 35127 15660
rect 35069 15651 35127 15657
rect 35342 15648 35348 15660
rect 35400 15648 35406 15700
rect 40218 15688 40224 15700
rect 40179 15660 40224 15688
rect 40218 15648 40224 15660
rect 40276 15648 40282 15700
rect 41138 15688 41144 15700
rect 41051 15660 41144 15688
rect 41138 15648 41144 15660
rect 41196 15688 41202 15700
rect 42058 15688 42064 15700
rect 41196 15660 42064 15688
rect 41196 15648 41202 15660
rect 42058 15648 42064 15660
rect 42116 15648 42122 15700
rect 25682 15580 25688 15632
rect 25740 15620 25746 15632
rect 31389 15623 31447 15629
rect 31389 15620 31401 15623
rect 25740 15592 31401 15620
rect 25740 15580 25746 15592
rect 31389 15589 31401 15592
rect 31435 15589 31447 15623
rect 31389 15583 31447 15589
rect 34054 15580 34060 15632
rect 34112 15620 34118 15632
rect 36446 15620 36452 15632
rect 34112 15592 36452 15620
rect 34112 15580 34118 15592
rect 36446 15580 36452 15592
rect 36504 15620 36510 15632
rect 36541 15623 36599 15629
rect 36541 15620 36553 15623
rect 36504 15592 36553 15620
rect 36504 15580 36510 15592
rect 36541 15589 36553 15592
rect 36587 15589 36599 15623
rect 36541 15583 36599 15589
rect 36906 15580 36912 15632
rect 36964 15620 36970 15632
rect 42610 15620 42616 15632
rect 36964 15592 42616 15620
rect 36964 15580 36970 15592
rect 42610 15580 42616 15592
rect 42668 15580 42674 15632
rect 26878 15512 26884 15564
rect 26936 15552 26942 15564
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 26936 15524 26985 15552
rect 26936 15512 26942 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 29362 15552 29368 15564
rect 26973 15515 27031 15521
rect 27264 15524 29368 15552
rect 27264 15496 27292 15524
rect 29362 15512 29368 15524
rect 29420 15512 29426 15564
rect 30650 15512 30656 15564
rect 30708 15552 30714 15564
rect 31665 15555 31723 15561
rect 30708 15524 31432 15552
rect 30708 15512 30714 15524
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 24302 15484 24308 15496
rect 23615 15456 24308 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 23400 15416 23428 15447
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 25590 15484 25596 15496
rect 25551 15456 25596 15484
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 26099 15456 26188 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 26160 15428 26188 15456
rect 26418 15444 26424 15496
rect 26476 15484 26482 15496
rect 27157 15487 27215 15493
rect 27157 15484 27169 15487
rect 26476 15456 27169 15484
rect 26476 15444 26482 15456
rect 27157 15453 27169 15456
rect 27203 15453 27215 15487
rect 27157 15447 27215 15453
rect 27246 15444 27252 15496
rect 27304 15484 27310 15496
rect 27304 15456 27397 15484
rect 27304 15444 27310 15456
rect 28810 15444 28816 15496
rect 28868 15484 28874 15496
rect 28905 15487 28963 15493
rect 28905 15484 28917 15487
rect 28868 15456 28917 15484
rect 28868 15444 28874 15456
rect 28905 15453 28917 15456
rect 28951 15453 28963 15487
rect 28905 15447 28963 15453
rect 29086 15444 29092 15496
rect 29144 15484 29150 15496
rect 31404 15484 31432 15524
rect 31665 15521 31677 15555
rect 31711 15552 31723 15555
rect 32401 15555 32459 15561
rect 32401 15552 32413 15555
rect 31711 15524 32413 15552
rect 31711 15521 31723 15524
rect 31665 15515 31723 15521
rect 32401 15521 32413 15524
rect 32447 15521 32459 15555
rect 32401 15515 32459 15521
rect 32490 15512 32496 15564
rect 32548 15552 32554 15564
rect 32769 15555 32827 15561
rect 32548 15524 32720 15552
rect 32548 15512 32554 15524
rect 31938 15484 31944 15496
rect 29144 15456 29189 15484
rect 31404 15456 31754 15484
rect 31899 15456 31944 15484
rect 29144 15444 29150 15456
rect 23934 15416 23940 15428
rect 23400 15388 23940 15416
rect 23934 15376 23940 15388
rect 23992 15416 23998 15428
rect 23992 15388 24978 15416
rect 23992 15376 23998 15388
rect 26142 15376 26148 15428
rect 26200 15376 26206 15428
rect 26878 15376 26884 15428
rect 26936 15416 26942 15428
rect 27801 15419 27859 15425
rect 27801 15416 27813 15419
rect 26936 15388 27813 15416
rect 26936 15376 26942 15388
rect 27801 15385 27813 15388
rect 27847 15416 27859 15419
rect 29638 15416 29644 15428
rect 27847 15388 29644 15416
rect 27847 15385 27859 15388
rect 27801 15379 27859 15385
rect 29638 15376 29644 15388
rect 29696 15376 29702 15428
rect 30469 15419 30527 15425
rect 30469 15385 30481 15419
rect 30515 15385 30527 15419
rect 30650 15416 30656 15428
rect 30611 15388 30656 15416
rect 30469 15379 30527 15385
rect 23474 15348 23480 15360
rect 23435 15320 23480 15348
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 26970 15348 26976 15360
rect 26931 15320 26976 15348
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 30285 15351 30343 15357
rect 30285 15348 30297 15351
rect 29052 15320 30297 15348
rect 29052 15308 29058 15320
rect 30285 15317 30297 15320
rect 30331 15317 30343 15351
rect 30484 15348 30512 15379
rect 30650 15376 30656 15388
rect 30708 15376 30714 15428
rect 31726 15416 31754 15456
rect 31938 15444 31944 15456
rect 31996 15444 32002 15496
rect 32582 15484 32588 15496
rect 32543 15456 32588 15484
rect 32582 15444 32588 15456
rect 32640 15444 32646 15496
rect 32692 15484 32720 15524
rect 32769 15521 32781 15555
rect 32815 15552 32827 15555
rect 33134 15552 33140 15564
rect 32815 15524 33140 15552
rect 32815 15521 32827 15524
rect 32769 15515 32827 15521
rect 33134 15512 33140 15524
rect 33192 15552 33198 15564
rect 33686 15552 33692 15564
rect 33192 15524 33692 15552
rect 33192 15512 33198 15524
rect 33686 15512 33692 15524
rect 33744 15512 33750 15564
rect 35618 15512 35624 15564
rect 35676 15552 35682 15564
rect 37461 15555 37519 15561
rect 35676 15524 37044 15552
rect 35676 15512 35682 15524
rect 32861 15487 32919 15493
rect 32861 15484 32873 15487
rect 32692 15456 32873 15484
rect 32861 15453 32873 15456
rect 32907 15453 32919 15487
rect 32861 15447 32919 15453
rect 33318 15444 33324 15496
rect 33376 15484 33382 15496
rect 33781 15487 33839 15493
rect 33781 15484 33793 15487
rect 33376 15456 33793 15484
rect 33376 15444 33382 15456
rect 33781 15453 33793 15456
rect 33827 15453 33839 15487
rect 33962 15484 33968 15496
rect 33923 15456 33968 15484
rect 33781 15447 33839 15453
rect 33962 15444 33968 15456
rect 34020 15444 34026 15496
rect 34057 15487 34115 15493
rect 34057 15453 34069 15487
rect 34103 15453 34115 15487
rect 35986 15484 35992 15496
rect 34057 15447 34115 15453
rect 35820 15456 35992 15484
rect 33597 15419 33655 15425
rect 33597 15416 33609 15419
rect 31726 15388 33609 15416
rect 33597 15385 33609 15388
rect 33643 15385 33655 15419
rect 33597 15379 33655 15385
rect 31018 15348 31024 15360
rect 30484 15320 31024 15348
rect 30285 15311 30343 15317
rect 31018 15308 31024 15320
rect 31076 15348 31082 15360
rect 33042 15348 33048 15360
rect 31076 15320 33048 15348
rect 31076 15308 31082 15320
rect 33042 15308 33048 15320
rect 33100 15308 33106 15360
rect 34072 15348 34100 15447
rect 34698 15376 34704 15428
rect 34756 15416 34762 15428
rect 35253 15419 35311 15425
rect 35253 15416 35265 15419
rect 34756 15388 35265 15416
rect 34756 15376 34762 15388
rect 35253 15385 35265 15388
rect 35299 15416 35311 15419
rect 35820 15416 35848 15456
rect 35986 15444 35992 15456
rect 36044 15444 36050 15496
rect 36354 15444 36360 15496
rect 36412 15484 36418 15496
rect 36449 15487 36507 15493
rect 36449 15484 36461 15487
rect 36412 15456 36461 15484
rect 36412 15444 36418 15456
rect 36449 15453 36461 15456
rect 36495 15453 36507 15487
rect 36449 15447 36507 15453
rect 36725 15487 36783 15493
rect 36725 15453 36737 15487
rect 36771 15484 36783 15487
rect 36906 15484 36912 15496
rect 36771 15456 36912 15484
rect 36771 15453 36783 15456
rect 36725 15447 36783 15453
rect 36906 15444 36912 15456
rect 36964 15444 36970 15496
rect 37016 15484 37044 15524
rect 37461 15521 37473 15555
rect 37507 15552 37519 15555
rect 38381 15555 38439 15561
rect 38381 15552 38393 15555
rect 37507 15524 38393 15552
rect 37507 15521 37519 15524
rect 37461 15515 37519 15521
rect 38381 15521 38393 15524
rect 38427 15552 38439 15555
rect 40126 15552 40132 15564
rect 38427 15524 40132 15552
rect 38427 15521 38439 15524
rect 38381 15515 38439 15521
rect 40126 15512 40132 15524
rect 40184 15512 40190 15564
rect 40310 15552 40316 15564
rect 40271 15524 40316 15552
rect 40310 15512 40316 15524
rect 40368 15512 40374 15564
rect 42794 15512 42800 15564
rect 42852 15552 42858 15564
rect 43073 15555 43131 15561
rect 43073 15552 43085 15555
rect 42852 15524 43085 15552
rect 42852 15512 42858 15524
rect 43073 15521 43085 15524
rect 43119 15521 43131 15555
rect 43898 15552 43904 15564
rect 43859 15524 43904 15552
rect 43073 15515 43131 15521
rect 43898 15512 43904 15524
rect 43956 15512 43962 15564
rect 45094 15512 45100 15564
rect 45152 15552 45158 15564
rect 46293 15555 46351 15561
rect 46293 15552 46305 15555
rect 45152 15524 45600 15552
rect 45152 15512 45158 15524
rect 37274 15484 37280 15496
rect 37016 15456 37280 15484
rect 37274 15444 37280 15456
rect 37332 15484 37338 15496
rect 37553 15487 37611 15493
rect 37553 15484 37565 15487
rect 37332 15456 37565 15484
rect 37332 15444 37338 15456
rect 37553 15453 37565 15456
rect 37599 15453 37611 15487
rect 37553 15447 37611 15453
rect 37645 15487 37703 15493
rect 37645 15453 37657 15487
rect 37691 15453 37703 15487
rect 37645 15447 37703 15453
rect 37737 15487 37795 15493
rect 37737 15453 37749 15487
rect 37783 15484 37795 15487
rect 38286 15484 38292 15496
rect 37783 15456 38292 15484
rect 37783 15453 37795 15456
rect 37737 15447 37795 15453
rect 35299 15388 35848 15416
rect 35299 15385 35311 15388
rect 35253 15379 35311 15385
rect 35894 15376 35900 15428
rect 35952 15416 35958 15428
rect 37660 15416 37688 15447
rect 38286 15444 38292 15456
rect 38344 15444 38350 15496
rect 40589 15487 40647 15493
rect 40589 15453 40601 15487
rect 40635 15484 40647 15487
rect 41138 15484 41144 15496
rect 40635 15456 41144 15484
rect 40635 15453 40647 15456
rect 40589 15447 40647 15453
rect 41138 15444 41144 15456
rect 41196 15444 41202 15496
rect 42518 15484 42524 15496
rect 42479 15456 42524 15484
rect 42518 15444 42524 15456
rect 42576 15444 42582 15496
rect 43257 15487 43315 15493
rect 43257 15453 43269 15487
rect 43303 15453 43315 15487
rect 43806 15484 43812 15496
rect 43767 15456 43812 15484
rect 43257 15447 43315 15453
rect 35952 15388 37688 15416
rect 35952 15376 35958 15388
rect 35053 15351 35111 15357
rect 35053 15348 35065 15351
rect 34072 15320 35065 15348
rect 35053 15317 35065 15320
rect 35099 15348 35111 15351
rect 36170 15348 36176 15360
rect 35099 15320 36176 15348
rect 35099 15317 35111 15320
rect 35053 15311 35111 15317
rect 36170 15308 36176 15320
rect 36228 15308 36234 15360
rect 36354 15308 36360 15360
rect 36412 15348 36418 15360
rect 37277 15351 37335 15357
rect 37277 15348 37289 15351
rect 36412 15320 37289 15348
rect 36412 15308 36418 15320
rect 37277 15317 37289 15320
rect 37323 15317 37335 15351
rect 37660 15348 37688 15388
rect 38102 15376 38108 15428
rect 38160 15416 38166 15428
rect 42613 15419 42671 15425
rect 42613 15416 42625 15419
rect 38160 15388 42625 15416
rect 38160 15376 38166 15388
rect 42613 15385 42625 15388
rect 42659 15385 42671 15419
rect 43272 15416 43300 15447
rect 43806 15444 43812 15456
rect 43864 15444 43870 15496
rect 45462 15484 45468 15496
rect 45423 15456 45468 15484
rect 45462 15444 45468 15456
rect 45520 15444 45526 15496
rect 45572 15493 45600 15524
rect 45664 15524 46305 15552
rect 45664 15496 45692 15524
rect 46293 15521 46305 15524
rect 46339 15521 46351 15555
rect 46293 15515 46351 15521
rect 45557 15487 45615 15493
rect 45557 15453 45569 15487
rect 45603 15453 45615 15487
rect 45557 15447 45615 15453
rect 45646 15444 45652 15496
rect 45704 15484 45710 15496
rect 45704 15456 45749 15484
rect 45704 15444 45710 15456
rect 45830 15444 45836 15496
rect 45888 15484 45894 15496
rect 45888 15456 45933 15484
rect 45888 15444 45894 15456
rect 45189 15419 45247 15425
rect 45189 15416 45201 15419
rect 43272 15388 45201 15416
rect 42613 15379 42671 15385
rect 45189 15385 45201 15388
rect 45235 15385 45247 15419
rect 45189 15379 45247 15385
rect 38838 15348 38844 15360
rect 37660 15320 38844 15348
rect 37277 15311 37335 15317
rect 38838 15308 38844 15320
rect 38896 15308 38902 15360
rect 40034 15348 40040 15360
rect 39995 15320 40040 15348
rect 40034 15308 40040 15320
rect 40092 15308 40098 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 25590 15104 25596 15156
rect 25648 15144 25654 15156
rect 26053 15147 26111 15153
rect 26053 15144 26065 15147
rect 25648 15116 26065 15144
rect 25648 15104 25654 15116
rect 26053 15113 26065 15116
rect 26099 15113 26111 15147
rect 29178 15144 29184 15156
rect 26053 15107 26111 15113
rect 28184 15116 29184 15144
rect 27246 15076 27252 15088
rect 26068 15048 27252 15076
rect 23934 15008 23940 15020
rect 23895 14980 23940 15008
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 24302 15008 24308 15020
rect 24263 14980 24308 15008
rect 24302 14968 24308 14980
rect 24360 14968 24366 15020
rect 26068 15017 26096 15048
rect 27246 15036 27252 15048
rect 27304 15036 27310 15088
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26970 15008 26976 15020
rect 26467 14980 26976 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 27525 15011 27583 15017
rect 27525 14977 27537 15011
rect 27571 15008 27583 15011
rect 27982 15008 27988 15020
rect 27571 14980 27988 15008
rect 27571 14977 27583 14980
rect 27525 14971 27583 14977
rect 25869 14943 25927 14949
rect 25869 14909 25881 14943
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 24210 14872 24216 14884
rect 24171 14844 24216 14872
rect 24210 14832 24216 14844
rect 24268 14832 24274 14884
rect 25884 14872 25912 14903
rect 26142 14900 26148 14952
rect 26200 14940 26206 14952
rect 27154 14940 27160 14952
rect 26200 14912 27160 14940
rect 26200 14900 26206 14912
rect 27154 14900 27160 14912
rect 27212 14900 27218 14952
rect 27356 14940 27384 14971
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28184 15017 28212 15116
rect 29178 15104 29184 15116
rect 29236 15144 29242 15156
rect 30282 15144 30288 15156
rect 29236 15116 30288 15144
rect 29236 15104 29242 15116
rect 30282 15104 30288 15116
rect 30340 15144 30346 15156
rect 31294 15144 31300 15156
rect 30340 15116 31300 15144
rect 30340 15104 30346 15116
rect 31294 15104 31300 15116
rect 31352 15104 31358 15156
rect 31665 15147 31723 15153
rect 31665 15113 31677 15147
rect 31711 15144 31723 15147
rect 32582 15144 32588 15156
rect 31711 15116 32588 15144
rect 31711 15113 31723 15116
rect 31665 15107 31723 15113
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 33042 15144 33048 15156
rect 33003 15116 33048 15144
rect 33042 15104 33048 15116
rect 33100 15104 33106 15156
rect 33686 15144 33692 15156
rect 33647 15116 33692 15144
rect 33686 15104 33692 15116
rect 33744 15104 33750 15156
rect 35250 15104 35256 15156
rect 35308 15144 35314 15156
rect 36170 15144 36176 15156
rect 35308 15116 36176 15144
rect 35308 15104 35314 15116
rect 36170 15104 36176 15116
rect 36228 15104 36234 15156
rect 36354 15144 36360 15156
rect 36280 15116 36360 15144
rect 28994 15076 29000 15088
rect 28552 15048 29000 15076
rect 28552 15017 28580 15048
rect 28994 15036 29000 15048
rect 29052 15036 29058 15088
rect 30558 15076 30564 15088
rect 29840 15048 30564 15076
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28537 15011 28595 15017
rect 28537 14977 28549 15011
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28813 15011 28871 15017
rect 28813 14977 28825 15011
rect 28859 14977 28871 15011
rect 28813 14971 28871 14977
rect 27798 14940 27804 14952
rect 27356 14912 27804 14940
rect 27798 14900 27804 14912
rect 27856 14940 27862 14952
rect 28353 14943 28411 14949
rect 28353 14940 28365 14943
rect 27856 14912 28365 14940
rect 27856 14900 27862 14912
rect 28353 14909 28365 14912
rect 28399 14909 28411 14943
rect 28353 14903 28411 14909
rect 26418 14872 26424 14884
rect 25884 14844 26424 14872
rect 26418 14832 26424 14844
rect 26476 14832 26482 14884
rect 28166 14832 28172 14884
rect 28224 14872 28230 14884
rect 28828 14872 28856 14971
rect 28902 14968 28908 15020
rect 28960 15008 28966 15020
rect 29840 15017 29868 15048
rect 30558 15036 30564 15048
rect 30616 15036 30622 15088
rect 31772 15048 32720 15076
rect 29825 15011 29883 15017
rect 28960 14980 29005 15008
rect 28960 14968 28966 14980
rect 29825 14977 29837 15011
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 30285 15011 30343 15017
rect 30285 14977 30297 15011
rect 30331 14977 30343 15011
rect 30285 14971 30343 14977
rect 30469 15011 30527 15017
rect 30469 14977 30481 15011
rect 30515 15008 30527 15011
rect 30650 15008 30656 15020
rect 30515 14980 30656 15008
rect 30515 14977 30527 14980
rect 30469 14971 30527 14977
rect 30300 14940 30328 14971
rect 30650 14968 30656 14980
rect 30708 14968 30714 15020
rect 31772 15017 31800 15048
rect 32692 15020 32720 15048
rect 32766 15036 32772 15088
rect 32824 15076 32830 15088
rect 36280 15076 36308 15116
rect 36354 15104 36360 15116
rect 36412 15104 36418 15156
rect 36446 15104 36452 15156
rect 36504 15104 36510 15156
rect 36725 15147 36783 15153
rect 36725 15113 36737 15147
rect 36771 15144 36783 15147
rect 42426 15144 42432 15156
rect 36771 15116 42432 15144
rect 36771 15113 36783 15116
rect 36725 15107 36783 15113
rect 42426 15104 42432 15116
rect 42484 15104 42490 15156
rect 44082 15144 44088 15156
rect 44043 15116 44088 15144
rect 44082 15104 44088 15116
rect 44140 15104 44146 15156
rect 36464 15076 36492 15104
rect 32824 15048 36308 15076
rect 36372 15048 36492 15076
rect 32824 15036 32830 15048
rect 31757 15011 31815 15017
rect 31757 14977 31769 15011
rect 31803 14977 31815 15011
rect 31757 14971 31815 14977
rect 32549 15011 32607 15017
rect 32549 14977 32561 15011
rect 32595 14977 32607 15011
rect 32674 15008 32680 15020
rect 32635 14980 32680 15008
rect 32549 14971 32607 14977
rect 32214 14940 32220 14952
rect 30300 14912 32220 14940
rect 32214 14900 32220 14912
rect 32272 14940 32278 14952
rect 32564 14940 32592 14971
rect 32674 14968 32680 14980
rect 32732 14968 32738 15020
rect 32861 15011 32919 15017
rect 32861 14977 32873 15011
rect 32907 15008 32919 15011
rect 33042 15008 33048 15020
rect 32907 14980 33048 15008
rect 32907 14977 32919 14980
rect 32861 14971 32919 14977
rect 33042 14968 33048 14980
rect 33100 15008 33106 15020
rect 33796 15017 33824 15048
rect 33597 15011 33655 15017
rect 33597 15008 33609 15011
rect 33100 14980 33609 15008
rect 33100 14968 33106 14980
rect 33597 14977 33609 14980
rect 33643 14977 33655 15011
rect 33597 14971 33655 14977
rect 33781 15011 33839 15017
rect 33781 14977 33793 15011
rect 33827 14977 33839 15011
rect 33781 14971 33839 14977
rect 34698 14968 34704 15020
rect 34756 15008 34762 15020
rect 35069 15011 35127 15017
rect 35069 15008 35081 15011
rect 34756 14980 35081 15008
rect 34756 14968 34762 14980
rect 35069 14977 35081 14980
rect 35115 14977 35127 15011
rect 35250 15008 35256 15020
rect 35211 14980 35256 15008
rect 35069 14971 35127 14977
rect 35250 14968 35256 14980
rect 35308 14968 35314 15020
rect 35434 15008 35440 15020
rect 35395 14980 35440 15008
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 35618 15008 35624 15020
rect 35579 14980 35624 15008
rect 35618 14968 35624 14980
rect 35676 14968 35682 15020
rect 35894 14968 35900 15020
rect 35952 15008 35958 15020
rect 36078 15008 36084 15020
rect 35952 14980 36084 15008
rect 35952 14968 35958 14980
rect 36078 14968 36084 14980
rect 36136 14968 36142 15020
rect 36262 15008 36268 15020
rect 36223 14980 36268 15008
rect 36262 14968 36268 14980
rect 36320 14968 36326 15020
rect 36372 15017 36400 15048
rect 36906 15036 36912 15088
rect 36964 15076 36970 15088
rect 37553 15079 37611 15085
rect 37553 15076 37565 15079
rect 36964 15048 37565 15076
rect 36964 15036 36970 15048
rect 37553 15045 37565 15048
rect 37599 15076 37611 15079
rect 38105 15079 38163 15085
rect 38105 15076 38117 15079
rect 37599 15048 38117 15076
rect 37599 15045 37611 15048
rect 37553 15039 37611 15045
rect 38105 15045 38117 15048
rect 38151 15076 38163 15079
rect 38562 15076 38568 15088
rect 38151 15048 38568 15076
rect 38151 15045 38163 15048
rect 38105 15039 38163 15045
rect 38562 15036 38568 15048
rect 38620 15036 38626 15088
rect 40957 15079 41015 15085
rect 38948 15048 40908 15076
rect 36357 15011 36415 15017
rect 36357 14977 36369 15011
rect 36403 14977 36415 15011
rect 36357 14971 36415 14977
rect 36449 15011 36507 15017
rect 36449 14977 36461 15011
rect 36495 15008 36507 15011
rect 37734 15008 37740 15020
rect 36495 14980 37740 15008
rect 36495 14977 36507 14980
rect 36449 14971 36507 14977
rect 37734 14968 37740 14980
rect 37792 14968 37798 15020
rect 38470 14968 38476 15020
rect 38528 15008 38534 15020
rect 38948 15017 38976 15048
rect 38841 15011 38899 15017
rect 38841 15008 38853 15011
rect 38528 14980 38853 15008
rect 38528 14968 38534 14980
rect 38841 14977 38853 14980
rect 38887 14977 38899 15011
rect 38841 14971 38899 14977
rect 38933 15011 38991 15017
rect 38933 14977 38945 15011
rect 38979 14977 38991 15011
rect 38933 14971 38991 14977
rect 33134 14940 33140 14952
rect 32272 14912 33140 14940
rect 32272 14900 32278 14912
rect 33134 14900 33140 14912
rect 33192 14900 33198 14952
rect 35342 14940 35348 14952
rect 35303 14912 35348 14940
rect 35342 14900 35348 14912
rect 35400 14900 35406 14952
rect 38856 14940 38884 14971
rect 39022 14968 39028 15020
rect 39080 15008 39086 15020
rect 39209 15011 39267 15017
rect 39080 14980 39125 15008
rect 39080 14968 39086 14980
rect 39209 14977 39221 15011
rect 39255 15008 39267 15011
rect 39298 15008 39304 15020
rect 39255 14980 39304 15008
rect 39255 14977 39267 14980
rect 39209 14971 39267 14977
rect 39298 14968 39304 14980
rect 39356 14968 39362 15020
rect 39574 14968 39580 15020
rect 39632 15008 39638 15020
rect 39761 15011 39819 15017
rect 39761 15008 39773 15011
rect 39632 14980 39773 15008
rect 39632 14968 39638 14980
rect 39761 14977 39773 14980
rect 39807 14977 39819 15011
rect 40034 15008 40040 15020
rect 39995 14980 40040 15008
rect 39761 14971 39819 14977
rect 40034 14968 40040 14980
rect 40092 14968 40098 15020
rect 40678 15008 40684 15020
rect 40639 14980 40684 15008
rect 40678 14968 40684 14980
rect 40736 14968 40742 15020
rect 40773 15011 40831 15017
rect 40773 14977 40785 15011
rect 40819 14977 40831 15011
rect 40773 14971 40831 14977
rect 39666 14940 39672 14952
rect 38856 14912 39672 14940
rect 39666 14900 39672 14912
rect 39724 14940 39730 14952
rect 39853 14943 39911 14949
rect 39853 14940 39865 14943
rect 39724 14912 39865 14940
rect 39724 14900 39730 14912
rect 39853 14909 39865 14912
rect 39899 14909 39911 14943
rect 39853 14903 39911 14909
rect 39945 14943 40003 14949
rect 39945 14909 39957 14943
rect 39991 14940 40003 14943
rect 40218 14940 40224 14952
rect 39991 14912 40224 14940
rect 39991 14909 40003 14912
rect 39945 14903 40003 14909
rect 40218 14900 40224 14912
rect 40276 14900 40282 14952
rect 40402 14900 40408 14952
rect 40460 14940 40466 14952
rect 40788 14940 40816 14971
rect 40460 14912 40816 14940
rect 40460 14900 40466 14912
rect 32766 14881 32772 14884
rect 30377 14875 30435 14881
rect 30377 14872 30389 14875
rect 28224 14844 30389 14872
rect 28224 14832 28230 14844
rect 30377 14841 30389 14844
rect 30423 14841 30435 14875
rect 32765 14872 32772 14881
rect 32727 14844 32772 14872
rect 30377 14835 30435 14841
rect 32765 14835 32772 14844
rect 32766 14832 32772 14835
rect 32824 14832 32830 14884
rect 32950 14832 32956 14884
rect 33008 14872 33014 14884
rect 36078 14872 36084 14884
rect 33008 14844 36084 14872
rect 33008 14832 33014 14844
rect 36078 14832 36084 14844
rect 36136 14872 36142 14884
rect 37366 14872 37372 14884
rect 36136 14844 37372 14872
rect 36136 14832 36142 14844
rect 37366 14832 37372 14844
rect 37424 14872 37430 14884
rect 38562 14872 38568 14884
rect 37424 14844 38424 14872
rect 38523 14844 38568 14872
rect 37424 14832 37430 14844
rect 29638 14804 29644 14816
rect 29599 14776 29644 14804
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 34330 14804 34336 14816
rect 34291 14776 34336 14804
rect 34330 14764 34336 14776
rect 34388 14764 34394 14816
rect 34885 14807 34943 14813
rect 34885 14773 34897 14807
rect 34931 14804 34943 14807
rect 35342 14804 35348 14816
rect 34931 14776 35348 14804
rect 34931 14773 34943 14776
rect 34885 14767 34943 14773
rect 35342 14764 35348 14776
rect 35400 14764 35406 14816
rect 38396 14804 38424 14844
rect 38562 14832 38568 14844
rect 38620 14832 38626 14884
rect 40880 14872 40908 15048
rect 40957 15045 40969 15079
rect 41003 15076 41015 15079
rect 41506 15076 41512 15088
rect 41003 15048 41512 15076
rect 41003 15045 41015 15048
rect 40957 15039 41015 15045
rect 41506 15036 41512 15048
rect 41564 15036 41570 15088
rect 42061 15079 42119 15085
rect 42061 15045 42073 15079
rect 42107 15076 42119 15079
rect 42107 15048 43208 15076
rect 42107 15045 42119 15048
rect 42061 15039 42119 15045
rect 41598 15008 41604 15020
rect 41511 14980 41604 15008
rect 41598 14968 41604 14980
rect 41656 14968 41662 15020
rect 41782 15008 41788 15020
rect 41743 14980 41788 15008
rect 41782 14968 41788 14980
rect 41840 14968 41846 15020
rect 41877 15011 41935 15017
rect 41877 14977 41889 15011
rect 41923 15008 41935 15011
rect 42150 15008 42156 15020
rect 41923 14980 42156 15008
rect 41923 14977 41935 14980
rect 41877 14971 41935 14977
rect 42150 14968 42156 14980
rect 42208 14968 42214 15020
rect 42702 15008 42708 15020
rect 42663 14980 42708 15008
rect 42702 14968 42708 14980
rect 42760 14968 42766 15020
rect 42794 14968 42800 15020
rect 42852 15008 42858 15020
rect 43180 15017 43208 15048
rect 42981 15011 43039 15017
rect 42981 15008 42993 15011
rect 42852 14980 42993 15008
rect 42852 14968 42858 14980
rect 42981 14977 42993 14980
rect 43027 14977 43039 15011
rect 42981 14971 43039 14977
rect 43165 15011 43223 15017
rect 43165 14977 43177 15011
rect 43211 14977 43223 15011
rect 44450 15008 44456 15020
rect 44411 14980 44456 15008
rect 43165 14971 43223 14977
rect 44450 14968 44456 14980
rect 44508 14968 44514 15020
rect 41616 14872 41644 14968
rect 41966 14940 41972 14952
rect 41879 14912 41972 14940
rect 41966 14900 41972 14912
rect 42024 14940 42030 14952
rect 42886 14940 42892 14952
rect 42024 14912 42892 14940
rect 42024 14900 42030 14912
rect 42886 14900 42892 14912
rect 42944 14900 42950 14952
rect 43441 14943 43499 14949
rect 43441 14909 43453 14943
rect 43487 14909 43499 14943
rect 43441 14903 43499 14909
rect 42702 14872 42708 14884
rect 40880 14844 41552 14872
rect 41616 14844 42708 14872
rect 38930 14804 38936 14816
rect 38396 14776 38936 14804
rect 38930 14764 38936 14776
rect 38988 14764 38994 14816
rect 39298 14764 39304 14816
rect 39356 14804 39362 14816
rect 40221 14807 40279 14813
rect 40221 14804 40233 14807
rect 39356 14776 40233 14804
rect 39356 14764 39362 14776
rect 40221 14773 40233 14776
rect 40267 14773 40279 14807
rect 40221 14767 40279 14773
rect 40957 14807 41015 14813
rect 40957 14773 40969 14807
rect 41003 14804 41015 14807
rect 41046 14804 41052 14816
rect 41003 14776 41052 14804
rect 41003 14773 41015 14776
rect 40957 14767 41015 14773
rect 41046 14764 41052 14776
rect 41104 14764 41110 14816
rect 41524 14804 41552 14844
rect 42702 14832 42708 14844
rect 42760 14832 42766 14884
rect 43346 14872 43352 14884
rect 43307 14844 43352 14872
rect 43346 14832 43352 14844
rect 43404 14832 43410 14884
rect 43456 14872 43484 14903
rect 43901 14875 43959 14881
rect 43901 14872 43913 14875
rect 43456 14844 43913 14872
rect 43901 14841 43913 14844
rect 43947 14841 43959 14875
rect 43901 14835 43959 14841
rect 41690 14804 41696 14816
rect 41524 14776 41696 14804
rect 41690 14764 41696 14776
rect 41748 14804 41754 14816
rect 42150 14804 42156 14816
rect 41748 14776 42156 14804
rect 41748 14764 41754 14776
rect 42150 14764 42156 14776
rect 42208 14764 42214 14816
rect 43806 14764 43812 14816
rect 43864 14804 43870 14816
rect 44085 14807 44143 14813
rect 44085 14804 44097 14807
rect 43864 14776 44097 14804
rect 43864 14764 43870 14776
rect 44085 14773 44097 14776
rect 44131 14773 44143 14807
rect 44085 14767 44143 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 25317 14603 25375 14609
rect 25317 14569 25329 14603
rect 25363 14600 25375 14603
rect 26142 14600 26148 14612
rect 25363 14572 26148 14600
rect 25363 14569 25375 14572
rect 25317 14563 25375 14569
rect 26142 14560 26148 14572
rect 26200 14560 26206 14612
rect 26421 14603 26479 14609
rect 26421 14569 26433 14603
rect 26467 14600 26479 14603
rect 26878 14600 26884 14612
rect 26467 14572 26884 14600
rect 26467 14569 26479 14572
rect 26421 14563 26479 14569
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 26973 14603 27031 14609
rect 26973 14569 26985 14603
rect 27019 14600 27031 14603
rect 27522 14600 27528 14612
rect 27019 14572 27528 14600
rect 27019 14569 27031 14572
rect 26973 14563 27031 14569
rect 27522 14560 27528 14572
rect 27580 14600 27586 14612
rect 27706 14600 27712 14612
rect 27580 14572 27712 14600
rect 27580 14560 27586 14572
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 27982 14600 27988 14612
rect 27943 14572 27988 14600
rect 27982 14560 27988 14572
rect 28040 14560 28046 14612
rect 29178 14600 29184 14612
rect 29139 14572 29184 14600
rect 29178 14560 29184 14572
rect 29236 14560 29242 14612
rect 30006 14560 30012 14612
rect 30064 14600 30070 14612
rect 30193 14603 30251 14609
rect 30193 14600 30205 14603
rect 30064 14572 30205 14600
rect 30064 14560 30070 14572
rect 30193 14569 30205 14572
rect 30239 14569 30251 14603
rect 31386 14600 31392 14612
rect 31347 14572 31392 14600
rect 30193 14563 30251 14569
rect 31386 14560 31392 14572
rect 31444 14560 31450 14612
rect 33962 14560 33968 14612
rect 34020 14600 34026 14612
rect 34241 14603 34299 14609
rect 34241 14600 34253 14603
rect 34020 14572 34253 14600
rect 34020 14560 34026 14572
rect 34241 14569 34253 14572
rect 34287 14600 34299 14603
rect 36538 14600 36544 14612
rect 34287 14572 36544 14600
rect 34287 14569 34299 14572
rect 34241 14563 34299 14569
rect 36538 14560 36544 14572
rect 36596 14600 36602 14612
rect 36909 14603 36967 14609
rect 36909 14600 36921 14603
rect 36596 14572 36921 14600
rect 36596 14560 36602 14572
rect 36909 14569 36921 14572
rect 36955 14569 36967 14603
rect 39298 14600 39304 14612
rect 36909 14563 36967 14569
rect 37108 14572 39304 14600
rect 27614 14492 27620 14544
rect 27672 14532 27678 14544
rect 32585 14535 32643 14541
rect 32585 14532 32597 14535
rect 27672 14504 32597 14532
rect 27672 14492 27678 14504
rect 32585 14501 32597 14504
rect 32631 14501 32643 14535
rect 32585 14495 32643 14501
rect 34974 14492 34980 14544
rect 35032 14532 35038 14544
rect 35437 14535 35495 14541
rect 35437 14532 35449 14535
rect 35032 14504 35449 14532
rect 35032 14492 35038 14504
rect 35437 14501 35449 14504
rect 35483 14501 35495 14535
rect 35986 14532 35992 14544
rect 35437 14495 35495 14501
rect 35912 14504 35992 14532
rect 28166 14464 28172 14476
rect 28127 14436 28172 14464
rect 28166 14424 28172 14436
rect 28224 14424 28230 14476
rect 28261 14467 28319 14473
rect 28261 14433 28273 14467
rect 28307 14464 28319 14467
rect 28994 14464 29000 14476
rect 28307 14436 29000 14464
rect 28307 14433 28319 14436
rect 28261 14427 28319 14433
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 30837 14467 30895 14473
rect 30837 14433 30849 14467
rect 30883 14464 30895 14467
rect 31202 14464 31208 14476
rect 30883 14436 31208 14464
rect 30883 14433 30895 14436
rect 30837 14427 30895 14433
rect 31202 14424 31208 14436
rect 31260 14424 31266 14476
rect 35710 14424 35716 14476
rect 35768 14424 35774 14476
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 24210 14396 24216 14408
rect 23891 14368 24216 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14396 25099 14399
rect 25590 14396 25596 14408
rect 25087 14368 25596 14396
rect 25087 14365 25099 14368
rect 25041 14359 25099 14365
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 27525 14399 27583 14405
rect 27525 14365 27537 14399
rect 27571 14396 27583 14399
rect 28353 14399 28411 14405
rect 28353 14396 28365 14399
rect 27571 14368 28365 14396
rect 27571 14365 27583 14368
rect 27525 14359 27583 14365
rect 28353 14365 28365 14368
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28445 14399 28503 14405
rect 28445 14365 28457 14399
rect 28491 14396 28503 14399
rect 28902 14396 28908 14408
rect 28491 14368 28908 14396
rect 28491 14365 28503 14368
rect 28445 14359 28503 14365
rect 28368 14328 28396 14359
rect 28902 14356 28908 14368
rect 28960 14356 28966 14408
rect 30558 14396 30564 14408
rect 30519 14368 30564 14396
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 31389 14399 31447 14405
rect 31389 14396 31401 14399
rect 31036 14368 31401 14396
rect 29178 14328 29184 14340
rect 28368 14300 29184 14328
rect 29178 14288 29184 14300
rect 29236 14288 29242 14340
rect 31036 14272 31064 14368
rect 31389 14365 31401 14368
rect 31435 14365 31447 14399
rect 31570 14396 31576 14408
rect 31531 14368 31576 14396
rect 31389 14359 31447 14365
rect 31570 14356 31576 14368
rect 31628 14356 31634 14408
rect 34054 14396 34060 14408
rect 34015 14368 34060 14396
rect 34054 14356 34060 14368
rect 34112 14356 34118 14408
rect 34330 14396 34336 14408
rect 34243 14368 34336 14396
rect 34330 14356 34336 14368
rect 34388 14396 34394 14408
rect 35621 14399 35679 14405
rect 34388 14368 34928 14396
rect 34388 14356 34394 14368
rect 32766 14328 32772 14340
rect 32727 14300 32772 14328
rect 32766 14288 32772 14300
rect 32824 14288 32830 14340
rect 32950 14328 32956 14340
rect 32911 14300 32956 14328
rect 32950 14288 32956 14300
rect 33008 14288 33014 14340
rect 34900 14337 34928 14368
rect 35621 14365 35633 14399
rect 35667 14396 35679 14399
rect 35728 14396 35756 14424
rect 35667 14368 35756 14396
rect 35805 14399 35863 14405
rect 35667 14365 35679 14368
rect 35621 14359 35679 14365
rect 35805 14365 35817 14399
rect 35851 14396 35863 14399
rect 35912 14396 35940 14504
rect 35986 14492 35992 14504
rect 36044 14492 36050 14544
rect 36262 14464 36268 14476
rect 36004 14436 36268 14464
rect 36004 14405 36032 14436
rect 36262 14424 36268 14436
rect 36320 14424 36326 14476
rect 35851 14368 35940 14396
rect 35989 14399 36047 14405
rect 35851 14365 35863 14368
rect 35805 14359 35863 14365
rect 35989 14365 36001 14399
rect 36035 14365 36047 14399
rect 35989 14359 36047 14365
rect 36078 14356 36084 14408
rect 36136 14396 36142 14408
rect 36136 14368 36181 14396
rect 36136 14356 36142 14368
rect 36906 14356 36912 14408
rect 36964 14396 36970 14408
rect 37001 14399 37059 14405
rect 37001 14396 37013 14399
rect 36964 14368 37013 14396
rect 36964 14356 36970 14368
rect 37001 14365 37013 14368
rect 37047 14365 37059 14399
rect 37001 14359 37059 14365
rect 34885 14331 34943 14337
rect 34885 14297 34897 14331
rect 34931 14328 34943 14331
rect 35713 14331 35771 14337
rect 34931 14300 35480 14328
rect 34931 14297 34943 14300
rect 34885 14291 34943 14297
rect 23750 14260 23756 14272
rect 23711 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 25406 14220 25412 14272
rect 25464 14260 25470 14272
rect 25501 14263 25559 14269
rect 25501 14260 25513 14263
rect 25464 14232 25513 14260
rect 25464 14220 25470 14232
rect 25501 14229 25513 14232
rect 25547 14229 25559 14263
rect 25501 14223 25559 14229
rect 30653 14263 30711 14269
rect 30653 14229 30665 14263
rect 30699 14260 30711 14263
rect 31018 14260 31024 14272
rect 30699 14232 31024 14260
rect 30699 14229 30711 14232
rect 30653 14223 30711 14229
rect 31018 14220 31024 14232
rect 31076 14220 31082 14272
rect 33870 14260 33876 14272
rect 33831 14232 33876 14260
rect 33870 14220 33876 14232
rect 33928 14220 33934 14272
rect 35452 14260 35480 14300
rect 35713 14297 35725 14331
rect 35759 14328 35771 14331
rect 36354 14328 36360 14340
rect 35759 14300 36360 14328
rect 35759 14297 35771 14300
rect 35713 14291 35771 14297
rect 36354 14288 36360 14300
rect 36412 14288 36418 14340
rect 37108 14260 37136 14572
rect 39298 14560 39304 14572
rect 39356 14560 39362 14612
rect 39393 14603 39451 14609
rect 39393 14569 39405 14603
rect 39439 14600 39451 14603
rect 39574 14600 39580 14612
rect 39439 14572 39580 14600
rect 39439 14569 39451 14572
rect 39393 14563 39451 14569
rect 39574 14560 39580 14572
rect 39632 14560 39638 14612
rect 39850 14560 39856 14612
rect 39908 14600 39914 14612
rect 40037 14603 40095 14609
rect 40037 14600 40049 14603
rect 39908 14572 40049 14600
rect 39908 14560 39914 14572
rect 40037 14569 40049 14572
rect 40083 14569 40095 14603
rect 40037 14563 40095 14569
rect 42889 14603 42947 14609
rect 42889 14569 42901 14603
rect 42935 14600 42947 14603
rect 43438 14600 43444 14612
rect 42935 14572 43444 14600
rect 42935 14569 42947 14572
rect 42889 14563 42947 14569
rect 43438 14560 43444 14572
rect 43496 14600 43502 14612
rect 43806 14600 43812 14612
rect 43496 14572 43812 14600
rect 43496 14560 43502 14572
rect 43806 14560 43812 14572
rect 43864 14560 43870 14612
rect 45281 14603 45339 14609
rect 45281 14569 45293 14603
rect 45327 14600 45339 14603
rect 45370 14600 45376 14612
rect 45327 14572 45376 14600
rect 45327 14569 45339 14572
rect 45281 14563 45339 14569
rect 38286 14532 38292 14544
rect 38028 14504 38292 14532
rect 38028 14473 38056 14504
rect 38286 14492 38292 14504
rect 38344 14492 38350 14544
rect 38470 14492 38476 14544
rect 38528 14532 38534 14544
rect 43346 14532 43352 14544
rect 38528 14504 43352 14532
rect 38528 14492 38534 14504
rect 43346 14492 43352 14504
rect 43404 14492 43410 14544
rect 37921 14467 37979 14473
rect 37921 14464 37933 14467
rect 37661 14436 37933 14464
rect 37185 14399 37243 14405
rect 37185 14365 37197 14399
rect 37231 14396 37243 14399
rect 37550 14396 37556 14408
rect 37231 14368 37556 14396
rect 37231 14365 37243 14368
rect 37185 14359 37243 14365
rect 37550 14356 37556 14368
rect 37608 14356 37614 14408
rect 37661 14328 37689 14436
rect 37921 14433 37933 14436
rect 37967 14433 37979 14467
rect 37921 14427 37979 14433
rect 38013 14467 38071 14473
rect 38013 14433 38025 14467
rect 38059 14433 38071 14467
rect 38013 14427 38071 14433
rect 38378 14424 38384 14476
rect 38436 14464 38442 14476
rect 39482 14464 39488 14476
rect 38436 14436 39488 14464
rect 38436 14424 38442 14436
rect 39482 14424 39488 14436
rect 39540 14424 39546 14476
rect 40678 14464 40684 14476
rect 40639 14436 40684 14464
rect 40678 14424 40684 14436
rect 40736 14424 40742 14476
rect 41966 14464 41972 14476
rect 41524 14436 41972 14464
rect 37826 14396 37832 14408
rect 37787 14368 37832 14396
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 38105 14399 38163 14405
rect 38105 14365 38117 14399
rect 38151 14396 38163 14399
rect 40865 14399 40923 14405
rect 38151 14368 38240 14396
rect 38151 14365 38163 14368
rect 38105 14359 38163 14365
rect 38212 14340 38240 14368
rect 38396 14368 39344 14396
rect 38010 14328 38016 14340
rect 37661 14300 38016 14328
rect 38010 14288 38016 14300
rect 38068 14288 38074 14340
rect 38194 14288 38200 14340
rect 38252 14328 38258 14340
rect 38396 14328 38424 14368
rect 38252 14300 38424 14328
rect 38252 14288 38258 14300
rect 38562 14288 38568 14340
rect 38620 14328 38626 14340
rect 38620 14300 38884 14328
rect 38620 14288 38626 14300
rect 37642 14260 37648 14272
rect 35452 14232 37136 14260
rect 37603 14232 37648 14260
rect 37642 14220 37648 14232
rect 37700 14220 37706 14272
rect 38286 14220 38292 14272
rect 38344 14260 38350 14272
rect 38654 14260 38660 14272
rect 38344 14232 38660 14260
rect 38344 14220 38350 14232
rect 38654 14220 38660 14232
rect 38712 14220 38718 14272
rect 38856 14260 38884 14300
rect 38930 14288 38936 14340
rect 38988 14328 38994 14340
rect 39025 14331 39083 14337
rect 39025 14328 39037 14331
rect 38988 14300 39037 14328
rect 38988 14288 38994 14300
rect 39025 14297 39037 14300
rect 39071 14297 39083 14331
rect 39206 14328 39212 14340
rect 39167 14300 39212 14328
rect 39025 14291 39083 14297
rect 39206 14288 39212 14300
rect 39264 14288 39270 14340
rect 39316 14328 39344 14368
rect 40865 14365 40877 14399
rect 40911 14396 40923 14399
rect 40954 14396 40960 14408
rect 40911 14368 40960 14396
rect 40911 14365 40923 14368
rect 40865 14359 40923 14365
rect 40954 14356 40960 14368
rect 41012 14356 41018 14408
rect 41046 14356 41052 14408
rect 41104 14396 41110 14408
rect 41524 14405 41552 14436
rect 41966 14424 41972 14436
rect 42024 14424 42030 14476
rect 42150 14464 42156 14476
rect 42111 14436 42156 14464
rect 42150 14424 42156 14436
rect 42208 14424 42214 14476
rect 41509 14399 41567 14405
rect 41104 14368 41149 14396
rect 41104 14356 41110 14368
rect 41509 14365 41521 14399
rect 41555 14365 41567 14399
rect 41509 14359 41567 14365
rect 41524 14328 41552 14359
rect 41598 14356 41604 14408
rect 41656 14396 41662 14408
rect 41877 14399 41935 14405
rect 41877 14396 41889 14399
rect 41656 14368 41889 14396
rect 41656 14356 41662 14368
rect 41877 14365 41889 14368
rect 41923 14365 41935 14399
rect 41877 14359 41935 14365
rect 42610 14356 42616 14408
rect 42668 14396 42674 14408
rect 42889 14399 42947 14405
rect 42889 14396 42901 14399
rect 42668 14368 42901 14396
rect 42668 14356 42674 14368
rect 42889 14365 42901 14368
rect 42935 14365 42947 14399
rect 42889 14359 42947 14365
rect 43073 14399 43131 14405
rect 43073 14365 43085 14399
rect 43119 14396 43131 14399
rect 43530 14396 43536 14408
rect 43119 14368 43536 14396
rect 43119 14365 43131 14368
rect 43073 14359 43131 14365
rect 43530 14356 43536 14368
rect 43588 14356 43594 14408
rect 44361 14399 44419 14405
rect 44361 14365 44373 14399
rect 44407 14396 44419 14399
rect 44450 14396 44456 14408
rect 44407 14368 44456 14396
rect 44407 14365 44419 14368
rect 44361 14359 44419 14365
rect 44450 14356 44456 14368
rect 44508 14356 44514 14408
rect 44545 14399 44603 14405
rect 44545 14365 44557 14399
rect 44591 14396 44603 14399
rect 45296 14396 45324 14563
rect 45370 14560 45376 14572
rect 45428 14560 45434 14612
rect 44591 14368 45324 14396
rect 44591 14365 44603 14368
rect 44545 14359 44603 14365
rect 39316 14300 41552 14328
rect 41322 14260 41328 14272
rect 38856 14232 41328 14260
rect 41322 14220 41328 14232
rect 41380 14220 41386 14272
rect 44266 14220 44272 14272
rect 44324 14260 44330 14272
rect 44453 14263 44511 14269
rect 44453 14260 44465 14263
rect 44324 14232 44465 14260
rect 44324 14220 44330 14232
rect 44453 14229 44465 14232
rect 44499 14229 44511 14263
rect 44453 14223 44511 14229
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23750 14056 23756 14068
rect 23523 14028 23756 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 26053 14059 26111 14065
rect 26053 14056 26065 14059
rect 23900 14028 26065 14056
rect 23900 14016 23906 14028
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 24670 13988 24676 14000
rect 22879 13960 24676 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 24670 13948 24676 13960
rect 24728 13948 24734 14000
rect 22741 13923 22799 13929
rect 22741 13889 22753 13923
rect 22787 13920 22799 13923
rect 22925 13923 22983 13929
rect 22787 13892 22876 13920
rect 22787 13889 22799 13892
rect 22741 13883 22799 13889
rect 22848 13784 22876 13892
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 23382 13920 23388 13932
rect 23343 13892 23388 13920
rect 22925 13883 22983 13889
rect 22940 13852 22968 13883
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23661 13923 23719 13929
rect 23661 13920 23673 13923
rect 23532 13892 23673 13920
rect 23532 13880 23538 13892
rect 23661 13889 23673 13892
rect 23707 13889 23719 13923
rect 24394 13920 24400 13932
rect 24355 13892 24400 13920
rect 23661 13883 23719 13889
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 24581 13923 24639 13929
rect 24581 13889 24593 13923
rect 24627 13920 24639 13923
rect 24780 13920 24808 14028
rect 26053 14025 26065 14028
rect 26099 14025 26111 14059
rect 27798 14056 27804 14068
rect 26053 14019 26111 14025
rect 26252 14028 27804 14056
rect 25406 13948 25412 14000
rect 25464 13988 25470 14000
rect 26145 13991 26203 13997
rect 26145 13988 26157 13991
rect 25464 13960 25633 13988
rect 25464 13948 25470 13960
rect 25605 13954 25633 13960
rect 25700 13960 26157 13988
rect 25700 13954 25728 13960
rect 24627 13892 24808 13920
rect 25317 13923 25375 13929
rect 24627 13889 24639 13892
rect 24581 13883 24639 13889
rect 25317 13889 25329 13923
rect 25363 13889 25375 13923
rect 25498 13920 25504 13932
rect 25459 13892 25504 13920
rect 25317 13883 25375 13889
rect 23492 13852 23520 13880
rect 23842 13852 23848 13864
rect 22940 13824 23520 13852
rect 23584 13824 23848 13852
rect 23584 13784 23612 13824
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 24302 13852 24308 13864
rect 24263 13824 24308 13852
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 24412 13852 24440 13880
rect 25130 13852 25136 13864
rect 24412 13824 25136 13852
rect 25130 13812 25136 13824
rect 25188 13812 25194 13864
rect 25332 13852 25360 13883
rect 25498 13880 25504 13892
rect 25556 13880 25562 13932
rect 25605 13929 25728 13954
rect 26145 13957 26157 13960
rect 26191 13957 26203 13991
rect 26145 13951 26203 13957
rect 25593 13926 25728 13929
rect 25593 13923 25651 13926
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 25774 13880 25780 13932
rect 25832 13920 25838 13932
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 25832 13892 26065 13920
rect 25832 13880 25838 13892
rect 26053 13889 26065 13892
rect 26099 13920 26111 13923
rect 26252 13920 26280 14028
rect 27798 14016 27804 14028
rect 27856 14016 27862 14068
rect 29273 14059 29331 14065
rect 29273 14025 29285 14059
rect 29319 14025 29331 14059
rect 29638 14056 29644 14068
rect 29599 14028 29644 14056
rect 29273 14019 29331 14025
rect 28721 13991 28779 13997
rect 28721 13957 28733 13991
rect 28767 13988 28779 13991
rect 29178 13988 29184 14000
rect 28767 13960 29184 13988
rect 28767 13957 28779 13960
rect 28721 13951 28779 13957
rect 29178 13948 29184 13960
rect 29236 13948 29242 14000
rect 26099 13892 26280 13920
rect 26329 13923 26387 13929
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 26375 13892 26409 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 26344 13852 26372 13883
rect 27246 13880 27252 13932
rect 27304 13920 27310 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 27304 13892 27353 13920
rect 27304 13880 27310 13892
rect 27341 13889 27353 13892
rect 27387 13920 27399 13923
rect 28353 13923 28411 13929
rect 28353 13920 28365 13923
rect 27387 13892 28365 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 28353 13889 28365 13892
rect 28399 13889 28411 13923
rect 28534 13920 28540 13932
rect 28495 13892 28540 13920
rect 28353 13883 28411 13889
rect 28534 13880 28540 13892
rect 28592 13880 28598 13932
rect 28813 13923 28871 13929
rect 28813 13889 28825 13923
rect 28859 13920 28871 13923
rect 29288 13920 29316 14019
rect 29638 14016 29644 14028
rect 29696 14016 29702 14068
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 31113 14059 31171 14065
rect 31113 14056 31125 14059
rect 30892 14028 31125 14056
rect 30892 14016 30898 14028
rect 31113 14025 31125 14028
rect 31159 14025 31171 14059
rect 31113 14019 31171 14025
rect 31202 14016 31208 14068
rect 31260 14056 31266 14068
rect 32769 14059 32827 14065
rect 31260 14028 31305 14056
rect 31260 14016 31266 14028
rect 32769 14025 32781 14059
rect 32815 14056 32827 14059
rect 32950 14056 32956 14068
rect 32815 14028 32956 14056
rect 32815 14025 32827 14028
rect 32769 14019 32827 14025
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 34333 14059 34391 14065
rect 34333 14025 34345 14059
rect 34379 14056 34391 14059
rect 34422 14056 34428 14068
rect 34379 14028 34428 14056
rect 34379 14025 34391 14028
rect 34333 14019 34391 14025
rect 34422 14016 34428 14028
rect 34480 14016 34486 14068
rect 36446 14056 36452 14068
rect 36407 14028 36452 14056
rect 36446 14016 36452 14028
rect 36504 14016 36510 14068
rect 36538 14016 36544 14068
rect 36596 14056 36602 14068
rect 40310 14056 40316 14068
rect 36596 14028 40316 14056
rect 36596 14016 36602 14028
rect 40310 14016 40316 14028
rect 40368 14016 40374 14068
rect 40770 14016 40776 14068
rect 40828 14056 40834 14068
rect 40957 14059 41015 14065
rect 40957 14056 40969 14059
rect 40828 14028 40969 14056
rect 40828 14016 40834 14028
rect 40957 14025 40969 14028
rect 41003 14025 41015 14059
rect 41874 14056 41880 14068
rect 40957 14019 41015 14025
rect 41708 14028 41880 14056
rect 29733 13991 29791 13997
rect 29733 13957 29745 13991
rect 29779 13988 29791 13991
rect 31481 13991 31539 13997
rect 31481 13988 31493 13991
rect 29779 13960 31493 13988
rect 29779 13957 29791 13960
rect 29733 13951 29791 13957
rect 31128 13932 31156 13960
rect 31481 13957 31493 13960
rect 31527 13988 31539 13991
rect 31846 13988 31852 14000
rect 31527 13960 31852 13988
rect 31527 13957 31539 13960
rect 31481 13951 31539 13957
rect 31846 13948 31852 13960
rect 31904 13948 31910 14000
rect 35084 13960 35572 13988
rect 28859 13892 29316 13920
rect 28859 13889 28871 13892
rect 28813 13883 28871 13889
rect 30558 13880 30564 13932
rect 30616 13920 30622 13932
rect 30929 13923 30987 13929
rect 30929 13920 30941 13923
rect 30616 13892 30941 13920
rect 30616 13880 30622 13892
rect 30929 13889 30941 13892
rect 30975 13889 30987 13923
rect 30929 13883 30987 13889
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 31294 13920 31300 13932
rect 31255 13892 31300 13920
rect 31294 13880 31300 13892
rect 31352 13880 31358 13932
rect 33042 13920 33048 13932
rect 33003 13892 33048 13920
rect 33042 13880 33048 13892
rect 33100 13880 33106 13932
rect 33226 13920 33232 13932
rect 33187 13892 33232 13920
rect 33226 13880 33232 13892
rect 33284 13920 33290 13932
rect 33778 13920 33784 13932
rect 33284 13892 33784 13920
rect 33284 13880 33290 13892
rect 33778 13880 33784 13892
rect 33836 13880 33842 13932
rect 34974 13920 34980 13932
rect 34935 13892 34980 13920
rect 34974 13880 34980 13892
rect 35032 13880 35038 13932
rect 35084 13929 35112 13960
rect 35069 13923 35127 13929
rect 35069 13889 35081 13923
rect 35115 13889 35127 13923
rect 35250 13920 35256 13932
rect 35211 13892 35256 13920
rect 35069 13883 35127 13889
rect 35250 13880 35256 13892
rect 35308 13880 35314 13932
rect 35342 13880 35348 13932
rect 35400 13920 35406 13932
rect 35544 13920 35572 13960
rect 35710 13948 35716 14000
rect 35768 13988 35774 14000
rect 37737 13991 37795 13997
rect 37737 13988 37749 13991
rect 35768 13960 37749 13988
rect 35768 13948 35774 13960
rect 37737 13957 37749 13960
rect 37783 13957 37795 13991
rect 37737 13951 37795 13957
rect 37826 13948 37832 14000
rect 37884 13988 37890 14000
rect 38378 13988 38384 14000
rect 37884 13960 38384 13988
rect 37884 13948 37890 13960
rect 36447 13923 36505 13929
rect 36447 13920 36459 13923
rect 35400 13892 35445 13920
rect 35544 13892 36459 13920
rect 35400 13880 35406 13892
rect 36447 13889 36459 13892
rect 36493 13920 36505 13923
rect 36630 13920 36636 13932
rect 36493 13892 36636 13920
rect 36493 13889 36505 13892
rect 36447 13883 36505 13889
rect 36630 13880 36636 13892
rect 36688 13880 36694 13932
rect 37274 13880 37280 13932
rect 37332 13920 37338 13932
rect 37918 13920 37924 13932
rect 37332 13892 37780 13920
rect 37879 13892 37924 13920
rect 37332 13880 37338 13892
rect 26786 13852 26792 13864
rect 25332 13824 26792 13852
rect 26786 13812 26792 13824
rect 26844 13812 26850 13864
rect 27433 13855 27491 13861
rect 27433 13821 27445 13855
rect 27479 13852 27491 13855
rect 27982 13852 27988 13864
rect 27479 13824 27752 13852
rect 27479 13821 27491 13824
rect 27433 13815 27491 13821
rect 22848 13756 23612 13784
rect 23400 13728 23428 13756
rect 24026 13744 24032 13796
rect 24084 13784 24090 13796
rect 24762 13784 24768 13796
rect 24084 13756 24768 13784
rect 24084 13744 24090 13756
rect 24762 13744 24768 13756
rect 24820 13744 24826 13796
rect 27724 13784 27752 13824
rect 27908 13824 27988 13852
rect 27908 13784 27936 13824
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 29917 13855 29975 13861
rect 29917 13821 29929 13855
rect 29963 13821 29975 13855
rect 29917 13815 29975 13821
rect 27724 13756 27936 13784
rect 23382 13676 23388 13728
rect 23440 13676 23446 13728
rect 23842 13716 23848 13728
rect 23803 13688 23848 13716
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 27157 13719 27215 13725
rect 27157 13716 27169 13719
rect 26292 13688 27169 13716
rect 26292 13676 26298 13688
rect 27157 13685 27169 13688
rect 27203 13685 27215 13719
rect 29932 13716 29960 13815
rect 32858 13812 32864 13864
rect 32916 13852 32922 13864
rect 32953 13855 33011 13861
rect 32953 13852 32965 13855
rect 32916 13824 32965 13852
rect 32916 13812 32922 13824
rect 32953 13821 32965 13824
rect 32999 13821 33011 13855
rect 33134 13852 33140 13864
rect 33095 13824 33140 13852
rect 32953 13815 33011 13821
rect 33134 13812 33140 13824
rect 33192 13812 33198 13864
rect 34054 13812 34060 13864
rect 34112 13852 34118 13864
rect 36909 13855 36967 13861
rect 36909 13852 36921 13855
rect 34112 13824 36921 13852
rect 34112 13812 34118 13824
rect 36909 13821 36921 13824
rect 36955 13852 36967 13855
rect 37642 13852 37648 13864
rect 36955 13824 37648 13852
rect 36955 13821 36967 13824
rect 36909 13815 36967 13821
rect 37642 13812 37648 13824
rect 37700 13812 37706 13864
rect 37752 13852 37780 13892
rect 37918 13880 37924 13892
rect 37976 13880 37982 13932
rect 38028 13929 38056 13960
rect 38378 13948 38384 13960
rect 38436 13948 38442 14000
rect 38841 13991 38899 13997
rect 38841 13957 38853 13991
rect 38887 13988 38899 13991
rect 39206 13988 39212 14000
rect 38887 13960 39212 13988
rect 38887 13957 38899 13960
rect 38841 13951 38899 13957
rect 39206 13948 39212 13960
rect 39264 13988 39270 14000
rect 41138 13988 41144 14000
rect 39264 13960 41144 13988
rect 39264 13948 39270 13960
rect 38013 13923 38071 13929
rect 38013 13889 38025 13923
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 38102 13880 38108 13932
rect 38160 13920 38166 13932
rect 39684 13929 39712 13960
rect 41138 13948 41144 13960
rect 41196 13948 41202 14000
rect 41708 13997 41736 14028
rect 41874 14016 41880 14028
rect 41932 14056 41938 14068
rect 42058 14056 42064 14068
rect 41932 14028 42064 14056
rect 41932 14016 41938 14028
rect 42058 14016 42064 14028
rect 42116 14016 42122 14068
rect 44174 14016 44180 14068
rect 44232 14056 44238 14068
rect 44232 14028 45232 14056
rect 44232 14016 44238 14028
rect 41693 13991 41751 13997
rect 41693 13957 41705 13991
rect 41739 13957 41751 13991
rect 42978 13988 42984 14000
rect 42939 13960 42984 13988
rect 41693 13951 41751 13957
rect 42978 13948 42984 13960
rect 43036 13948 43042 14000
rect 44450 13948 44456 14000
rect 44508 13988 44514 14000
rect 44508 13960 44588 13988
rect 44508 13948 44514 13960
rect 38749 13923 38807 13929
rect 38749 13920 38761 13923
rect 38160 13892 38761 13920
rect 38160 13880 38166 13892
rect 38749 13889 38761 13892
rect 38795 13889 38807 13923
rect 38749 13883 38807 13889
rect 39669 13923 39727 13929
rect 39669 13889 39681 13923
rect 39715 13889 39727 13923
rect 39669 13883 39727 13889
rect 40678 13880 40684 13932
rect 40736 13920 40742 13932
rect 40822 13926 40880 13929
rect 40954 13926 40960 13932
rect 40822 13923 40960 13926
rect 40736 13892 40781 13920
rect 40736 13880 40742 13892
rect 40822 13889 40834 13923
rect 40868 13898 40960 13923
rect 40868 13892 40885 13898
rect 40868 13889 40880 13892
rect 40822 13883 40880 13889
rect 40954 13880 40960 13898
rect 41012 13880 41018 13932
rect 41049 13923 41107 13929
rect 41049 13889 41061 13923
rect 41095 13920 41107 13923
rect 41322 13920 41328 13932
rect 41095 13892 41328 13920
rect 41095 13889 41107 13892
rect 41049 13883 41107 13889
rect 41322 13880 41328 13892
rect 41380 13880 41386 13932
rect 41877 13923 41935 13929
rect 41877 13889 41889 13923
rect 41923 13920 41935 13923
rect 41966 13920 41972 13932
rect 41923 13892 41972 13920
rect 41923 13889 41935 13892
rect 41877 13883 41935 13889
rect 41966 13880 41972 13892
rect 42024 13880 42030 13932
rect 42610 13920 42616 13932
rect 42523 13892 42616 13920
rect 42610 13880 42616 13892
rect 42668 13880 42674 13932
rect 42889 13923 42947 13929
rect 42889 13889 42901 13923
rect 42935 13918 42947 13923
rect 43530 13920 43536 13932
rect 43042 13918 43536 13920
rect 42935 13892 43536 13918
rect 42935 13890 43070 13892
rect 42935 13889 42947 13890
rect 42889 13883 42947 13889
rect 43530 13880 43536 13892
rect 43588 13880 43594 13932
rect 44082 13920 44088 13932
rect 44043 13892 44088 13920
rect 44082 13880 44088 13892
rect 44140 13880 44146 13932
rect 44266 13920 44272 13932
rect 44227 13892 44272 13920
rect 44266 13880 44272 13892
rect 44324 13880 44330 13932
rect 44358 13880 44364 13932
rect 44416 13920 44422 13932
rect 44560 13929 44588 13960
rect 44545 13923 44603 13929
rect 44416 13892 44509 13920
rect 44416 13880 44422 13892
rect 44545 13889 44557 13923
rect 44591 13889 44603 13923
rect 44545 13883 44603 13889
rect 44634 13880 44640 13932
rect 44692 13920 44698 13932
rect 45204 13929 45232 14028
rect 45005 13923 45063 13929
rect 45005 13920 45017 13923
rect 44692 13892 45017 13920
rect 44692 13880 44698 13892
rect 45005 13889 45017 13892
rect 45051 13889 45063 13923
rect 45005 13883 45063 13889
rect 45189 13923 45247 13929
rect 45189 13889 45201 13923
rect 45235 13920 45247 13923
rect 45462 13920 45468 13932
rect 45235 13892 45468 13920
rect 45235 13889 45247 13892
rect 45189 13883 45247 13889
rect 45462 13880 45468 13892
rect 45520 13880 45526 13932
rect 40310 13852 40316 13864
rect 37752 13824 40316 13852
rect 40310 13812 40316 13824
rect 40368 13812 40374 13864
rect 41138 13812 41144 13864
rect 41196 13852 41202 13864
rect 42628 13852 42656 13880
rect 41196 13824 42656 13852
rect 41196 13812 41202 13824
rect 42702 13812 42708 13864
rect 42760 13852 42766 13864
rect 44177 13855 44235 13861
rect 44177 13852 44189 13855
rect 42760 13824 44189 13852
rect 42760 13812 42766 13824
rect 44177 13821 44189 13824
rect 44223 13821 44235 13855
rect 44376 13852 44404 13880
rect 45738 13852 45744 13864
rect 44376 13824 45744 13852
rect 44177 13815 44235 13821
rect 45738 13812 45744 13824
rect 45796 13812 45802 13864
rect 30374 13744 30380 13796
rect 30432 13784 30438 13796
rect 30650 13784 30656 13796
rect 30432 13756 30656 13784
rect 30432 13744 30438 13756
rect 30650 13744 30656 13756
rect 30708 13744 30714 13796
rect 36817 13787 36875 13793
rect 36817 13753 36829 13787
rect 36863 13784 36875 13787
rect 43622 13784 43628 13796
rect 36863 13756 43628 13784
rect 36863 13753 36875 13756
rect 36817 13747 36875 13753
rect 43622 13744 43628 13756
rect 43680 13744 43686 13796
rect 44450 13744 44456 13796
rect 44508 13784 44514 13796
rect 45646 13784 45652 13796
rect 44508 13756 45652 13784
rect 44508 13744 44514 13756
rect 45646 13744 45652 13756
rect 45704 13744 45710 13796
rect 33870 13716 33876 13728
rect 29932 13688 33876 13716
rect 27157 13679 27215 13685
rect 33870 13676 33876 13688
rect 33928 13676 33934 13728
rect 34790 13716 34796 13728
rect 34751 13688 34796 13716
rect 34790 13676 34796 13688
rect 34848 13676 34854 13728
rect 36265 13719 36323 13725
rect 36265 13685 36277 13719
rect 36311 13716 36323 13719
rect 36354 13716 36360 13728
rect 36311 13688 36360 13716
rect 36311 13685 36323 13688
rect 36265 13679 36323 13685
rect 36354 13676 36360 13688
rect 36412 13676 36418 13728
rect 37734 13716 37740 13728
rect 37695 13688 37740 13716
rect 37734 13676 37740 13688
rect 37792 13676 37798 13728
rect 39298 13676 39304 13728
rect 39356 13716 39362 13728
rect 39485 13719 39543 13725
rect 39485 13716 39497 13719
rect 39356 13688 39497 13716
rect 39356 13676 39362 13688
rect 39485 13685 39497 13688
rect 39531 13685 39543 13719
rect 39485 13679 39543 13685
rect 40681 13719 40739 13725
rect 40681 13685 40693 13719
rect 40727 13716 40739 13719
rect 41230 13716 41236 13728
rect 40727 13688 41236 13716
rect 40727 13685 40739 13688
rect 40681 13679 40739 13685
rect 41230 13676 41236 13688
rect 41288 13676 41294 13728
rect 41506 13716 41512 13728
rect 41467 13688 41512 13716
rect 41506 13676 41512 13688
rect 41564 13676 41570 13728
rect 42150 13676 42156 13728
rect 42208 13716 42214 13728
rect 43901 13719 43959 13725
rect 43901 13716 43913 13719
rect 42208 13688 43913 13716
rect 42208 13676 42214 13688
rect 43901 13685 43913 13688
rect 43947 13685 43959 13719
rect 45002 13716 45008 13728
rect 44963 13688 45008 13716
rect 43901 13679 43959 13685
rect 45002 13676 45008 13688
rect 45060 13676 45066 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 28534 13472 28540 13524
rect 28592 13512 28598 13524
rect 28905 13515 28963 13521
rect 28905 13512 28917 13515
rect 28592 13484 28917 13512
rect 28592 13472 28598 13484
rect 28905 13481 28917 13484
rect 28951 13481 28963 13515
rect 28905 13475 28963 13481
rect 29825 13515 29883 13521
rect 29825 13481 29837 13515
rect 29871 13512 29883 13515
rect 30466 13512 30472 13524
rect 29871 13484 30472 13512
rect 29871 13481 29883 13484
rect 29825 13475 29883 13481
rect 30466 13472 30472 13484
rect 30524 13472 30530 13524
rect 31018 13512 31024 13524
rect 30979 13484 31024 13512
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 32766 13472 32772 13524
rect 32824 13512 32830 13524
rect 32861 13515 32919 13521
rect 32861 13512 32873 13515
rect 32824 13484 32873 13512
rect 32824 13472 32830 13484
rect 32861 13481 32873 13484
rect 32907 13481 32919 13515
rect 32861 13475 32919 13481
rect 33042 13472 33048 13524
rect 33100 13512 33106 13524
rect 33597 13515 33655 13521
rect 33597 13512 33609 13515
rect 33100 13484 33609 13512
rect 33100 13472 33106 13484
rect 33597 13481 33609 13484
rect 33643 13481 33655 13515
rect 33597 13475 33655 13481
rect 33873 13515 33931 13521
rect 33873 13481 33885 13515
rect 33919 13512 33931 13515
rect 35526 13512 35532 13524
rect 33919 13484 35532 13512
rect 33919 13481 33931 13484
rect 33873 13475 33931 13481
rect 35526 13472 35532 13484
rect 35584 13472 35590 13524
rect 36446 13512 36452 13524
rect 36407 13484 36452 13512
rect 36446 13472 36452 13484
rect 36504 13472 36510 13524
rect 38841 13515 38899 13521
rect 36924 13484 38056 13512
rect 26786 13444 26792 13456
rect 26747 13416 26792 13444
rect 26786 13404 26792 13416
rect 26844 13404 26850 13456
rect 30377 13447 30435 13453
rect 30377 13444 30389 13447
rect 26988 13416 30389 13444
rect 23750 13376 23756 13388
rect 23711 13348 23756 13376
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 25130 13376 25136 13388
rect 25091 13348 25136 13376
rect 25130 13336 25136 13348
rect 25188 13336 25194 13388
rect 23382 13308 23388 13320
rect 23343 13280 23388 13308
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13308 23535 13311
rect 24394 13308 24400 13320
rect 23523 13280 24400 13308
rect 23523 13277 23535 13280
rect 23477 13271 23535 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 25225 13311 25283 13317
rect 24811 13280 25176 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 25148 13240 25176 13280
rect 25225 13277 25237 13311
rect 25271 13308 25283 13311
rect 25866 13308 25872 13320
rect 25271 13280 25872 13308
rect 25271 13277 25283 13280
rect 25225 13271 25283 13277
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13308 26111 13311
rect 26234 13308 26240 13320
rect 26099 13280 26240 13308
rect 26099 13277 26111 13280
rect 26053 13271 26111 13277
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26326 13268 26332 13320
rect 26384 13308 26390 13320
rect 26988 13308 27016 13416
rect 30377 13413 30389 13416
rect 30423 13413 30435 13447
rect 30377 13407 30435 13413
rect 32490 13404 32496 13456
rect 32548 13444 32554 13456
rect 32950 13444 32956 13456
rect 32548 13416 32956 13444
rect 32548 13404 32554 13416
rect 32950 13404 32956 13416
rect 33008 13404 33014 13456
rect 35618 13404 35624 13456
rect 35676 13404 35682 13456
rect 36262 13404 36268 13456
rect 36320 13444 36326 13456
rect 36630 13444 36636 13456
rect 36320 13416 36636 13444
rect 36320 13404 36326 13416
rect 36630 13404 36636 13416
rect 36688 13444 36694 13456
rect 36817 13447 36875 13453
rect 36817 13444 36829 13447
rect 36688 13416 36829 13444
rect 36688 13404 36694 13416
rect 36817 13413 36829 13416
rect 36863 13413 36875 13447
rect 36817 13407 36875 13413
rect 27246 13376 27252 13388
rect 27207 13348 27252 13376
rect 27246 13336 27252 13348
rect 27304 13336 27310 13388
rect 27801 13379 27859 13385
rect 27801 13345 27813 13379
rect 27847 13376 27859 13379
rect 27890 13376 27896 13388
rect 27847 13348 27896 13376
rect 27847 13345 27859 13348
rect 27801 13339 27859 13345
rect 27890 13336 27896 13348
rect 27948 13376 27954 13388
rect 31018 13376 31024 13388
rect 27948 13348 31024 13376
rect 27948 13336 27954 13348
rect 31018 13336 31024 13348
rect 31076 13376 31082 13388
rect 31757 13379 31815 13385
rect 31757 13376 31769 13379
rect 31076 13348 31769 13376
rect 31076 13336 31082 13348
rect 31757 13345 31769 13348
rect 31803 13345 31815 13379
rect 31757 13339 31815 13345
rect 33226 13336 33232 13388
rect 33284 13376 33290 13388
rect 33284 13348 33916 13376
rect 33284 13336 33290 13348
rect 27154 13308 27160 13320
rect 26384 13280 27016 13308
rect 27115 13280 27160 13308
rect 26384 13268 26390 13280
rect 27154 13268 27160 13280
rect 27212 13268 27218 13320
rect 27985 13311 28043 13317
rect 27985 13277 27997 13311
rect 28031 13277 28043 13311
rect 28353 13311 28411 13317
rect 28353 13308 28365 13311
rect 27985 13271 28043 13277
rect 28092 13280 28365 13308
rect 23768 13212 24992 13240
rect 25148 13212 25912 13240
rect 23566 13172 23572 13184
rect 23527 13144 23572 13172
rect 23566 13132 23572 13144
rect 23624 13132 23630 13184
rect 23768 13181 23796 13212
rect 23753 13175 23811 13181
rect 23753 13141 23765 13175
rect 23799 13141 23811 13175
rect 23753 13135 23811 13141
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 24964 13181 24992 13212
rect 24857 13175 24915 13181
rect 24857 13172 24869 13175
rect 24728 13144 24869 13172
rect 24728 13132 24734 13144
rect 24857 13141 24869 13144
rect 24903 13141 24915 13175
rect 24857 13135 24915 13141
rect 24949 13175 25007 13181
rect 24949 13141 24961 13175
rect 24995 13141 25007 13175
rect 25406 13172 25412 13184
rect 25367 13144 25412 13172
rect 24949 13135 25007 13141
rect 25406 13132 25412 13144
rect 25464 13132 25470 13184
rect 25884 13181 25912 13212
rect 27246 13200 27252 13252
rect 27304 13240 27310 13252
rect 28000 13240 28028 13271
rect 27304 13212 28028 13240
rect 27304 13200 27310 13212
rect 25869 13175 25927 13181
rect 25869 13141 25881 13175
rect 25915 13141 25927 13175
rect 25869 13135 25927 13141
rect 26237 13175 26295 13181
rect 26237 13141 26249 13175
rect 26283 13172 26295 13175
rect 26418 13172 26424 13184
rect 26283 13144 26424 13172
rect 26283 13141 26295 13144
rect 26237 13135 26295 13141
rect 26418 13132 26424 13144
rect 26476 13172 26482 13184
rect 26878 13172 26884 13184
rect 26476 13144 26884 13172
rect 26476 13132 26482 13144
rect 26878 13132 26884 13144
rect 26936 13132 26942 13184
rect 27522 13132 27528 13184
rect 27580 13172 27586 13184
rect 28092 13172 28120 13280
rect 28353 13277 28365 13280
rect 28399 13277 28411 13311
rect 28353 13271 28411 13277
rect 28997 13311 29055 13317
rect 28997 13277 29009 13311
rect 29043 13308 29055 13311
rect 29454 13308 29460 13320
rect 29043 13280 29460 13308
rect 29043 13277 29055 13280
rect 28997 13271 29055 13277
rect 29454 13268 29460 13280
rect 29512 13308 29518 13320
rect 30190 13308 30196 13320
rect 29512 13280 30196 13308
rect 29512 13268 29518 13280
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13308 30343 13311
rect 30374 13308 30380 13320
rect 30331 13280 30380 13308
rect 30331 13277 30343 13280
rect 30285 13271 30343 13277
rect 30374 13268 30380 13280
rect 30432 13268 30438 13320
rect 30469 13311 30527 13317
rect 30469 13277 30481 13311
rect 30515 13308 30527 13311
rect 30742 13308 30748 13320
rect 30515 13280 30748 13308
rect 30515 13277 30527 13280
rect 30469 13271 30527 13277
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 31294 13308 31300 13320
rect 31255 13280 31300 13308
rect 31294 13268 31300 13280
rect 31352 13268 31358 13320
rect 32585 13311 32643 13317
rect 32585 13277 32597 13311
rect 32631 13308 32643 13311
rect 33042 13308 33048 13320
rect 32631 13280 33048 13308
rect 32631 13277 32643 13280
rect 32585 13271 32643 13277
rect 33042 13268 33048 13280
rect 33100 13268 33106 13320
rect 33781 13311 33839 13317
rect 33781 13277 33793 13311
rect 33827 13277 33839 13311
rect 33888 13308 33916 13348
rect 33962 13336 33968 13388
rect 34020 13376 34026 13388
rect 34238 13376 34244 13388
rect 34020 13348 34244 13376
rect 34020 13336 34026 13348
rect 34238 13336 34244 13348
rect 34296 13336 34302 13388
rect 35161 13379 35219 13385
rect 35161 13345 35173 13379
rect 35207 13376 35219 13379
rect 35636 13376 35664 13404
rect 36722 13376 36728 13388
rect 35207 13348 35664 13376
rect 36683 13348 36728 13376
rect 35207 13345 35219 13348
rect 35161 13339 35219 13345
rect 36722 13336 36728 13348
rect 36780 13336 36786 13388
rect 36924 13376 36952 13484
rect 37734 13404 37740 13456
rect 37792 13444 37798 13456
rect 37829 13447 37887 13453
rect 37829 13444 37841 13447
rect 37792 13416 37841 13444
rect 37792 13404 37798 13416
rect 37829 13413 37841 13416
rect 37875 13413 37887 13447
rect 37829 13407 37887 13413
rect 38028 13444 38056 13484
rect 38841 13481 38853 13515
rect 38887 13512 38899 13515
rect 39022 13512 39028 13524
rect 38887 13484 39028 13512
rect 38887 13481 38899 13484
rect 38841 13475 38899 13481
rect 39022 13472 39028 13484
rect 39080 13472 39086 13524
rect 40034 13472 40040 13524
rect 40092 13512 40098 13524
rect 40681 13515 40739 13521
rect 40681 13512 40693 13515
rect 40092 13484 40693 13512
rect 40092 13472 40098 13484
rect 40681 13481 40693 13484
rect 40727 13481 40739 13515
rect 40681 13475 40739 13481
rect 40770 13472 40776 13524
rect 40828 13512 40834 13524
rect 41417 13515 41475 13521
rect 41417 13512 41429 13515
rect 40828 13484 41429 13512
rect 40828 13472 40834 13484
rect 41417 13481 41429 13484
rect 41463 13512 41475 13515
rect 41463 13484 44128 13512
rect 41463 13481 41475 13484
rect 41417 13475 41475 13481
rect 38930 13444 38936 13456
rect 38028 13416 38936 13444
rect 36832 13348 36952 13376
rect 34149 13311 34207 13317
rect 34149 13308 34161 13311
rect 33888 13280 34161 13308
rect 33781 13271 33839 13277
rect 34149 13277 34161 13280
rect 34195 13308 34207 13311
rect 34422 13308 34428 13320
rect 34195 13280 34428 13308
rect 34195 13277 34207 13280
rect 34149 13271 34207 13277
rect 30558 13200 30564 13252
rect 30616 13240 30622 13252
rect 30926 13240 30932 13252
rect 30616 13212 30932 13240
rect 30616 13200 30622 13212
rect 30926 13200 30932 13212
rect 30984 13240 30990 13252
rect 31021 13243 31079 13249
rect 31021 13240 31033 13243
rect 30984 13212 31033 13240
rect 30984 13200 30990 13212
rect 31021 13209 31033 13212
rect 31067 13209 31079 13243
rect 32858 13240 32864 13252
rect 32819 13212 32864 13240
rect 31021 13203 31079 13209
rect 32858 13200 32864 13212
rect 32916 13200 32922 13252
rect 33796 13240 33824 13271
rect 34422 13268 34428 13280
rect 34480 13268 34486 13320
rect 35069 13311 35127 13317
rect 35069 13277 35081 13311
rect 35115 13277 35127 13311
rect 35069 13271 35127 13277
rect 35621 13311 35679 13317
rect 35621 13277 35633 13311
rect 35667 13308 35679 13311
rect 36633 13311 36691 13317
rect 36633 13308 36645 13311
rect 35667 13280 36645 13308
rect 35667 13277 35679 13280
rect 35621 13271 35679 13277
rect 36633 13277 36645 13280
rect 36679 13308 36691 13311
rect 36832 13308 36860 13348
rect 37458 13336 37464 13388
rect 37516 13376 37522 13388
rect 37921 13379 37979 13385
rect 37921 13376 37933 13379
rect 37516 13348 37933 13376
rect 37516 13336 37522 13348
rect 37921 13345 37933 13348
rect 37967 13345 37979 13379
rect 37921 13339 37979 13345
rect 36679 13280 36860 13308
rect 36909 13311 36967 13317
rect 36679 13277 36691 13280
rect 36633 13271 36691 13277
rect 36909 13277 36921 13311
rect 36955 13308 36967 13311
rect 37553 13311 37611 13317
rect 37553 13308 37565 13311
rect 36955 13280 37565 13308
rect 36955 13277 36967 13280
rect 36909 13271 36967 13277
rect 37553 13277 37565 13280
rect 37599 13277 37611 13311
rect 37734 13308 37740 13320
rect 37695 13280 37740 13308
rect 37553 13271 37611 13277
rect 34514 13240 34520 13252
rect 33796 13212 34520 13240
rect 34514 13200 34520 13212
rect 34572 13200 34578 13252
rect 27580 13144 28120 13172
rect 28261 13175 28319 13181
rect 27580 13132 27586 13144
rect 28261 13141 28273 13175
rect 28307 13172 28319 13175
rect 28534 13172 28540 13184
rect 28307 13144 28540 13172
rect 28307 13141 28319 13144
rect 28261 13135 28319 13141
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 30834 13132 30840 13184
rect 30892 13172 30898 13184
rect 31205 13175 31263 13181
rect 31205 13172 31217 13175
rect 30892 13144 31217 13172
rect 30892 13132 30898 13144
rect 31205 13141 31217 13144
rect 31251 13141 31263 13175
rect 31205 13135 31263 13141
rect 32677 13175 32735 13181
rect 32677 13141 32689 13175
rect 32723 13172 32735 13175
rect 33134 13172 33140 13184
rect 32723 13144 33140 13172
rect 32723 13141 32735 13144
rect 32677 13135 32735 13141
rect 33134 13132 33140 13144
rect 33192 13132 33198 13184
rect 35084 13172 35112 13271
rect 37568 13240 37596 13271
rect 37734 13268 37740 13280
rect 37792 13268 37798 13320
rect 38028 13317 38056 13416
rect 38930 13404 38936 13416
rect 38988 13404 38994 13456
rect 39206 13404 39212 13456
rect 39264 13444 39270 13456
rect 41969 13447 42027 13453
rect 41969 13444 41981 13447
rect 39264 13416 41981 13444
rect 39264 13404 39270 13416
rect 41969 13413 41981 13416
rect 42015 13413 42027 13447
rect 43254 13444 43260 13456
rect 43215 13416 43260 13444
rect 41969 13407 42027 13413
rect 43254 13404 43260 13416
rect 43312 13404 43318 13456
rect 43349 13447 43407 13453
rect 43349 13413 43361 13447
rect 43395 13444 43407 13447
rect 43993 13447 44051 13453
rect 43993 13444 44005 13447
rect 43395 13416 44005 13444
rect 43395 13413 43407 13416
rect 43349 13407 43407 13413
rect 43993 13413 44005 13416
rect 44039 13413 44051 13447
rect 43993 13407 44051 13413
rect 38746 13376 38752 13388
rect 38120 13348 38752 13376
rect 38013 13311 38071 13317
rect 38013 13277 38025 13311
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 38120 13240 38148 13348
rect 38746 13336 38752 13348
rect 38804 13336 38810 13388
rect 38838 13336 38844 13388
rect 38896 13336 38902 13388
rect 40494 13336 40500 13388
rect 40552 13376 40558 13388
rect 41233 13379 41291 13385
rect 41233 13376 41245 13379
rect 40552 13348 41245 13376
rect 40552 13336 40558 13348
rect 41233 13345 41245 13348
rect 41279 13345 41291 13379
rect 41233 13339 41291 13345
rect 42058 13336 42064 13388
rect 42116 13376 42122 13388
rect 42794 13376 42800 13388
rect 42116 13348 42800 13376
rect 42116 13336 42122 13348
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13308 38715 13311
rect 38856 13308 38884 13336
rect 40310 13308 40316 13320
rect 38703 13280 38884 13308
rect 40223 13280 40316 13308
rect 38703 13277 38715 13280
rect 38657 13271 38715 13277
rect 40310 13268 40316 13280
rect 40368 13308 40374 13320
rect 40368 13280 40632 13308
rect 40368 13268 40374 13280
rect 37568 13212 38148 13240
rect 38746 13200 38752 13252
rect 38804 13249 38810 13252
rect 38804 13243 38826 13249
rect 38814 13209 38826 13243
rect 38930 13240 38936 13252
rect 38891 13212 38936 13240
rect 38804 13203 38826 13209
rect 38804 13200 38810 13203
rect 38930 13200 38936 13212
rect 38988 13200 38994 13252
rect 40402 13240 40408 13252
rect 40363 13212 40408 13240
rect 40402 13200 40408 13212
rect 40460 13200 40466 13252
rect 37734 13172 37740 13184
rect 35084 13144 37740 13172
rect 37734 13132 37740 13144
rect 37792 13132 37798 13184
rect 37826 13132 37832 13184
rect 37884 13172 37890 13184
rect 38197 13175 38255 13181
rect 38197 13172 38209 13175
rect 37884 13144 38209 13172
rect 37884 13132 37890 13144
rect 38197 13141 38209 13144
rect 38243 13141 38255 13175
rect 38197 13135 38255 13141
rect 39666 13132 39672 13184
rect 39724 13172 39730 13184
rect 40037 13175 40095 13181
rect 40037 13172 40049 13175
rect 39724 13144 40049 13172
rect 39724 13132 39730 13144
rect 40037 13141 40049 13144
rect 40083 13141 40095 13175
rect 40037 13135 40095 13141
rect 40126 13132 40132 13184
rect 40184 13172 40190 13184
rect 40494 13172 40500 13184
rect 40184 13144 40500 13172
rect 40184 13132 40190 13144
rect 40494 13132 40500 13144
rect 40552 13132 40558 13184
rect 40604 13172 40632 13280
rect 40770 13268 40776 13320
rect 40828 13308 40834 13320
rect 40828 13280 40873 13308
rect 40828 13268 40834 13280
rect 40954 13268 40960 13320
rect 41012 13308 41018 13320
rect 41509 13311 41567 13317
rect 41012 13280 41368 13308
rect 41012 13268 41018 13280
rect 41046 13200 41052 13252
rect 41104 13240 41110 13252
rect 41233 13243 41291 13249
rect 41233 13240 41245 13243
rect 41104 13212 41245 13240
rect 41104 13200 41110 13212
rect 41233 13209 41245 13212
rect 41279 13209 41291 13243
rect 41340 13240 41368 13280
rect 41509 13277 41521 13311
rect 41555 13308 41567 13311
rect 41874 13308 41880 13320
rect 41555 13280 41880 13308
rect 41555 13277 41567 13280
rect 41509 13271 41567 13277
rect 41874 13268 41880 13280
rect 41932 13268 41938 13320
rect 42150 13308 42156 13320
rect 42111 13280 42156 13308
rect 42150 13268 42156 13280
rect 42208 13268 42214 13320
rect 42260 13317 42288 13348
rect 42794 13336 42800 13348
rect 42852 13336 42858 13388
rect 44100 13376 44128 13484
rect 44008 13348 44128 13376
rect 44008 13320 44036 13348
rect 42245 13311 42303 13317
rect 42245 13277 42257 13311
rect 42291 13277 42303 13311
rect 42426 13308 42432 13320
rect 42387 13280 42432 13308
rect 42245 13271 42303 13277
rect 42426 13268 42432 13280
rect 42484 13268 42490 13320
rect 42521 13311 42579 13317
rect 42521 13277 42533 13311
rect 42567 13308 42579 13311
rect 42981 13311 43039 13317
rect 42981 13308 42993 13311
rect 42567 13280 42993 13308
rect 42567 13277 42579 13280
rect 42521 13271 42579 13277
rect 42981 13277 42993 13280
rect 43027 13277 43039 13311
rect 42981 13271 43039 13277
rect 43165 13311 43223 13317
rect 43165 13277 43177 13311
rect 43211 13277 43223 13311
rect 43438 13308 43444 13320
rect 43399 13280 43444 13308
rect 43165 13271 43223 13277
rect 43180 13240 43208 13271
rect 43438 13268 43444 13280
rect 43496 13268 43502 13320
rect 43990 13308 43996 13320
rect 43951 13280 43996 13308
rect 43990 13268 43996 13280
rect 44048 13268 44054 13320
rect 44174 13308 44180 13320
rect 44135 13280 44180 13308
rect 44174 13268 44180 13280
rect 44232 13268 44238 13320
rect 41340 13212 43208 13240
rect 41233 13203 41291 13209
rect 42242 13172 42248 13184
rect 40604 13144 42248 13172
rect 42242 13132 42248 13144
rect 42300 13132 42306 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 25866 12968 25872 12980
rect 25827 12940 25872 12968
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 26037 12971 26095 12977
rect 26037 12937 26049 12971
rect 26083 12968 26095 12971
rect 26142 12968 26148 12980
rect 26083 12940 26148 12968
rect 26083 12937 26095 12940
rect 26037 12931 26095 12937
rect 26142 12928 26148 12940
rect 26200 12928 26206 12980
rect 28905 12971 28963 12977
rect 28905 12937 28917 12971
rect 28951 12968 28963 12971
rect 30466 12968 30472 12980
rect 28951 12940 30472 12968
rect 28951 12937 28963 12940
rect 28905 12931 28963 12937
rect 30466 12928 30472 12940
rect 30524 12968 30530 12980
rect 30524 12940 30696 12968
rect 30524 12928 30530 12940
rect 30668 12912 30696 12940
rect 33134 12928 33140 12980
rect 33192 12968 33198 12980
rect 33502 12968 33508 12980
rect 33192 12940 33508 12968
rect 33192 12928 33198 12940
rect 33502 12928 33508 12940
rect 33560 12968 33566 12980
rect 33873 12971 33931 12977
rect 33873 12968 33885 12971
rect 33560 12940 33885 12968
rect 33560 12928 33566 12940
rect 33873 12937 33885 12940
rect 33919 12968 33931 12971
rect 34517 12971 34575 12977
rect 34517 12968 34529 12971
rect 33919 12940 34529 12968
rect 33919 12937 33931 12940
rect 33873 12931 33931 12937
rect 34517 12937 34529 12940
rect 34563 12937 34575 12971
rect 34517 12931 34575 12937
rect 35342 12928 35348 12980
rect 35400 12968 35406 12980
rect 35437 12971 35495 12977
rect 35437 12968 35449 12971
rect 35400 12940 35449 12968
rect 35400 12928 35406 12940
rect 35437 12937 35449 12940
rect 35483 12937 35495 12971
rect 36630 12968 36636 12980
rect 36591 12940 36636 12968
rect 35437 12931 35495 12937
rect 36630 12928 36636 12940
rect 36688 12928 36694 12980
rect 38286 12968 38292 12980
rect 38247 12940 38292 12968
rect 38286 12928 38292 12940
rect 38344 12928 38350 12980
rect 38746 12968 38752 12980
rect 38626 12940 38752 12968
rect 26237 12903 26295 12909
rect 26237 12869 26249 12903
rect 26283 12900 26295 12903
rect 26418 12900 26424 12912
rect 26283 12872 26424 12900
rect 26283 12869 26295 12872
rect 26237 12863 26295 12869
rect 26418 12860 26424 12872
rect 26476 12860 26482 12912
rect 27246 12900 27252 12912
rect 27207 12872 27252 12900
rect 27246 12860 27252 12872
rect 27304 12860 27310 12912
rect 27522 12909 27528 12912
rect 27465 12903 27528 12909
rect 27465 12869 27477 12903
rect 27511 12869 27528 12903
rect 27465 12863 27528 12869
rect 27522 12860 27528 12863
rect 27580 12860 27586 12912
rect 29086 12900 29092 12912
rect 28920 12872 29092 12900
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12832 23719 12835
rect 23842 12832 23848 12844
rect 23707 12804 23848 12832
rect 23707 12801 23719 12804
rect 23661 12795 23719 12801
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 24302 12832 24308 12844
rect 24263 12804 24308 12832
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 28350 12832 28356 12844
rect 27632 12804 28356 12832
rect 27632 12705 27660 12804
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 28920 12841 28948 12872
rect 29086 12860 29092 12872
rect 29144 12900 29150 12912
rect 30558 12900 30564 12912
rect 29144 12872 30564 12900
rect 29144 12860 29150 12872
rect 30558 12860 30564 12872
rect 30616 12860 30622 12912
rect 30650 12860 30656 12912
rect 30708 12900 30714 12912
rect 30929 12903 30987 12909
rect 30929 12900 30941 12903
rect 30708 12872 30941 12900
rect 30708 12860 30714 12872
rect 30929 12869 30941 12872
rect 30975 12869 30987 12903
rect 31110 12900 31116 12912
rect 31071 12872 31116 12900
rect 30929 12863 30987 12869
rect 31110 12860 31116 12872
rect 31168 12860 31174 12912
rect 31294 12860 31300 12912
rect 31352 12900 31358 12912
rect 34790 12900 34796 12912
rect 31352 12872 34796 12900
rect 31352 12860 31358 12872
rect 28905 12835 28963 12841
rect 28905 12801 28917 12835
rect 28951 12801 28963 12835
rect 28905 12795 28963 12801
rect 28994 12792 29000 12844
rect 29052 12832 29058 12844
rect 29178 12832 29184 12844
rect 29052 12804 29184 12832
rect 29052 12792 29058 12804
rect 29178 12792 29184 12804
rect 29236 12832 29242 12844
rect 29917 12835 29975 12841
rect 29917 12832 29929 12835
rect 29236 12804 29929 12832
rect 29236 12792 29242 12804
rect 29917 12801 29929 12804
rect 29963 12801 29975 12835
rect 30742 12832 30748 12844
rect 30703 12804 30748 12832
rect 29917 12795 29975 12801
rect 30742 12792 30748 12804
rect 30800 12792 30806 12844
rect 31570 12832 31576 12844
rect 31531 12804 31576 12832
rect 31570 12792 31576 12804
rect 31628 12792 31634 12844
rect 32692 12841 32720 12872
rect 34790 12860 34796 12872
rect 34848 12860 34854 12912
rect 35894 12900 35900 12912
rect 35636 12872 35900 12900
rect 31757 12835 31815 12841
rect 31757 12801 31769 12835
rect 31803 12801 31815 12835
rect 31757 12795 31815 12801
rect 32677 12835 32735 12841
rect 32677 12801 32689 12835
rect 32723 12801 32735 12835
rect 32677 12795 32735 12801
rect 28445 12767 28503 12773
rect 28445 12733 28457 12767
rect 28491 12764 28503 12767
rect 28534 12764 28540 12776
rect 28491 12736 28540 12764
rect 28491 12733 28503 12736
rect 28445 12727 28503 12733
rect 28534 12724 28540 12736
rect 28592 12724 28598 12776
rect 29840 12767 29898 12773
rect 29840 12733 29852 12767
rect 29886 12764 29898 12767
rect 29886 12736 30052 12764
rect 29886 12733 29898 12736
rect 29840 12727 29898 12733
rect 30024 12708 30052 12736
rect 30190 12724 30196 12776
rect 30248 12764 30254 12776
rect 30285 12767 30343 12773
rect 30285 12764 30297 12767
rect 30248 12736 30297 12764
rect 30248 12724 30254 12736
rect 30285 12733 30297 12736
rect 30331 12733 30343 12767
rect 30285 12727 30343 12733
rect 30834 12724 30840 12776
rect 30892 12764 30898 12776
rect 31386 12764 31392 12776
rect 30892 12736 31392 12764
rect 30892 12724 30898 12736
rect 31386 12724 31392 12736
rect 31444 12764 31450 12776
rect 31772 12764 31800 12795
rect 32950 12792 32956 12844
rect 33008 12832 33014 12844
rect 33689 12835 33747 12841
rect 33689 12832 33701 12835
rect 33008 12804 33701 12832
rect 33008 12792 33014 12804
rect 33689 12801 33701 12804
rect 33735 12801 33747 12835
rect 34422 12832 34428 12844
rect 34383 12804 34428 12832
rect 33689 12795 33747 12801
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 34701 12835 34759 12841
rect 34701 12832 34713 12835
rect 34532 12804 34713 12832
rect 32582 12764 32588 12776
rect 31444 12736 31800 12764
rect 32543 12736 32588 12764
rect 31444 12724 31450 12736
rect 32582 12724 32588 12736
rect 32640 12724 32646 12776
rect 34532 12708 34560 12804
rect 34701 12801 34713 12804
rect 34747 12832 34759 12835
rect 35526 12832 35532 12844
rect 34747 12804 35532 12832
rect 34747 12801 34759 12804
rect 34701 12795 34759 12801
rect 35526 12792 35532 12804
rect 35584 12792 35590 12844
rect 35636 12841 35664 12872
rect 35894 12860 35900 12872
rect 35952 12900 35958 12912
rect 38626 12900 38654 12940
rect 38746 12928 38752 12940
rect 38804 12968 38810 12980
rect 40310 12968 40316 12980
rect 38804 12940 40316 12968
rect 38804 12928 38810 12940
rect 40310 12928 40316 12940
rect 40368 12928 40374 12980
rect 40494 12928 40500 12980
rect 40552 12968 40558 12980
rect 41785 12971 41843 12977
rect 41785 12968 41797 12971
rect 40552 12940 41797 12968
rect 40552 12928 40558 12940
rect 41785 12937 41797 12940
rect 41831 12968 41843 12971
rect 44450 12968 44456 12980
rect 41831 12940 44456 12968
rect 41831 12937 41843 12940
rect 41785 12931 41843 12937
rect 44450 12928 44456 12940
rect 44508 12928 44514 12980
rect 35952 12872 38654 12900
rect 35952 12860 35958 12872
rect 38930 12860 38936 12912
rect 38988 12900 38994 12912
rect 40862 12900 40868 12912
rect 38988 12872 39804 12900
rect 40823 12872 40868 12900
rect 38988 12860 38994 12872
rect 35621 12835 35679 12841
rect 35621 12801 35633 12835
rect 35667 12801 35679 12835
rect 35621 12795 35679 12801
rect 36170 12792 36176 12844
rect 36228 12832 36234 12844
rect 36541 12835 36599 12841
rect 36541 12832 36553 12835
rect 36228 12804 36553 12832
rect 36228 12792 36234 12804
rect 36541 12801 36553 12804
rect 36587 12801 36599 12835
rect 36541 12795 36599 12801
rect 36722 12792 36728 12844
rect 36780 12832 36786 12844
rect 36906 12832 36912 12844
rect 36780 12804 36912 12832
rect 36780 12792 36786 12804
rect 36906 12792 36912 12804
rect 36964 12792 36970 12844
rect 37645 12835 37703 12841
rect 37645 12801 37657 12835
rect 37691 12801 37703 12835
rect 37826 12832 37832 12844
rect 37787 12804 37832 12832
rect 37645 12795 37703 12801
rect 35897 12767 35955 12773
rect 35897 12733 35909 12767
rect 35943 12764 35955 12767
rect 36814 12764 36820 12776
rect 35943 12736 36820 12764
rect 35943 12733 35955 12736
rect 35897 12727 35955 12733
rect 36814 12724 36820 12736
rect 36872 12724 36878 12776
rect 37660 12764 37688 12795
rect 37826 12792 37832 12804
rect 37884 12792 37890 12844
rect 39408 12841 39436 12872
rect 39393 12835 39451 12841
rect 39393 12801 39405 12835
rect 39439 12801 39451 12835
rect 39666 12832 39672 12844
rect 39627 12804 39672 12832
rect 39393 12795 39451 12801
rect 39666 12792 39672 12804
rect 39724 12792 39730 12844
rect 39776 12832 39804 12872
rect 40862 12860 40868 12872
rect 40920 12860 40926 12912
rect 41138 12900 41144 12912
rect 41064 12872 41144 12900
rect 40954 12832 40960 12844
rect 39776 12804 40960 12832
rect 40954 12792 40960 12804
rect 41012 12792 41018 12844
rect 41064 12841 41092 12872
rect 41138 12860 41144 12872
rect 41196 12860 41202 12912
rect 41874 12860 41880 12912
rect 41932 12900 41938 12912
rect 42613 12903 42671 12909
rect 42613 12900 42625 12903
rect 41932 12872 42625 12900
rect 41932 12860 41938 12872
rect 42613 12869 42625 12872
rect 42659 12869 42671 12903
rect 42613 12863 42671 12869
rect 41049 12835 41107 12841
rect 41049 12801 41061 12835
rect 41095 12801 41107 12835
rect 41230 12832 41236 12844
rect 41143 12804 41236 12832
rect 41049 12795 41107 12801
rect 39209 12767 39267 12773
rect 39209 12764 39221 12767
rect 37660 12736 39221 12764
rect 39209 12733 39221 12736
rect 39255 12733 39267 12767
rect 39209 12727 39267 12733
rect 39485 12767 39543 12773
rect 39485 12733 39497 12767
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 39577 12767 39635 12773
rect 39577 12733 39589 12767
rect 39623 12764 39635 12767
rect 41064 12764 41092 12795
rect 41230 12792 41236 12804
rect 41288 12792 41294 12844
rect 41325 12835 41383 12841
rect 41325 12801 41337 12835
rect 41371 12832 41383 12835
rect 41506 12832 41512 12844
rect 41371 12804 41512 12832
rect 41371 12801 41383 12804
rect 41325 12795 41383 12801
rect 41506 12792 41512 12804
rect 41564 12792 41570 12844
rect 39623 12736 41092 12764
rect 39623 12733 39635 12736
rect 39577 12727 39635 12733
rect 27617 12699 27675 12705
rect 27617 12665 27629 12699
rect 27663 12665 27675 12699
rect 27617 12659 27675 12665
rect 30006 12656 30012 12708
rect 30064 12696 30070 12708
rect 32309 12699 32367 12705
rect 32309 12696 32321 12699
rect 30064 12668 32321 12696
rect 30064 12656 30070 12668
rect 32309 12665 32321 12668
rect 32355 12665 32367 12699
rect 32309 12659 32367 12665
rect 34514 12656 34520 12708
rect 34572 12656 34578 12708
rect 35802 12696 35808 12708
rect 35715 12668 35808 12696
rect 35802 12656 35808 12668
rect 35860 12696 35866 12708
rect 39500 12696 39528 12727
rect 41248 12696 41276 12792
rect 45002 12696 45008 12708
rect 35860 12668 38424 12696
rect 39500 12668 41276 12696
rect 41386 12668 45008 12696
rect 35860 12656 35866 12668
rect 24946 12628 24952 12640
rect 24907 12600 24952 12628
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 26053 12631 26111 12637
rect 26053 12597 26065 12631
rect 26099 12628 26111 12631
rect 26326 12628 26332 12640
rect 26099 12600 26332 12628
rect 26099 12597 26111 12600
rect 26053 12591 26111 12597
rect 26326 12588 26332 12600
rect 26384 12588 26390 12640
rect 27433 12631 27491 12637
rect 27433 12597 27445 12631
rect 27479 12628 27491 12631
rect 27890 12628 27896 12640
rect 27479 12600 27896 12628
rect 27479 12597 27491 12600
rect 27433 12591 27491 12597
rect 27890 12588 27896 12600
rect 27948 12588 27954 12640
rect 29641 12631 29699 12637
rect 29641 12597 29653 12631
rect 29687 12628 29699 12631
rect 29914 12628 29920 12640
rect 29687 12600 29920 12628
rect 29687 12597 29699 12600
rect 29641 12591 29699 12597
rect 29914 12588 29920 12600
rect 29972 12588 29978 12640
rect 31294 12588 31300 12640
rect 31352 12628 31358 12640
rect 31573 12631 31631 12637
rect 31573 12628 31585 12631
rect 31352 12600 31585 12628
rect 31352 12588 31358 12600
rect 31573 12597 31585 12600
rect 31619 12597 31631 12631
rect 34698 12628 34704 12640
rect 34659 12600 34704 12628
rect 31573 12591 31631 12597
rect 34698 12588 34704 12600
rect 34756 12588 34762 12640
rect 36630 12588 36636 12640
rect 36688 12628 36694 12640
rect 37645 12631 37703 12637
rect 37645 12628 37657 12631
rect 36688 12600 37657 12628
rect 36688 12588 36694 12600
rect 37645 12597 37657 12600
rect 37691 12597 37703 12631
rect 38396 12628 38424 12668
rect 41386 12628 41414 12668
rect 45002 12656 45008 12668
rect 45060 12656 45066 12708
rect 38396 12600 41414 12628
rect 37645 12591 37703 12597
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 28534 12424 28540 12436
rect 28495 12396 28540 12424
rect 28534 12384 28540 12396
rect 28592 12384 28598 12436
rect 28905 12427 28963 12433
rect 28905 12393 28917 12427
rect 28951 12424 28963 12427
rect 28994 12424 29000 12436
rect 28951 12396 29000 12424
rect 28951 12393 28963 12396
rect 28905 12387 28963 12393
rect 28994 12384 29000 12396
rect 29052 12384 29058 12436
rect 30006 12424 30012 12436
rect 29840 12396 30012 12424
rect 29840 12365 29868 12396
rect 30006 12384 30012 12396
rect 30064 12384 30070 12436
rect 30190 12424 30196 12436
rect 30151 12396 30196 12424
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 32582 12424 32588 12436
rect 32543 12396 32588 12424
rect 32582 12384 32588 12396
rect 32640 12384 32646 12436
rect 32766 12384 32772 12436
rect 32824 12424 32830 12436
rect 35621 12427 35679 12433
rect 32824 12396 35480 12424
rect 32824 12384 32830 12396
rect 26881 12359 26939 12365
rect 26881 12325 26893 12359
rect 26927 12356 26939 12359
rect 29825 12359 29883 12365
rect 26927 12328 27292 12356
rect 26927 12325 26939 12328
rect 26881 12319 26939 12325
rect 27264 12300 27292 12328
rect 29825 12325 29837 12359
rect 29871 12325 29883 12359
rect 32674 12356 32680 12368
rect 29825 12319 29883 12325
rect 29932 12328 32680 12356
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24912 12260 25053 12288
rect 24912 12248 24918 12260
rect 25041 12257 25053 12260
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 27246 12248 27252 12300
rect 27304 12288 27310 12300
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27304 12260 27813 12288
rect 27304 12248 27310 12260
rect 27801 12257 27813 12260
rect 27847 12257 27859 12291
rect 27801 12251 27859 12257
rect 27890 12248 27896 12300
rect 27948 12288 27954 12300
rect 28629 12291 28687 12297
rect 27948 12260 27993 12288
rect 27948 12248 27954 12260
rect 28629 12257 28641 12291
rect 28675 12288 28687 12291
rect 29086 12288 29092 12300
rect 28675 12260 29092 12288
rect 28675 12257 28687 12260
rect 28629 12251 28687 12257
rect 29086 12248 29092 12260
rect 29144 12248 29150 12300
rect 25222 12220 25228 12232
rect 25183 12192 25228 12220
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 25869 12223 25927 12229
rect 25869 12220 25881 12223
rect 25740 12192 25881 12220
rect 25740 12180 25746 12192
rect 25869 12189 25881 12192
rect 25915 12189 25927 12223
rect 26142 12220 26148 12232
rect 26103 12192 26148 12220
rect 25869 12183 25927 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 27706 12220 27712 12232
rect 27667 12192 27712 12220
rect 27706 12180 27712 12192
rect 27764 12180 27770 12232
rect 28350 12180 28356 12232
rect 28408 12220 28414 12232
rect 28537 12223 28595 12229
rect 28537 12220 28549 12223
rect 28408 12192 28549 12220
rect 28408 12180 28414 12192
rect 28537 12189 28549 12192
rect 28583 12189 28595 12223
rect 28537 12183 28595 12189
rect 28994 12180 29000 12232
rect 29052 12220 29058 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29052 12192 29745 12220
rect 29052 12180 29058 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 27430 12112 27436 12164
rect 27488 12152 27494 12164
rect 29932 12152 29960 12328
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 33134 12356 33140 12368
rect 32968 12328 33140 12356
rect 32030 12288 32036 12300
rect 30944 12260 32036 12288
rect 30009 12223 30067 12229
rect 30009 12189 30021 12223
rect 30055 12220 30067 12223
rect 30650 12220 30656 12232
rect 30055 12192 30656 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 30650 12180 30656 12192
rect 30708 12220 30714 12232
rect 30944 12229 30972 12260
rect 32030 12248 32036 12260
rect 32088 12248 32094 12300
rect 32968 12297 32996 12328
rect 33134 12316 33140 12328
rect 33192 12356 33198 12368
rect 35342 12356 35348 12368
rect 33192 12328 35348 12356
rect 33192 12316 33198 12328
rect 35342 12316 35348 12328
rect 35400 12316 35406 12368
rect 32861 12291 32919 12297
rect 32861 12288 32873 12291
rect 32324 12260 32873 12288
rect 30929 12223 30987 12229
rect 30929 12220 30941 12223
rect 30708 12192 30941 12220
rect 30708 12180 30714 12192
rect 30929 12189 30941 12192
rect 30975 12189 30987 12223
rect 31113 12223 31171 12229
rect 31113 12220 31125 12223
rect 30929 12183 30987 12189
rect 31036 12192 31125 12220
rect 27488 12124 29960 12152
rect 27488 12112 27494 12124
rect 30374 12112 30380 12164
rect 30432 12152 30438 12164
rect 31036 12152 31064 12192
rect 31113 12189 31125 12192
rect 31159 12189 31171 12223
rect 31205 12223 31263 12229
rect 31205 12210 31217 12223
rect 31251 12210 31263 12223
rect 31113 12183 31171 12189
rect 31202 12158 31208 12210
rect 31260 12158 31266 12210
rect 31294 12180 31300 12232
rect 31352 12220 31358 12232
rect 31352 12192 31397 12220
rect 31352 12180 31358 12192
rect 31478 12180 31484 12232
rect 31536 12220 31542 12232
rect 32324 12220 32352 12260
rect 32861 12257 32873 12260
rect 32907 12257 32919 12291
rect 32861 12251 32919 12257
rect 32953 12291 33011 12297
rect 32953 12257 32965 12291
rect 32999 12257 33011 12291
rect 32953 12251 33011 12257
rect 33502 12248 33508 12300
rect 33560 12288 33566 12300
rect 33965 12291 34023 12297
rect 33965 12288 33977 12291
rect 33560 12260 33977 12288
rect 33560 12248 33566 12260
rect 33965 12257 33977 12260
rect 34011 12257 34023 12291
rect 33965 12251 34023 12257
rect 34057 12291 34115 12297
rect 34057 12257 34069 12291
rect 34103 12288 34115 12291
rect 34422 12288 34428 12300
rect 34103 12260 34428 12288
rect 34103 12257 34115 12260
rect 34057 12251 34115 12257
rect 34422 12248 34428 12260
rect 34480 12288 34486 12300
rect 34790 12288 34796 12300
rect 34480 12260 34796 12288
rect 34480 12248 34486 12260
rect 34790 12248 34796 12260
rect 34848 12248 34854 12300
rect 35452 12288 35480 12396
rect 35621 12393 35633 12427
rect 35667 12393 35679 12427
rect 35621 12387 35679 12393
rect 35526 12316 35532 12368
rect 35584 12356 35590 12368
rect 35636 12356 35664 12387
rect 36722 12384 36728 12436
rect 36780 12424 36786 12436
rect 37001 12427 37059 12433
rect 37001 12424 37013 12427
rect 36780 12396 37013 12424
rect 36780 12384 36786 12396
rect 37001 12393 37013 12396
rect 37047 12424 37059 12427
rect 40770 12424 40776 12436
rect 37047 12396 40776 12424
rect 37047 12393 37059 12396
rect 37001 12387 37059 12393
rect 40770 12384 40776 12396
rect 40828 12424 40834 12436
rect 40865 12427 40923 12433
rect 40865 12424 40877 12427
rect 40828 12396 40877 12424
rect 40828 12384 40834 12396
rect 40865 12393 40877 12396
rect 40911 12393 40923 12427
rect 40865 12387 40923 12393
rect 41693 12427 41751 12433
rect 41693 12393 41705 12427
rect 41739 12424 41751 12427
rect 41874 12424 41880 12436
rect 41739 12396 41880 12424
rect 41739 12393 41751 12396
rect 41693 12387 41751 12393
rect 41874 12384 41880 12396
rect 41932 12384 41938 12436
rect 36357 12359 36415 12365
rect 36357 12356 36369 12359
rect 35584 12328 36369 12356
rect 35584 12316 35590 12328
rect 36357 12325 36369 12328
rect 36403 12356 36415 12359
rect 39114 12356 39120 12368
rect 36403 12328 39120 12356
rect 36403 12325 36415 12328
rect 36357 12319 36415 12325
rect 39114 12316 39120 12328
rect 39172 12316 39178 12368
rect 36541 12291 36599 12297
rect 36541 12288 36553 12291
rect 35452 12260 36553 12288
rect 32766 12220 32772 12232
rect 31536 12192 32352 12220
rect 32727 12192 32772 12220
rect 31536 12180 31542 12192
rect 32766 12180 32772 12192
rect 32824 12180 32830 12232
rect 33042 12180 33048 12232
rect 33100 12220 33106 12232
rect 33100 12192 33145 12220
rect 33100 12180 33106 12192
rect 33594 12180 33600 12232
rect 33652 12220 33658 12232
rect 33870 12220 33876 12232
rect 33652 12192 33876 12220
rect 33652 12180 33658 12192
rect 33870 12180 33876 12192
rect 33928 12180 33934 12232
rect 34149 12223 34207 12229
rect 34149 12189 34161 12223
rect 34195 12220 34207 12223
rect 34330 12220 34336 12232
rect 34195 12192 34336 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 34330 12180 34336 12192
rect 34388 12220 34394 12232
rect 34606 12220 34612 12232
rect 34388 12192 34612 12220
rect 34388 12180 34394 12192
rect 34606 12180 34612 12192
rect 34664 12180 34670 12232
rect 35452 12229 35480 12260
rect 36541 12257 36553 12260
rect 36587 12288 36599 12291
rect 36630 12288 36636 12300
rect 36587 12260 36636 12288
rect 36587 12257 36599 12260
rect 36541 12251 36599 12257
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 35437 12223 35495 12229
rect 35437 12189 35449 12223
rect 35483 12189 35495 12223
rect 35437 12183 35495 12189
rect 35529 12223 35587 12229
rect 35529 12189 35541 12223
rect 35575 12220 35587 12223
rect 36265 12223 36323 12229
rect 36265 12220 36277 12223
rect 35575 12192 36277 12220
rect 35575 12189 35587 12192
rect 35529 12183 35587 12189
rect 36265 12189 36277 12192
rect 36311 12189 36323 12223
rect 36265 12183 36323 12189
rect 37737 12223 37795 12229
rect 37737 12189 37749 12223
rect 37783 12220 37795 12223
rect 39206 12220 39212 12232
rect 37783 12192 39212 12220
rect 37783 12189 37795 12192
rect 37737 12183 37795 12189
rect 33502 12152 33508 12164
rect 30432 12124 31064 12152
rect 31404 12124 33508 12152
rect 30432 12112 30438 12124
rect 25409 12087 25467 12093
rect 25409 12053 25421 12087
rect 25455 12084 25467 12087
rect 25498 12084 25504 12096
rect 25455 12056 25504 12084
rect 25455 12053 25467 12056
rect 25409 12047 25467 12053
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 27338 12084 27344 12096
rect 27299 12056 27344 12084
rect 27338 12044 27344 12056
rect 27396 12044 27402 12096
rect 27522 12044 27528 12096
rect 27580 12084 27586 12096
rect 30926 12084 30932 12096
rect 27580 12056 30932 12084
rect 27580 12044 27586 12056
rect 30926 12044 30932 12056
rect 30984 12084 30990 12096
rect 31404 12084 31432 12124
rect 33502 12112 33508 12124
rect 33560 12152 33566 12164
rect 35544 12152 35572 12183
rect 39206 12180 39212 12192
rect 39264 12180 39270 12232
rect 33560 12124 35572 12152
rect 33560 12112 33566 12124
rect 30984 12056 31432 12084
rect 30984 12044 30990 12056
rect 31478 12044 31484 12096
rect 31536 12084 31542 12096
rect 31573 12087 31631 12093
rect 31573 12084 31585 12087
rect 31536 12056 31585 12084
rect 31536 12044 31542 12056
rect 31573 12053 31585 12056
rect 31619 12053 31631 12087
rect 31573 12047 31631 12053
rect 32030 12044 32036 12096
rect 32088 12084 32094 12096
rect 34238 12084 34244 12096
rect 32088 12056 34244 12084
rect 32088 12044 32094 12056
rect 34238 12044 34244 12056
rect 34296 12044 34302 12096
rect 34333 12087 34391 12093
rect 34333 12053 34345 12087
rect 34379 12084 34391 12087
rect 34422 12084 34428 12096
rect 34379 12056 34428 12084
rect 34379 12053 34391 12056
rect 34333 12047 34391 12053
rect 34422 12044 34428 12056
rect 34480 12044 34486 12096
rect 35802 12084 35808 12096
rect 35763 12056 35808 12084
rect 35802 12044 35808 12056
rect 35860 12044 35866 12096
rect 36538 12084 36544 12096
rect 36499 12056 36544 12084
rect 36538 12044 36544 12056
rect 36596 12044 36602 12096
rect 37182 12044 37188 12096
rect 37240 12084 37246 12096
rect 37645 12087 37703 12093
rect 37645 12084 37657 12087
rect 37240 12056 37657 12084
rect 37240 12044 37246 12056
rect 37645 12053 37657 12056
rect 37691 12053 37703 12087
rect 37645 12047 37703 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 25682 11880 25688 11892
rect 25643 11852 25688 11880
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 26142 11880 26148 11892
rect 26103 11852 26148 11880
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 27338 11840 27344 11892
rect 27396 11880 27402 11892
rect 27617 11883 27675 11889
rect 27617 11880 27629 11883
rect 27396 11852 27629 11880
rect 27396 11840 27402 11852
rect 27617 11849 27629 11852
rect 27663 11849 27675 11883
rect 28810 11880 28816 11892
rect 28771 11852 28816 11880
rect 27617 11843 27675 11849
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 30469 11883 30527 11889
rect 30469 11880 30481 11883
rect 30432 11852 30481 11880
rect 30432 11840 30438 11852
rect 30469 11849 30481 11852
rect 30515 11849 30527 11883
rect 30469 11843 30527 11849
rect 31113 11883 31171 11889
rect 31113 11849 31125 11883
rect 31159 11880 31171 11883
rect 31202 11880 31208 11892
rect 31159 11852 31208 11880
rect 31159 11849 31171 11852
rect 31113 11843 31171 11849
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 31386 11840 31392 11892
rect 31444 11880 31450 11892
rect 31481 11883 31539 11889
rect 31481 11880 31493 11883
rect 31444 11852 31493 11880
rect 31444 11840 31450 11852
rect 31481 11849 31493 11852
rect 31527 11849 31539 11883
rect 31481 11843 31539 11849
rect 32769 11883 32827 11889
rect 32769 11849 32781 11883
rect 32815 11880 32827 11883
rect 33134 11880 33140 11892
rect 32815 11852 33140 11880
rect 32815 11849 32827 11852
rect 32769 11843 32827 11849
rect 33134 11840 33140 11852
rect 33192 11840 33198 11892
rect 33502 11880 33508 11892
rect 33463 11852 33508 11880
rect 33502 11840 33508 11852
rect 33560 11840 33566 11892
rect 34238 11840 34244 11892
rect 34296 11880 34302 11892
rect 34296 11852 35572 11880
rect 34296 11840 34302 11852
rect 35544 11824 35572 11852
rect 29086 11812 29092 11824
rect 26206 11784 27844 11812
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 1903 11716 2421 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2409 11713 2421 11716
rect 2455 11744 2467 11747
rect 18598 11744 18604 11756
rect 2455 11716 18604 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 25498 11744 25504 11756
rect 25459 11716 25504 11744
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 26206 11688 26234 11784
rect 26329 11747 26387 11753
rect 26329 11713 26341 11747
rect 26375 11744 26387 11747
rect 27522 11744 27528 11756
rect 26375 11716 27200 11744
rect 27483 11716 27528 11744
rect 26375 11713 26387 11716
rect 26329 11707 26387 11713
rect 25041 11679 25099 11685
rect 25041 11645 25053 11679
rect 25087 11676 25099 11679
rect 25222 11676 25228 11688
rect 25087 11648 25228 11676
rect 25087 11645 25099 11648
rect 25041 11639 25099 11645
rect 25222 11636 25228 11648
rect 25280 11676 25286 11688
rect 26206 11676 26240 11688
rect 25280 11648 26240 11676
rect 25280 11636 25286 11648
rect 26234 11636 26240 11648
rect 26292 11636 26298 11688
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 27172 11617 27200 11716
rect 27522 11704 27528 11716
rect 27580 11704 27586 11756
rect 27816 11685 27844 11784
rect 28552 11784 29092 11812
rect 27801 11679 27859 11685
rect 27801 11645 27813 11679
rect 27847 11676 27859 11679
rect 28552 11676 28580 11784
rect 29086 11772 29092 11784
rect 29144 11772 29150 11824
rect 30006 11772 30012 11824
rect 30064 11812 30070 11824
rect 32585 11815 32643 11821
rect 32585 11812 32597 11815
rect 30064 11784 32597 11812
rect 30064 11772 30070 11784
rect 32585 11781 32597 11784
rect 32631 11812 32643 11815
rect 33042 11812 33048 11824
rect 32631 11784 33048 11812
rect 32631 11781 32643 11784
rect 32585 11775 32643 11781
rect 33042 11772 33048 11784
rect 33100 11812 33106 11824
rect 34422 11812 34428 11824
rect 33100 11784 33364 11812
rect 34383 11784 34428 11812
rect 33100 11772 33106 11784
rect 28994 11744 29000 11756
rect 28955 11716 29000 11744
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 30466 11744 30472 11756
rect 30427 11716 30472 11744
rect 30466 11704 30472 11716
rect 30524 11704 30530 11756
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11744 30711 11747
rect 31110 11744 31116 11756
rect 30699 11716 31116 11744
rect 30699 11713 30711 11716
rect 30653 11707 30711 11713
rect 31110 11704 31116 11716
rect 31168 11704 31174 11756
rect 31297 11747 31355 11753
rect 31297 11713 31309 11747
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 29178 11676 29184 11688
rect 27847 11648 28580 11676
rect 29139 11648 29184 11676
rect 27847 11645 27859 11648
rect 27801 11639 27859 11645
rect 29178 11636 29184 11648
rect 29236 11636 29242 11688
rect 30484 11676 30512 11704
rect 31312 11676 31340 11707
rect 31570 11704 31576 11756
rect 31628 11744 31634 11756
rect 31628 11716 31673 11744
rect 31628 11704 31634 11716
rect 32766 11704 32772 11756
rect 32824 11744 32830 11756
rect 33336 11753 33364 11784
rect 34422 11772 34428 11784
rect 34480 11772 34486 11824
rect 34609 11815 34667 11821
rect 34609 11781 34621 11815
rect 34655 11812 34667 11815
rect 34698 11812 34704 11824
rect 34655 11784 34704 11812
rect 34655 11781 34667 11784
rect 34609 11775 34667 11781
rect 34698 11772 34704 11784
rect 34756 11772 34762 11824
rect 35526 11812 35532 11824
rect 35439 11784 35532 11812
rect 35526 11772 35532 11784
rect 35584 11772 35590 11824
rect 35802 11821 35808 11824
rect 35745 11815 35808 11821
rect 35745 11781 35757 11815
rect 35791 11781 35808 11815
rect 35745 11775 35808 11781
rect 35802 11772 35808 11775
rect 35860 11772 35866 11824
rect 40586 11812 40592 11824
rect 36372 11784 38056 11812
rect 32861 11747 32919 11753
rect 32861 11744 32873 11747
rect 32824 11716 32873 11744
rect 32824 11704 32830 11716
rect 32861 11713 32873 11716
rect 32907 11713 32919 11747
rect 32861 11707 32919 11713
rect 33321 11747 33379 11753
rect 33321 11713 33333 11747
rect 33367 11713 33379 11747
rect 36262 11744 36268 11756
rect 33321 11707 33379 11713
rect 33428 11716 36268 11744
rect 30484 11648 31340 11676
rect 27157 11611 27215 11617
rect 27157 11577 27169 11611
rect 27203 11577 27215 11611
rect 27157 11571 27215 11577
rect 30009 11611 30067 11617
rect 30009 11577 30021 11611
rect 30055 11608 30067 11611
rect 30650 11608 30656 11620
rect 30055 11580 30656 11608
rect 30055 11577 30067 11580
rect 30009 11571 30067 11577
rect 30650 11568 30656 11580
rect 30708 11568 30714 11620
rect 31588 11608 31616 11704
rect 32674 11636 32680 11688
rect 32732 11676 32738 11688
rect 33428 11676 33456 11716
rect 36262 11704 36268 11716
rect 36320 11704 36326 11756
rect 36372 11676 36400 11784
rect 36722 11744 36728 11756
rect 36683 11716 36728 11744
rect 36722 11704 36728 11716
rect 36780 11704 36786 11756
rect 36906 11704 36912 11756
rect 36964 11744 36970 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36964 11716 37841 11744
rect 36964 11704 36970 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 38028 11685 38056 11784
rect 38488 11784 40592 11812
rect 38194 11744 38200 11756
rect 38155 11716 38200 11744
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 38488 11753 38516 11784
rect 40586 11772 40592 11784
rect 40644 11772 40650 11824
rect 38473 11747 38531 11753
rect 38473 11713 38485 11747
rect 38519 11713 38531 11747
rect 38473 11707 38531 11713
rect 38841 11747 38899 11753
rect 38841 11713 38853 11747
rect 38887 11744 38899 11747
rect 39206 11744 39212 11756
rect 38887 11716 39212 11744
rect 38887 11713 38899 11716
rect 38841 11707 38899 11713
rect 32732 11648 33456 11676
rect 34624 11648 36400 11676
rect 36633 11679 36691 11685
rect 32732 11636 32738 11648
rect 32585 11611 32643 11617
rect 32585 11608 32597 11611
rect 31588 11580 32597 11608
rect 32585 11577 32597 11580
rect 32631 11577 32643 11611
rect 32585 11571 32643 11577
rect 28442 11500 28448 11552
rect 28500 11540 28506 11552
rect 34624 11540 34652 11648
rect 36633 11645 36645 11679
rect 36679 11645 36691 11679
rect 36633 11639 36691 11645
rect 38013 11679 38071 11685
rect 38013 11645 38025 11679
rect 38059 11645 38071 11679
rect 38013 11639 38071 11645
rect 36538 11608 36544 11620
rect 35728 11580 36544 11608
rect 34790 11540 34796 11552
rect 28500 11512 34652 11540
rect 34751 11512 34796 11540
rect 28500 11500 28506 11512
rect 34790 11500 34796 11512
rect 34848 11500 34854 11552
rect 35728 11549 35756 11580
rect 36538 11568 36544 11580
rect 36596 11568 36602 11620
rect 36648 11608 36676 11639
rect 38488 11608 38516 11707
rect 39206 11704 39212 11716
rect 39264 11704 39270 11756
rect 39298 11704 39304 11756
rect 39356 11744 39362 11756
rect 39356 11716 39401 11744
rect 39356 11704 39362 11716
rect 36648 11580 38516 11608
rect 35713 11543 35771 11549
rect 35713 11509 35725 11543
rect 35759 11509 35771 11543
rect 35894 11540 35900 11552
rect 35855 11512 35900 11540
rect 35713 11503 35771 11509
rect 35894 11500 35900 11512
rect 35952 11500 35958 11552
rect 36354 11540 36360 11552
rect 36315 11512 36360 11540
rect 36354 11500 36360 11512
rect 36412 11500 36418 11552
rect 39114 11500 39120 11552
rect 39172 11540 39178 11552
rect 39393 11543 39451 11549
rect 39393 11540 39405 11543
rect 39172 11512 39405 11540
rect 39172 11500 39178 11512
rect 39393 11509 39405 11512
rect 39439 11509 39451 11543
rect 39758 11540 39764 11552
rect 39719 11512 39764 11540
rect 39393 11503 39451 11509
rect 39758 11500 39764 11512
rect 39816 11500 39822 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25685 11339 25743 11345
rect 25685 11336 25697 11339
rect 24912 11308 25697 11336
rect 24912 11296 24918 11308
rect 25685 11305 25697 11308
rect 25731 11336 25743 11339
rect 27430 11336 27436 11348
rect 25731 11308 26924 11336
rect 27391 11308 27436 11336
rect 25731 11305 25743 11308
rect 25685 11299 25743 11305
rect 26234 11228 26240 11280
rect 26292 11268 26298 11280
rect 26292 11240 26337 11268
rect 26292 11228 26298 11240
rect 26896 11073 26924 11308
rect 27430 11296 27436 11308
rect 27488 11296 27494 11348
rect 29270 11296 29276 11348
rect 29328 11336 29334 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 29328 11308 29929 11336
rect 29328 11296 29334 11308
rect 29917 11305 29929 11308
rect 29963 11305 29975 11339
rect 29917 11299 29975 11305
rect 30469 11339 30527 11345
rect 30469 11305 30481 11339
rect 30515 11336 30527 11339
rect 30558 11336 30564 11348
rect 30515 11308 30564 11336
rect 30515 11305 30527 11308
rect 30469 11299 30527 11305
rect 30558 11296 30564 11308
rect 30616 11296 30622 11348
rect 32953 11339 33011 11345
rect 32953 11305 32965 11339
rect 32999 11336 33011 11339
rect 33226 11336 33232 11348
rect 32999 11308 33232 11336
rect 32999 11305 33011 11308
rect 32953 11299 33011 11305
rect 33226 11296 33232 11308
rect 33284 11296 33290 11348
rect 33870 11296 33876 11348
rect 33928 11336 33934 11348
rect 34977 11339 35035 11345
rect 34977 11336 34989 11339
rect 33928 11308 34989 11336
rect 33928 11296 33934 11308
rect 34977 11305 34989 11308
rect 35023 11305 35035 11339
rect 34977 11299 35035 11305
rect 35526 11296 35532 11348
rect 35584 11336 35590 11348
rect 36173 11339 36231 11345
rect 36173 11336 36185 11339
rect 35584 11308 36185 11336
rect 35584 11296 35590 11308
rect 36173 11305 36185 11308
rect 36219 11336 36231 11339
rect 36219 11308 36492 11336
rect 36219 11305 36231 11308
rect 36173 11299 36231 11305
rect 28994 11268 29000 11280
rect 28552 11240 29000 11268
rect 28552 11209 28580 11240
rect 28994 11228 29000 11240
rect 29052 11268 29058 11280
rect 36354 11268 36360 11280
rect 29052 11240 36360 11268
rect 29052 11228 29058 11240
rect 36354 11228 36360 11240
rect 36412 11228 36418 11280
rect 36464 11268 36492 11308
rect 36722 11296 36728 11348
rect 36780 11336 36786 11348
rect 36817 11339 36875 11345
rect 36817 11336 36829 11339
rect 36780 11308 36829 11336
rect 36780 11296 36786 11308
rect 36817 11305 36829 11308
rect 36863 11305 36875 11339
rect 36817 11299 36875 11305
rect 36998 11296 37004 11348
rect 37056 11336 37062 11348
rect 37734 11336 37740 11348
rect 37056 11308 37740 11336
rect 37056 11296 37062 11308
rect 37734 11296 37740 11308
rect 37792 11336 37798 11348
rect 38194 11336 38200 11348
rect 37792 11308 38200 11336
rect 37792 11296 37798 11308
rect 38194 11296 38200 11308
rect 38252 11296 38258 11348
rect 58158 11336 58164 11348
rect 58119 11308 58164 11336
rect 58158 11296 58164 11308
rect 58216 11296 58222 11348
rect 39117 11271 39175 11277
rect 39117 11268 39129 11271
rect 36464 11240 39129 11268
rect 39117 11237 39129 11240
rect 39163 11268 39175 11271
rect 39298 11268 39304 11280
rect 39163 11240 39304 11268
rect 39163 11237 39175 11240
rect 39117 11231 39175 11237
rect 39298 11228 39304 11240
rect 39356 11228 39362 11280
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11169 28595 11203
rect 29178 11200 29184 11212
rect 28537 11163 28595 11169
rect 28644 11172 29184 11200
rect 28644 11141 28672 11172
rect 29178 11160 29184 11172
rect 29236 11200 29242 11212
rect 32306 11200 32312 11212
rect 29236 11172 32312 11200
rect 29236 11160 29242 11172
rect 32306 11160 32312 11172
rect 32364 11160 32370 11212
rect 32401 11203 32459 11209
rect 32401 11169 32413 11203
rect 32447 11200 32459 11203
rect 33226 11200 33232 11212
rect 32447 11172 33232 11200
rect 32447 11169 32459 11172
rect 32401 11163 32459 11169
rect 33226 11160 33232 11172
rect 33284 11160 33290 11212
rect 33873 11203 33931 11209
rect 33873 11169 33885 11203
rect 33919 11200 33931 11203
rect 33962 11200 33968 11212
rect 33919 11172 33968 11200
rect 33919 11169 33931 11172
rect 33873 11163 33931 11169
rect 33962 11160 33968 11172
rect 34020 11160 34026 11212
rect 36998 11200 37004 11212
rect 36959 11172 37004 11200
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 37093 11203 37151 11209
rect 37093 11169 37105 11203
rect 37139 11200 37151 11203
rect 37366 11200 37372 11212
rect 37139 11172 37372 11200
rect 37139 11169 37151 11172
rect 37093 11163 37151 11169
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11101 28687 11135
rect 29730 11132 29736 11144
rect 28629 11095 28687 11101
rect 29012 11104 29736 11132
rect 26881 11067 26939 11073
rect 26881 11033 26893 11067
rect 26927 11064 26939 11067
rect 26927 11036 28028 11064
rect 26927 11033 26939 11036
rect 26881 11027 26939 11033
rect 28000 11005 28028 11036
rect 27985 10999 28043 11005
rect 27985 10965 27997 10999
rect 28031 10996 28043 10999
rect 28718 10996 28724 11008
rect 28031 10968 28724 10996
rect 28031 10965 28043 10968
rect 27985 10959 28043 10965
rect 28718 10956 28724 10968
rect 28776 10956 28782 11008
rect 29012 11005 29040 11104
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 29914 11132 29920 11144
rect 29875 11104 29920 11132
rect 29914 11092 29920 11104
rect 29972 11092 29978 11144
rect 32125 11135 32183 11141
rect 32125 11101 32137 11135
rect 32171 11101 32183 11135
rect 32125 11095 32183 11101
rect 32217 11135 32275 11141
rect 32217 11101 32229 11135
rect 32263 11132 32275 11135
rect 33502 11132 33508 11144
rect 32263 11104 33508 11132
rect 32263 11101 32275 11104
rect 32217 11095 32275 11101
rect 32140 11064 32168 11095
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 33597 11135 33655 11141
rect 33597 11101 33609 11135
rect 33643 11101 33655 11135
rect 33597 11095 33655 11101
rect 33042 11064 33048 11076
rect 32140 11036 33048 11064
rect 33042 11024 33048 11036
rect 33100 11064 33106 11076
rect 33612 11064 33640 11095
rect 33686 11092 33692 11144
rect 33744 11132 33750 11144
rect 33744 11104 33789 11132
rect 33744 11092 33750 11104
rect 34422 11092 34428 11144
rect 34480 11132 34486 11144
rect 35069 11135 35127 11141
rect 35069 11132 35081 11135
rect 34480 11104 35081 11132
rect 34480 11092 34486 11104
rect 35069 11101 35081 11104
rect 35115 11132 35127 11135
rect 35529 11135 35587 11141
rect 35529 11132 35541 11135
rect 35115 11104 35541 11132
rect 35115 11101 35127 11104
rect 35069 11095 35127 11101
rect 35529 11101 35541 11104
rect 35575 11101 35587 11135
rect 35710 11132 35716 11144
rect 35671 11104 35716 11132
rect 35529 11095 35587 11101
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 36446 11092 36452 11144
rect 36504 11132 36510 11144
rect 36906 11132 36912 11144
rect 36504 11104 36912 11132
rect 36504 11092 36510 11104
rect 36906 11092 36912 11104
rect 36964 11132 36970 11144
rect 37185 11135 37243 11141
rect 37185 11132 37197 11135
rect 36964 11104 37197 11132
rect 36964 11092 36970 11104
rect 37185 11101 37197 11104
rect 37231 11101 37243 11135
rect 37185 11095 37243 11101
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37829 11135 37887 11141
rect 37829 11132 37841 11135
rect 37332 11104 37841 11132
rect 37332 11092 37338 11104
rect 37829 11101 37841 11104
rect 37875 11101 37887 11135
rect 37829 11095 37887 11101
rect 33870 11064 33876 11076
rect 33100 11036 33640 11064
rect 33831 11036 33876 11064
rect 33100 11024 33106 11036
rect 33870 11024 33876 11036
rect 33928 11024 33934 11076
rect 35621 11067 35679 11073
rect 35621 11033 35633 11067
rect 35667 11064 35679 11067
rect 38562 11064 38568 11076
rect 35667 11036 38568 11064
rect 35667 11033 35679 11036
rect 35621 11027 35679 11033
rect 38562 11024 38568 11036
rect 38620 11024 38626 11076
rect 57609 11067 57667 11073
rect 57609 11033 57621 11067
rect 57655 11064 57667 11067
rect 58250 11064 58256 11076
rect 57655 11036 58256 11064
rect 57655 11033 57667 11036
rect 57609 11027 57667 11033
rect 58250 11024 58256 11036
rect 58308 11024 58314 11076
rect 28997 10999 29055 11005
rect 28997 10965 29009 10999
rect 29043 10965 29055 10999
rect 28997 10959 29055 10965
rect 32401 10999 32459 11005
rect 32401 10965 32413 10999
rect 32447 10996 32459 10999
rect 32490 10996 32496 11008
rect 32447 10968 32496 10996
rect 32447 10965 32459 10968
rect 32401 10959 32459 10965
rect 32490 10956 32496 10968
rect 32548 10956 32554 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 28905 10795 28963 10801
rect 28905 10761 28917 10795
rect 28951 10761 28963 10795
rect 32306 10792 32312 10804
rect 32267 10764 32312 10792
rect 28905 10755 28963 10761
rect 27433 10727 27491 10733
rect 27433 10693 27445 10727
rect 27479 10724 27491 10727
rect 27706 10724 27712 10736
rect 27479 10696 27712 10724
rect 27479 10693 27491 10696
rect 27433 10687 27491 10693
rect 27706 10684 27712 10696
rect 27764 10684 27770 10736
rect 28718 10724 28724 10736
rect 28658 10696 28724 10724
rect 28718 10684 28724 10696
rect 28776 10684 28782 10736
rect 28920 10724 28948 10755
rect 32306 10752 32312 10764
rect 32364 10752 32370 10804
rect 32477 10795 32535 10801
rect 32477 10761 32489 10795
rect 32523 10792 32535 10795
rect 33137 10795 33195 10801
rect 33137 10792 33149 10795
rect 32523 10764 33149 10792
rect 32523 10761 32535 10764
rect 32477 10755 32535 10761
rect 33137 10761 33149 10764
rect 33183 10761 33195 10795
rect 33137 10755 33195 10761
rect 33686 10752 33692 10804
rect 33744 10792 33750 10804
rect 35437 10795 35495 10801
rect 35437 10792 35449 10795
rect 33744 10764 35449 10792
rect 33744 10752 33750 10764
rect 35437 10761 35449 10764
rect 35483 10761 35495 10795
rect 37274 10792 37280 10804
rect 35437 10755 35495 10761
rect 36280 10764 37280 10792
rect 36280 10736 36308 10764
rect 37274 10752 37280 10764
rect 37332 10792 37338 10804
rect 37461 10795 37519 10801
rect 37461 10792 37473 10795
rect 37332 10764 37473 10792
rect 37332 10752 37338 10764
rect 37461 10761 37473 10764
rect 37507 10761 37519 10795
rect 37461 10755 37519 10761
rect 30006 10724 30012 10736
rect 28920 10696 30012 10724
rect 30006 10684 30012 10696
rect 30064 10684 30070 10736
rect 31018 10684 31024 10736
rect 31076 10684 31082 10736
rect 31294 10684 31300 10736
rect 31352 10724 31358 10736
rect 32677 10727 32735 10733
rect 32677 10724 32689 10727
rect 31352 10696 32689 10724
rect 31352 10684 31358 10696
rect 32677 10693 32689 10696
rect 32723 10724 32735 10727
rect 34422 10724 34428 10736
rect 32723 10696 34428 10724
rect 32723 10693 32735 10696
rect 32677 10687 32735 10693
rect 34422 10684 34428 10696
rect 34480 10684 34486 10736
rect 34698 10684 34704 10736
rect 34756 10724 34762 10736
rect 35710 10724 35716 10736
rect 34756 10696 35716 10724
rect 34756 10684 34762 10696
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27120 10628 27169 10656
rect 27120 10616 27126 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 31757 10659 31815 10665
rect 31757 10625 31769 10659
rect 31803 10656 31815 10659
rect 33042 10656 33048 10668
rect 31803 10628 33048 10656
rect 31803 10625 31815 10628
rect 31757 10619 31815 10625
rect 33042 10616 33048 10628
rect 33100 10656 33106 10668
rect 33321 10659 33379 10665
rect 33321 10656 33333 10659
rect 33100 10628 33333 10656
rect 33100 10616 33106 10628
rect 33321 10625 33333 10628
rect 33367 10625 33379 10659
rect 33502 10656 33508 10668
rect 33463 10628 33508 10656
rect 33321 10619 33379 10625
rect 33502 10616 33508 10628
rect 33560 10656 33566 10668
rect 33560 10628 34468 10656
rect 33560 10616 33566 10628
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 34440 10597 34468 10628
rect 34606 10616 34612 10668
rect 34664 10656 34670 10668
rect 35544 10665 35572 10696
rect 35710 10684 35716 10696
rect 35768 10684 35774 10736
rect 36262 10724 36268 10736
rect 36223 10696 36268 10724
rect 36262 10684 36268 10696
rect 36320 10684 36326 10736
rect 36446 10724 36452 10736
rect 36407 10696 36452 10724
rect 36446 10684 36452 10696
rect 36504 10684 36510 10736
rect 39485 10727 39543 10733
rect 39485 10693 39497 10727
rect 39531 10724 39543 10727
rect 39758 10724 39764 10736
rect 39531 10696 39764 10724
rect 39531 10693 39543 10696
rect 39485 10687 39543 10693
rect 39758 10684 39764 10696
rect 39816 10684 39822 10736
rect 35345 10659 35403 10665
rect 35345 10656 35357 10659
rect 34664 10628 35357 10656
rect 34664 10616 34670 10628
rect 35345 10625 35357 10628
rect 35391 10625 35403 10659
rect 35345 10619 35403 10625
rect 35529 10659 35587 10665
rect 35529 10625 35541 10659
rect 35575 10625 35587 10659
rect 35529 10619 35587 10625
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29144 10560 29745 10588
rect 29144 10548 29150 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 34425 10591 34483 10597
rect 34425 10557 34437 10591
rect 34471 10557 34483 10591
rect 34698 10588 34704 10600
rect 34659 10560 34704 10588
rect 34425 10551 34483 10557
rect 34698 10548 34704 10560
rect 34756 10548 34762 10600
rect 34793 10591 34851 10597
rect 34793 10557 34805 10591
rect 34839 10557 34851 10591
rect 34793 10551 34851 10557
rect 33962 10480 33968 10532
rect 34020 10520 34026 10532
rect 34808 10520 34836 10551
rect 39114 10520 39120 10532
rect 34020 10492 34836 10520
rect 39075 10492 39120 10520
rect 34020 10480 34026 10492
rect 39114 10480 39120 10492
rect 39172 10480 39178 10532
rect 26418 10452 26424 10464
rect 26379 10424 26424 10452
rect 26418 10412 26424 10424
rect 26476 10412 26482 10464
rect 32490 10452 32496 10464
rect 32451 10424 32496 10452
rect 32490 10412 32496 10424
rect 32548 10412 32554 10464
rect 33226 10412 33232 10464
rect 33284 10452 33290 10464
rect 33321 10455 33379 10461
rect 33321 10452 33333 10455
rect 33284 10424 33333 10452
rect 33284 10412 33290 10424
rect 33321 10421 33333 10424
rect 33367 10421 33379 10455
rect 36078 10452 36084 10464
rect 36039 10424 36084 10452
rect 33321 10415 33379 10421
rect 36078 10412 36084 10424
rect 36136 10412 36142 10464
rect 38286 10412 38292 10464
rect 38344 10452 38350 10464
rect 39025 10455 39083 10461
rect 39025 10452 39037 10455
rect 38344 10424 39037 10452
rect 38344 10412 38350 10424
rect 39025 10421 39037 10424
rect 39071 10421 39083 10455
rect 39025 10415 39083 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 26881 10251 26939 10257
rect 26881 10217 26893 10251
rect 26927 10248 26939 10251
rect 27062 10248 27068 10260
rect 26927 10220 27068 10248
rect 26927 10217 26939 10220
rect 26881 10211 26939 10217
rect 27062 10208 27068 10220
rect 27120 10248 27126 10260
rect 29086 10248 29092 10260
rect 27120 10220 29092 10248
rect 27120 10208 27126 10220
rect 29086 10208 29092 10220
rect 29144 10208 29150 10260
rect 30282 10248 30288 10260
rect 29840 10220 30288 10248
rect 27433 10183 27491 10189
rect 27433 10149 27445 10183
rect 27479 10180 27491 10183
rect 29840 10180 29868 10220
rect 30282 10208 30288 10220
rect 30340 10248 30346 10260
rect 31297 10251 31355 10257
rect 31297 10248 31309 10251
rect 30340 10220 31309 10248
rect 30340 10208 30346 10220
rect 31297 10217 31309 10220
rect 31343 10248 31355 10251
rect 32490 10248 32496 10260
rect 31343 10220 32496 10248
rect 31343 10217 31355 10220
rect 31297 10211 31355 10217
rect 32490 10208 32496 10220
rect 32548 10208 32554 10260
rect 33226 10248 33232 10260
rect 33187 10220 33232 10248
rect 33226 10208 33232 10220
rect 33284 10208 33290 10260
rect 33686 10208 33692 10260
rect 33744 10248 33750 10260
rect 33873 10251 33931 10257
rect 33873 10248 33885 10251
rect 33744 10220 33885 10248
rect 33744 10208 33750 10220
rect 33873 10217 33885 10220
rect 33919 10217 33931 10251
rect 33873 10211 33931 10217
rect 27479 10152 29868 10180
rect 27479 10149 27491 10152
rect 27433 10143 27491 10149
rect 27908 10053 27936 10152
rect 29914 10140 29920 10192
rect 29972 10140 29978 10192
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 36817 10183 36875 10189
rect 36817 10180 36829 10183
rect 34572 10152 36829 10180
rect 34572 10140 34578 10152
rect 36817 10149 36829 10152
rect 36863 10149 36875 10183
rect 36817 10143 36875 10149
rect 29825 10115 29883 10121
rect 29825 10081 29837 10115
rect 29871 10112 29883 10115
rect 29932 10112 29960 10140
rect 29871 10084 29960 10112
rect 30285 10115 30343 10121
rect 29871 10081 29883 10084
rect 29825 10075 29883 10081
rect 30285 10081 30297 10115
rect 30331 10112 30343 10115
rect 31018 10112 31024 10124
rect 30331 10084 31024 10112
rect 30331 10081 30343 10084
rect 30285 10075 30343 10081
rect 31018 10072 31024 10084
rect 31076 10072 31082 10124
rect 36078 10112 36084 10124
rect 36039 10084 36084 10112
rect 36078 10072 36084 10084
rect 36136 10072 36142 10124
rect 37277 10115 37335 10121
rect 37277 10081 37289 10115
rect 37323 10112 37335 10115
rect 37458 10112 37464 10124
rect 37323 10084 37464 10112
rect 37323 10081 37335 10084
rect 37277 10075 37335 10081
rect 37458 10072 37464 10084
rect 37516 10072 37522 10124
rect 39114 10072 39120 10124
rect 39172 10112 39178 10124
rect 40129 10115 40187 10121
rect 40129 10112 40141 10115
rect 39172 10084 40141 10112
rect 39172 10072 39178 10084
rect 40129 10081 40141 10084
rect 40175 10081 40187 10115
rect 40129 10075 40187 10081
rect 27893 10047 27951 10053
rect 27893 10013 27905 10047
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 28077 10047 28135 10053
rect 28077 10013 28089 10047
rect 28123 10044 28135 10047
rect 28902 10044 28908 10056
rect 28123 10016 28908 10044
rect 28123 10013 28135 10016
rect 28077 10007 28135 10013
rect 28902 10004 28908 10016
rect 28960 10004 28966 10056
rect 29730 10004 29736 10056
rect 29788 10044 29794 10056
rect 29917 10047 29975 10053
rect 29917 10044 29929 10047
rect 29788 10016 29929 10044
rect 29788 10004 29794 10016
rect 29917 10013 29929 10016
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 31205 10047 31263 10053
rect 31205 10013 31217 10047
rect 31251 10044 31263 10047
rect 31294 10044 31300 10056
rect 31251 10016 31300 10044
rect 31251 10013 31263 10016
rect 31205 10007 31263 10013
rect 31294 10004 31300 10016
rect 31352 10004 31358 10056
rect 33042 10004 33048 10056
rect 33100 10044 33106 10056
rect 33873 10047 33931 10053
rect 33873 10044 33885 10047
rect 33100 10016 33885 10044
rect 33100 10004 33106 10016
rect 33873 10013 33885 10016
rect 33919 10013 33931 10047
rect 33873 10007 33931 10013
rect 33962 10004 33968 10056
rect 34020 10044 34026 10056
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 34020 10016 34069 10044
rect 34020 10004 34026 10016
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34057 10007 34115 10013
rect 35989 10047 36047 10053
rect 35989 10013 36001 10047
rect 36035 10013 36047 10047
rect 37182 10044 37188 10056
rect 37143 10016 37188 10044
rect 35989 10007 36047 10013
rect 36004 9976 36032 10007
rect 37182 10004 37188 10016
rect 37240 10004 37246 10056
rect 38286 10044 38292 10056
rect 38247 10016 38292 10044
rect 38286 10004 38292 10016
rect 38344 10004 38350 10056
rect 38562 10044 38568 10056
rect 38523 10016 38568 10044
rect 38562 10004 38568 10016
rect 38620 10004 38626 10056
rect 38749 10047 38807 10053
rect 38749 10013 38761 10047
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 37734 9976 37740 9988
rect 36004 9948 37740 9976
rect 37734 9936 37740 9948
rect 37792 9936 37798 9988
rect 38378 9936 38384 9988
rect 38436 9976 38442 9988
rect 38764 9976 38792 10007
rect 39758 10004 39764 10056
rect 39816 10044 39822 10056
rect 40221 10047 40279 10053
rect 40221 10044 40233 10047
rect 39816 10016 40233 10044
rect 39816 10004 39822 10016
rect 40221 10013 40233 10016
rect 40267 10013 40279 10047
rect 40221 10007 40279 10013
rect 38436 9948 38792 9976
rect 38436 9936 38442 9948
rect 27890 9908 27896 9920
rect 27851 9880 27896 9908
rect 27890 9868 27896 9880
rect 27948 9868 27954 9920
rect 28629 9911 28687 9917
rect 28629 9877 28641 9911
rect 28675 9908 28687 9911
rect 28718 9908 28724 9920
rect 28675 9880 28724 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 28718 9868 28724 9880
rect 28776 9868 28782 9920
rect 33686 9908 33692 9920
rect 33647 9880 33692 9908
rect 33686 9868 33692 9880
rect 33744 9868 33750 9920
rect 35621 9911 35679 9917
rect 35621 9877 35633 9911
rect 35667 9908 35679 9911
rect 35710 9908 35716 9920
rect 35667 9880 35716 9908
rect 35667 9877 35679 9880
rect 35621 9871 35679 9877
rect 35710 9868 35716 9880
rect 35768 9868 35774 9920
rect 37642 9868 37648 9920
rect 37700 9908 37706 9920
rect 38105 9911 38163 9917
rect 38105 9908 38117 9911
rect 37700 9880 38117 9908
rect 37700 9868 37706 9880
rect 38105 9877 38117 9880
rect 38151 9877 38163 9911
rect 38105 9871 38163 9877
rect 40589 9911 40647 9917
rect 40589 9877 40601 9911
rect 40635 9908 40647 9911
rect 57514 9908 57520 9920
rect 40635 9880 57520 9908
rect 40635 9877 40647 9880
rect 40589 9871 40647 9877
rect 57514 9868 57520 9880
rect 57572 9868 57578 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 28902 9704 28908 9716
rect 28863 9676 28908 9704
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 36906 9664 36912 9716
rect 36964 9704 36970 9716
rect 38378 9704 38384 9716
rect 36964 9676 38384 9704
rect 36964 9664 36970 9676
rect 28718 9636 28724 9648
rect 28658 9608 28724 9636
rect 28718 9596 28724 9608
rect 28776 9596 28782 9648
rect 28920 9636 28948 9664
rect 29641 9639 29699 9645
rect 29641 9636 29653 9639
rect 28920 9608 29653 9636
rect 29641 9605 29653 9608
rect 29687 9605 29699 9639
rect 29641 9599 29699 9605
rect 29825 9639 29883 9645
rect 29825 9605 29837 9639
rect 29871 9636 29883 9639
rect 30374 9636 30380 9648
rect 29871 9608 30380 9636
rect 29871 9605 29883 9608
rect 29825 9599 29883 9605
rect 30374 9596 30380 9608
rect 30432 9636 30438 9648
rect 31294 9636 31300 9648
rect 30432 9608 31300 9636
rect 30432 9596 30438 9608
rect 31294 9596 31300 9608
rect 31352 9596 31358 9648
rect 32490 9636 32496 9648
rect 32451 9608 32496 9636
rect 32490 9596 32496 9608
rect 32548 9636 32554 9648
rect 33042 9636 33048 9648
rect 32548 9608 33048 9636
rect 32548 9596 32554 9608
rect 33042 9596 33048 9608
rect 33100 9636 33106 9648
rect 37660 9645 37688 9676
rect 38378 9664 38384 9676
rect 38436 9664 38442 9716
rect 37645 9639 37703 9645
rect 33100 9608 34008 9636
rect 33100 9596 33106 9608
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9568 26663 9571
rect 27062 9568 27068 9580
rect 26651 9540 27068 9568
rect 26651 9537 26663 9540
rect 26605 9531 26663 9537
rect 27062 9528 27068 9540
rect 27120 9568 27126 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 27120 9540 27169 9568
rect 27120 9528 27126 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 31018 9568 31024 9580
rect 30979 9540 31024 9568
rect 27157 9531 27215 9537
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 33686 9568 33692 9580
rect 33647 9540 33692 9568
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 33870 9568 33876 9580
rect 33831 9540 33876 9568
rect 33870 9528 33876 9540
rect 33928 9528 33934 9580
rect 33980 9577 34008 9608
rect 35084 9608 35756 9636
rect 33965 9571 34023 9577
rect 33965 9537 33977 9571
rect 34011 9537 34023 9571
rect 33965 9531 34023 9537
rect 34425 9571 34483 9577
rect 34425 9537 34437 9571
rect 34471 9568 34483 9571
rect 34514 9568 34520 9580
rect 34471 9540 34520 9568
rect 34471 9537 34483 9540
rect 34425 9531 34483 9537
rect 34514 9528 34520 9540
rect 34572 9528 34578 9580
rect 34790 9528 34796 9580
rect 34848 9568 34854 9580
rect 35084 9577 35112 9608
rect 35728 9580 35756 9608
rect 37645 9605 37657 9639
rect 37691 9605 37703 9639
rect 37645 9599 37703 9605
rect 34885 9571 34943 9577
rect 34885 9568 34897 9571
rect 34848 9540 34897 9568
rect 34848 9528 34854 9540
rect 34885 9537 34897 9540
rect 34931 9537 34943 9571
rect 34885 9531 34943 9537
rect 35069 9571 35127 9577
rect 35069 9537 35081 9571
rect 35115 9537 35127 9571
rect 35526 9568 35532 9580
rect 35069 9531 35127 9537
rect 35176 9540 35532 9568
rect 27430 9500 27436 9512
rect 27391 9472 27436 9500
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 30558 9500 30564 9512
rect 30471 9472 30564 9500
rect 30558 9460 30564 9472
rect 30616 9500 30622 9512
rect 30926 9500 30932 9512
rect 30616 9472 30932 9500
rect 30616 9460 30622 9472
rect 30926 9460 30932 9472
rect 30984 9460 30990 9512
rect 31113 9503 31171 9509
rect 31113 9469 31125 9503
rect 31159 9500 31171 9503
rect 31202 9500 31208 9512
rect 31159 9472 31208 9500
rect 31159 9469 31171 9472
rect 31113 9463 31171 9469
rect 31202 9460 31208 9472
rect 31260 9460 31266 9512
rect 34900 9500 34928 9531
rect 35176 9500 35204 9540
rect 35526 9528 35532 9540
rect 35584 9528 35590 9580
rect 35710 9568 35716 9580
rect 35671 9540 35716 9568
rect 35710 9528 35716 9540
rect 35768 9528 35774 9580
rect 36909 9571 36967 9577
rect 36909 9537 36921 9571
rect 36955 9568 36967 9571
rect 37274 9568 37280 9580
rect 36955 9540 37280 9568
rect 36955 9537 36967 9540
rect 36909 9531 36967 9537
rect 37274 9528 37280 9540
rect 37332 9568 37338 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 37332 9540 37473 9568
rect 37332 9528 37338 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37734 9568 37740 9580
rect 37695 9540 37740 9568
rect 37461 9531 37519 9537
rect 37734 9528 37740 9540
rect 37792 9528 37798 9580
rect 38396 9568 38424 9664
rect 38565 9571 38623 9577
rect 38565 9568 38577 9571
rect 38396 9540 38577 9568
rect 38565 9537 38577 9540
rect 38611 9537 38623 9571
rect 38565 9531 38623 9537
rect 38470 9500 38476 9512
rect 34900 9472 35204 9500
rect 38431 9472 38476 9500
rect 38470 9460 38476 9472
rect 38528 9460 38534 9512
rect 38933 9503 38991 9509
rect 38933 9469 38945 9503
rect 38979 9500 38991 9503
rect 39114 9500 39120 9512
rect 38979 9472 39120 9500
rect 38979 9469 38991 9472
rect 38933 9463 38991 9469
rect 39114 9460 39120 9472
rect 39172 9460 39178 9512
rect 32950 9392 32956 9444
rect 33008 9432 33014 9444
rect 34333 9435 34391 9441
rect 34333 9432 34345 9435
rect 33008 9404 34345 9432
rect 33008 9392 33014 9404
rect 34333 9401 34345 9404
rect 34379 9401 34391 9435
rect 37458 9432 37464 9444
rect 37419 9404 37464 9432
rect 34333 9395 34391 9401
rect 37458 9392 37464 9404
rect 37516 9392 37522 9444
rect 30006 9364 30012 9376
rect 29967 9336 30012 9364
rect 30006 9324 30012 9336
rect 30064 9324 30070 9376
rect 31110 9364 31116 9376
rect 31071 9336 31116 9364
rect 31110 9324 31116 9336
rect 31168 9324 31174 9376
rect 31386 9364 31392 9376
rect 31347 9336 31392 9364
rect 31386 9324 31392 9336
rect 31444 9324 31450 9376
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 35069 9367 35127 9373
rect 35069 9364 35081 9367
rect 34848 9336 35081 9364
rect 34848 9324 34854 9336
rect 35069 9333 35081 9336
rect 35115 9333 35127 9367
rect 35618 9364 35624 9376
rect 35579 9336 35624 9364
rect 35069 9327 35127 9333
rect 35618 9324 35624 9336
rect 35676 9324 35682 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 27157 9163 27215 9169
rect 27157 9129 27169 9163
rect 27203 9160 27215 9163
rect 27430 9160 27436 9172
rect 27203 9132 27436 9160
rect 27203 9129 27215 9132
rect 27157 9123 27215 9129
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 28166 9120 28172 9172
rect 28224 9160 28230 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 28224 9132 28273 9160
rect 28224 9120 28230 9132
rect 28261 9129 28273 9132
rect 28307 9160 28319 9163
rect 28718 9160 28724 9172
rect 28307 9132 28724 9160
rect 28307 9129 28319 9132
rect 28261 9123 28319 9129
rect 28718 9120 28724 9132
rect 28776 9160 28782 9172
rect 29089 9163 29147 9169
rect 29089 9160 29101 9163
rect 28776 9132 29101 9160
rect 28776 9120 28782 9132
rect 29089 9129 29101 9132
rect 29135 9160 29147 9163
rect 30558 9160 30564 9172
rect 29135 9132 30564 9160
rect 29135 9129 29147 9132
rect 29089 9123 29147 9129
rect 30558 9120 30564 9132
rect 30616 9120 30622 9172
rect 30837 9163 30895 9169
rect 30837 9129 30849 9163
rect 30883 9160 30895 9163
rect 31110 9160 31116 9172
rect 30883 9132 31116 9160
rect 30883 9129 30895 9132
rect 30837 9123 30895 9129
rect 31110 9120 31116 9132
rect 31168 9160 31174 9172
rect 31389 9163 31447 9169
rect 31389 9160 31401 9163
rect 31168 9132 31401 9160
rect 31168 9120 31174 9132
rect 31389 9129 31401 9132
rect 31435 9129 31447 9163
rect 32950 9160 32956 9172
rect 32911 9132 32956 9160
rect 31389 9123 31447 9129
rect 32950 9120 32956 9132
rect 33008 9120 33014 9172
rect 29825 9095 29883 9101
rect 29825 9061 29837 9095
rect 29871 9092 29883 9095
rect 30650 9092 30656 9104
rect 29871 9064 30656 9092
rect 29871 9061 29883 9064
rect 29825 9055 29883 9061
rect 30650 9052 30656 9064
rect 30708 9052 30714 9104
rect 34241 9095 34299 9101
rect 34241 9092 34253 9095
rect 31496 9064 34253 9092
rect 31018 9024 31024 9036
rect 30668 8996 31024 9024
rect 26418 8916 26424 8968
rect 26476 8956 26482 8968
rect 26605 8959 26663 8965
rect 26605 8956 26617 8959
rect 26476 8928 26617 8956
rect 26476 8916 26482 8928
rect 26605 8925 26617 8928
rect 26651 8956 26663 8959
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 26651 8928 27077 8956
rect 26651 8925 26663 8928
rect 26605 8919 26663 8925
rect 27065 8925 27077 8928
rect 27111 8956 27123 8959
rect 27154 8956 27160 8968
rect 27111 8928 27160 8956
rect 27111 8925 27123 8928
rect 27065 8919 27123 8925
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8956 27307 8959
rect 27890 8956 27896 8968
rect 27295 8928 27896 8956
rect 27295 8925 27307 8928
rect 27249 8919 27307 8925
rect 27890 8916 27896 8928
rect 27948 8916 27954 8968
rect 30006 8956 30012 8968
rect 29967 8928 30012 8956
rect 30006 8916 30012 8928
rect 30064 8916 30070 8968
rect 30668 8965 30696 8996
rect 31018 8984 31024 8996
rect 31076 8984 31082 9036
rect 30653 8959 30711 8965
rect 30653 8925 30665 8959
rect 30699 8925 30711 8959
rect 30653 8919 30711 8925
rect 30929 8959 30987 8965
rect 30929 8925 30941 8959
rect 30975 8956 30987 8959
rect 31202 8956 31208 8968
rect 30975 8928 31208 8956
rect 30975 8925 30987 8928
rect 30929 8919 30987 8925
rect 31202 8916 31208 8928
rect 31260 8956 31266 8968
rect 31496 8956 31524 9064
rect 31573 9027 31631 9033
rect 31573 8993 31585 9027
rect 31619 9024 31631 9027
rect 32766 9024 32772 9036
rect 31619 8996 32772 9024
rect 31619 8993 31631 8996
rect 31573 8987 31631 8993
rect 32766 8984 32772 8996
rect 32824 8984 32830 9036
rect 32876 9033 32904 9064
rect 34241 9061 34253 9064
rect 34287 9061 34299 9095
rect 34241 9055 34299 9061
rect 32861 9027 32919 9033
rect 32861 8993 32873 9027
rect 32907 9024 32919 9027
rect 32950 9024 32956 9036
rect 32907 8996 32956 9024
rect 32907 8993 32919 8996
rect 32861 8987 32919 8993
rect 32950 8984 32956 8996
rect 33008 8984 33014 9036
rect 33686 8984 33692 9036
rect 33744 9024 33750 9036
rect 35621 9027 35679 9033
rect 33744 8996 34008 9024
rect 33744 8984 33750 8996
rect 31665 8959 31723 8965
rect 31665 8956 31677 8959
rect 31260 8928 31677 8956
rect 31260 8916 31266 8928
rect 31665 8925 31677 8928
rect 31711 8925 31723 8959
rect 31665 8919 31723 8925
rect 31757 8959 31815 8965
rect 31757 8925 31769 8959
rect 31803 8956 31815 8959
rect 32585 8959 32643 8965
rect 32585 8956 32597 8959
rect 31803 8928 32597 8956
rect 31803 8925 31815 8928
rect 31757 8919 31815 8925
rect 32585 8925 32597 8928
rect 32631 8925 32643 8959
rect 33870 8956 33876 8968
rect 33831 8928 33876 8956
rect 32585 8919 32643 8925
rect 27338 8848 27344 8900
rect 27396 8888 27402 8900
rect 27985 8891 28043 8897
rect 27985 8888 27997 8891
rect 27396 8860 27997 8888
rect 27396 8848 27402 8860
rect 27985 8857 27997 8860
rect 28031 8857 28043 8891
rect 27985 8851 28043 8857
rect 31478 8848 31484 8900
rect 31536 8888 31542 8900
rect 31772 8888 31800 8919
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 33980 8965 34008 8996
rect 35621 8993 35633 9027
rect 35667 9024 35679 9027
rect 35710 9024 35716 9036
rect 35667 8996 35716 9024
rect 35667 8993 35679 8996
rect 35621 8987 35679 8993
rect 35710 8984 35716 8996
rect 35768 8984 35774 9036
rect 33965 8959 34023 8965
rect 33965 8925 33977 8959
rect 34011 8925 34023 8959
rect 33965 8919 34023 8925
rect 34057 8959 34115 8965
rect 34057 8925 34069 8959
rect 34103 8956 34115 8959
rect 34514 8956 34520 8968
rect 34103 8928 34520 8956
rect 34103 8925 34115 8928
rect 34057 8919 34115 8925
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 35526 8956 35532 8968
rect 35487 8928 35532 8956
rect 35526 8916 35532 8928
rect 35584 8916 35590 8968
rect 37642 8956 37648 8968
rect 37603 8928 37648 8956
rect 37642 8916 37648 8928
rect 37700 8916 37706 8968
rect 37826 8916 37832 8968
rect 37884 8956 37890 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 37884 8928 38025 8956
rect 37884 8916 37890 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 31536 8860 31800 8888
rect 31536 8848 31542 8860
rect 33042 8848 33048 8900
rect 33100 8888 33106 8900
rect 33689 8891 33747 8897
rect 33689 8888 33701 8891
rect 33100 8860 33701 8888
rect 33100 8848 33106 8860
rect 33689 8857 33701 8860
rect 33735 8857 33747 8891
rect 33689 8851 33747 8857
rect 39485 8891 39543 8897
rect 39485 8857 39497 8891
rect 39531 8888 39543 8891
rect 57698 8888 57704 8900
rect 39531 8860 57704 8888
rect 39531 8857 39543 8860
rect 39485 8851 39543 8857
rect 57698 8848 57704 8860
rect 57756 8848 57762 8900
rect 30466 8820 30472 8832
rect 30427 8792 30472 8820
rect 30466 8780 30472 8792
rect 30524 8780 30530 8832
rect 33137 8823 33195 8829
rect 33137 8789 33149 8823
rect 33183 8820 33195 8823
rect 33870 8820 33876 8832
rect 33183 8792 33876 8820
rect 33183 8789 33195 8792
rect 33137 8783 33195 8789
rect 33870 8780 33876 8792
rect 33928 8780 33934 8832
rect 35897 8823 35955 8829
rect 35897 8789 35909 8823
rect 35943 8820 35955 8823
rect 36078 8820 36084 8832
rect 35943 8792 36084 8820
rect 35943 8789 35955 8792
rect 35897 8783 35955 8789
rect 36078 8780 36084 8792
rect 36136 8780 36142 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 27120 8588 27905 8616
rect 27120 8576 27126 8588
rect 27893 8585 27905 8588
rect 27939 8585 27951 8619
rect 27893 8579 27951 8585
rect 30193 8619 30251 8625
rect 30193 8585 30205 8619
rect 30239 8616 30251 8619
rect 30374 8616 30380 8628
rect 30239 8588 30380 8616
rect 30239 8585 30251 8588
rect 30193 8579 30251 8585
rect 27908 8480 27936 8579
rect 30374 8576 30380 8588
rect 30432 8576 30438 8628
rect 31113 8619 31171 8625
rect 31113 8585 31125 8619
rect 31159 8616 31171 8619
rect 31386 8616 31392 8628
rect 31159 8588 31392 8616
rect 31159 8585 31171 8588
rect 31113 8579 31171 8585
rect 31386 8576 31392 8588
rect 31444 8576 31450 8628
rect 32677 8619 32735 8625
rect 32677 8585 32689 8619
rect 32723 8616 32735 8619
rect 33781 8619 33839 8625
rect 33781 8616 33793 8619
rect 32723 8588 33793 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 33781 8585 33793 8588
rect 33827 8616 33839 8619
rect 34054 8616 34060 8628
rect 33827 8588 34060 8616
rect 33827 8585 33839 8588
rect 33781 8579 33839 8585
rect 34054 8576 34060 8588
rect 34112 8576 34118 8628
rect 35069 8619 35127 8625
rect 35069 8585 35081 8619
rect 35115 8616 35127 8619
rect 35618 8616 35624 8628
rect 35115 8588 35624 8616
rect 35115 8585 35127 8588
rect 35069 8579 35127 8585
rect 35618 8576 35624 8588
rect 35676 8576 35682 8628
rect 30558 8548 30564 8560
rect 29946 8520 30564 8548
rect 30558 8508 30564 8520
rect 30616 8508 30622 8560
rect 32858 8548 32864 8560
rect 32784 8520 32864 8548
rect 28445 8483 28503 8489
rect 28445 8480 28457 8483
rect 27908 8452 28457 8480
rect 28445 8449 28457 8452
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 30466 8440 30472 8492
rect 30524 8480 30530 8492
rect 30929 8483 30987 8489
rect 30929 8480 30941 8483
rect 30524 8452 30941 8480
rect 30524 8440 30530 8452
rect 30929 8449 30941 8452
rect 30975 8480 30987 8483
rect 31018 8480 31024 8492
rect 30975 8452 31024 8480
rect 30975 8449 30987 8452
rect 30929 8443 30987 8449
rect 31018 8440 31024 8452
rect 31076 8440 31082 8492
rect 31202 8480 31208 8492
rect 31163 8452 31208 8480
rect 31202 8440 31208 8452
rect 31260 8440 31266 8492
rect 31478 8440 31484 8492
rect 31536 8480 31542 8492
rect 32784 8489 32812 8520
rect 32858 8508 32864 8520
rect 32916 8508 32922 8560
rect 37642 8508 37648 8560
rect 37700 8548 37706 8560
rect 38013 8551 38071 8557
rect 38013 8548 38025 8551
rect 37700 8520 38025 8548
rect 37700 8508 37706 8520
rect 38013 8517 38025 8520
rect 38059 8517 38071 8551
rect 38013 8511 38071 8517
rect 32493 8483 32551 8489
rect 32493 8480 32505 8483
rect 31536 8452 32505 8480
rect 31536 8440 31542 8452
rect 32493 8449 32505 8452
rect 32539 8449 32551 8483
rect 32493 8443 32551 8449
rect 32769 8483 32827 8489
rect 32769 8449 32781 8483
rect 32815 8449 32827 8483
rect 32950 8480 32956 8492
rect 32911 8452 32956 8480
rect 32769 8443 32827 8449
rect 32950 8440 32956 8452
rect 33008 8440 33014 8492
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 27154 8372 27160 8424
rect 27212 8412 27218 8424
rect 28721 8415 28779 8421
rect 28721 8412 28733 8415
rect 27212 8384 28733 8412
rect 27212 8372 27218 8384
rect 28721 8381 28733 8384
rect 28767 8412 28779 8415
rect 28767 8384 29776 8412
rect 28767 8381 28779 8384
rect 28721 8375 28779 8381
rect 27338 8344 27344 8356
rect 27299 8316 27344 8344
rect 27338 8304 27344 8316
rect 27396 8304 27402 8356
rect 29748 8344 29776 8384
rect 30098 8372 30104 8424
rect 30156 8412 30162 8424
rect 30745 8415 30803 8421
rect 30745 8412 30757 8415
rect 30156 8384 30757 8412
rect 30156 8372 30162 8384
rect 30745 8381 30757 8384
rect 30791 8381 30803 8415
rect 33612 8412 33640 8443
rect 33870 8440 33876 8492
rect 33928 8480 33934 8492
rect 33928 8452 33973 8480
rect 33928 8440 33934 8452
rect 34790 8440 34796 8492
rect 34848 8480 34854 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34848 8452 34897 8480
rect 34848 8440 34854 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 35161 8483 35219 8489
rect 35161 8449 35173 8483
rect 35207 8480 35219 8483
rect 35894 8480 35900 8492
rect 35207 8452 35900 8480
rect 35207 8449 35219 8452
rect 35161 8443 35219 8449
rect 35894 8440 35900 8452
rect 35952 8440 35958 8492
rect 36078 8480 36084 8492
rect 36039 8452 36084 8480
rect 36078 8440 36084 8452
rect 36136 8440 36142 8492
rect 33962 8412 33968 8424
rect 33612 8384 33968 8412
rect 30745 8375 30803 8381
rect 33962 8372 33968 8384
rect 34020 8412 34026 8424
rect 34701 8415 34759 8421
rect 34701 8412 34713 8415
rect 34020 8384 34713 8412
rect 34020 8372 34026 8384
rect 34701 8381 34713 8384
rect 34747 8381 34759 8415
rect 34701 8375 34759 8381
rect 36909 8415 36967 8421
rect 36909 8381 36921 8415
rect 36955 8381 36967 8415
rect 36909 8375 36967 8381
rect 30650 8344 30656 8356
rect 29748 8316 30656 8344
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 36924 8344 36952 8375
rect 37737 8347 37795 8353
rect 37737 8344 37749 8347
rect 36924 8316 37749 8344
rect 37737 8313 37749 8316
rect 37783 8344 37795 8347
rect 37826 8344 37832 8356
rect 37783 8316 37832 8344
rect 37783 8313 37795 8316
rect 37737 8307 37795 8313
rect 37826 8304 37832 8316
rect 37884 8304 37890 8356
rect 33226 8236 33232 8288
rect 33284 8276 33290 8288
rect 33413 8279 33471 8285
rect 33413 8276 33425 8279
rect 33284 8248 33425 8276
rect 33284 8236 33290 8248
rect 33413 8245 33425 8248
rect 33459 8245 33471 8279
rect 37550 8276 37556 8288
rect 37511 8248 37556 8276
rect 33413 8239 33471 8245
rect 37550 8236 37556 8248
rect 37608 8236 37614 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 28166 8072 28172 8084
rect 28127 8044 28172 8072
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30650 8072 30656 8084
rect 30423 8044 30656 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30650 8032 30656 8044
rect 30708 8032 30714 8084
rect 33870 8032 33876 8084
rect 33928 8072 33934 8084
rect 33965 8075 34023 8081
rect 33965 8072 33977 8075
rect 33928 8044 33977 8072
rect 33928 8032 33934 8044
rect 33965 8041 33977 8044
rect 34011 8041 34023 8075
rect 33965 8035 34023 8041
rect 31386 8004 31392 8016
rect 31347 7976 31392 8004
rect 31386 7964 31392 7976
rect 31444 7964 31450 8016
rect 31018 7936 31024 7948
rect 30979 7908 31024 7936
rect 31018 7896 31024 7908
rect 31076 7896 31082 7948
rect 31202 7828 31208 7880
rect 31260 7868 31266 7880
rect 32861 7871 32919 7877
rect 32861 7868 32873 7871
rect 31260 7840 32873 7868
rect 31260 7828 31266 7840
rect 32861 7837 32873 7840
rect 32907 7837 32919 7871
rect 32861 7831 32919 7837
rect 33045 7871 33103 7877
rect 33045 7837 33057 7871
rect 33091 7837 33103 7871
rect 33226 7868 33232 7880
rect 33187 7840 33232 7868
rect 33045 7831 33103 7837
rect 33060 7800 33088 7831
rect 33226 7828 33232 7840
rect 33284 7828 33290 7880
rect 33321 7871 33379 7877
rect 33321 7837 33333 7871
rect 33367 7868 33379 7871
rect 33778 7868 33784 7880
rect 33367 7840 33784 7868
rect 33367 7837 33379 7840
rect 33321 7831 33379 7837
rect 33778 7828 33784 7840
rect 33836 7868 33842 7880
rect 37550 7868 37556 7880
rect 33836 7840 37556 7868
rect 33836 7828 33842 7840
rect 37550 7828 37556 7840
rect 37608 7828 37614 7880
rect 33134 7800 33140 7812
rect 33047 7772 33140 7800
rect 33134 7760 33140 7772
rect 33192 7800 33198 7812
rect 33962 7809 33968 7812
rect 33949 7803 33968 7809
rect 33192 7772 33824 7800
rect 33192 7760 33198 7772
rect 31386 7692 31392 7744
rect 31444 7732 31450 7744
rect 33796 7741 33824 7772
rect 33949 7769 33961 7803
rect 33949 7763 33968 7769
rect 33962 7760 33968 7763
rect 34020 7760 34026 7812
rect 34054 7760 34060 7812
rect 34112 7800 34118 7812
rect 34149 7803 34207 7809
rect 34149 7800 34161 7803
rect 34112 7772 34161 7800
rect 34112 7760 34118 7772
rect 34149 7769 34161 7772
rect 34195 7769 34207 7803
rect 34149 7763 34207 7769
rect 31481 7735 31539 7741
rect 31481 7732 31493 7735
rect 31444 7704 31493 7732
rect 31444 7692 31450 7704
rect 31481 7701 31493 7704
rect 31527 7701 31539 7735
rect 31481 7695 31539 7701
rect 33781 7735 33839 7741
rect 33781 7701 33793 7735
rect 33827 7701 33839 7735
rect 33781 7695 33839 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 31386 7392 31392 7404
rect 31347 7364 31392 7392
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 33686 7392 33692 7404
rect 33647 7364 33692 7392
rect 33686 7352 33692 7364
rect 33744 7352 33750 7404
rect 31202 7284 31208 7336
rect 31260 7324 31266 7336
rect 31297 7327 31355 7333
rect 31297 7324 31309 7327
rect 31260 7296 31309 7324
rect 31260 7284 31266 7296
rect 31297 7293 31309 7296
rect 31343 7293 31355 7327
rect 33778 7324 33784 7336
rect 33739 7296 33784 7324
rect 31297 7287 31355 7293
rect 33778 7284 33784 7296
rect 33836 7284 33842 7336
rect 33321 7259 33379 7265
rect 33321 7256 33333 7259
rect 26206 7228 33333 7256
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 26206 7188 26234 7228
rect 33321 7225 33333 7228
rect 33367 7225 33379 7259
rect 33321 7219 33379 7225
rect 22336 7160 26234 7188
rect 31757 7191 31815 7197
rect 22336 7148 22342 7160
rect 31757 7157 31769 7191
rect 31803 7188 31815 7191
rect 32950 7188 32956 7200
rect 31803 7160 32956 7188
rect 31803 7157 31815 7160
rect 31757 7151 31815 7157
rect 32950 7148 32956 7160
rect 33008 7148 33014 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 33686 6984 33692 6996
rect 33647 6956 33692 6984
rect 33686 6944 33692 6956
rect 33744 6944 33750 6996
rect 24946 6876 24952 6928
rect 25004 6916 25010 6928
rect 27706 6916 27712 6928
rect 25004 6888 27712 6916
rect 25004 6876 25010 6888
rect 27706 6876 27712 6888
rect 27764 6876 27770 6928
rect 33226 6876 33232 6928
rect 33284 6916 33290 6928
rect 33505 6919 33563 6925
rect 33505 6916 33517 6919
rect 33284 6888 33517 6916
rect 33284 6876 33290 6888
rect 33505 6885 33517 6888
rect 33551 6885 33563 6919
rect 33505 6879 33563 6885
rect 33134 6740 33140 6792
rect 33192 6780 33198 6792
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 33192 6752 33241 6780
rect 33192 6740 33198 6752
rect 33229 6749 33241 6752
rect 33275 6749 33287 6783
rect 33229 6743 33287 6749
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 57514 5896 57520 5908
rect 57475 5868 57520 5896
rect 57514 5856 57520 5868
rect 57572 5856 57578 5908
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2409 5695 2467 5701
rect 2409 5692 2421 5695
rect 1903 5664 2421 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2409 5661 2421 5664
rect 2455 5692 2467 5695
rect 20438 5692 20444 5704
rect 2455 5664 20444 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 57514 5652 57520 5704
rect 57572 5692 57578 5704
rect 58069 5695 58127 5701
rect 58069 5692 58081 5695
rect 57572 5664 58081 5692
rect 57572 5652 57578 5664
rect 58069 5661 58081 5664
rect 58115 5661 58127 5695
rect 58069 5655 58127 5661
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 58250 5556 58256 5568
rect 58211 5528 58256 5556
rect 58250 5516 58256 5528
rect 58308 5516 58314 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 27985 2635 28043 2641
rect 27985 2601 27997 2635
rect 28031 2632 28043 2635
rect 31662 2632 31668 2644
rect 28031 2604 31668 2632
rect 28031 2601 28043 2604
rect 27985 2595 28043 2601
rect 27338 2564 27344 2576
rect 6886 2536 27344 2564
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6886 2496 6914 2536
rect 27338 2524 27344 2536
rect 27396 2524 27402 2576
rect 14642 2496 14648 2508
rect 5767 2468 6914 2496
rect 10796 2468 14648 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 1872 2360 1900 2391
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5592 2400 6009 2428
rect 5592 2388 5598 2400
rect 5997 2397 6009 2400
rect 6043 2428 6055 2431
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6043 2400 6561 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 1872 2332 2421 2360
rect 2409 2329 2421 2332
rect 2455 2360 2467 2363
rect 10796 2360 10824 2468
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 17678 2496 17684 2508
rect 17639 2468 17684 2496
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 28000 2496 28028 2595
rect 31662 2592 31668 2604
rect 31720 2592 31726 2644
rect 37090 2592 37096 2644
rect 37148 2632 37154 2644
rect 37553 2635 37611 2641
rect 37553 2632 37565 2635
rect 37148 2604 37565 2632
rect 37148 2592 37154 2604
rect 37553 2601 37565 2604
rect 37599 2601 37611 2635
rect 44082 2632 44088 2644
rect 44043 2604 44088 2632
rect 37553 2595 37611 2601
rect 44082 2592 44088 2604
rect 44140 2592 44146 2644
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 44232 2604 51074 2632
rect 44232 2592 44238 2604
rect 34422 2524 34428 2576
rect 34480 2564 34486 2576
rect 34480 2536 48314 2564
rect 34480 2524 34486 2536
rect 43990 2496 43996 2508
rect 27448 2468 28028 2496
rect 31726 2468 43996 2496
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 17129 2431 17187 2437
rect 12023 2400 12572 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12544 2369 12572 2400
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17696 2428 17724 2456
rect 22278 2428 22284 2440
rect 17175 2400 17724 2428
rect 22239 2400 22284 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 27448 2437 27476 2468
rect 27433 2431 27491 2437
rect 25464 2400 27384 2428
rect 25464 2388 25470 2400
rect 2455 2332 10824 2360
rect 12529 2363 12587 2369
rect 2455 2329 2467 2332
rect 2409 2323 2467 2329
rect 12529 2329 12541 2363
rect 12575 2360 12587 2363
rect 22186 2360 22192 2372
rect 12575 2332 22192 2360
rect 12575 2329 12587 2332
rect 12529 2323 12587 2329
rect 22186 2320 22192 2332
rect 22244 2320 22250 2372
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11020 2264 11805 2292
rect 11020 2252 11026 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16172 2264 16957 2292
rect 16172 2252 16178 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21968 2264 22109 2292
rect 21968 2252 21974 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22097 2255 22155 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27249 2295 27307 2301
rect 27249 2292 27261 2295
rect 27120 2264 27261 2292
rect 27120 2252 27126 2264
rect 27249 2261 27261 2264
rect 27295 2261 27307 2295
rect 27356 2292 27384 2400
rect 27433 2397 27445 2431
rect 27479 2397 27491 2431
rect 27433 2391 27491 2397
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 31726 2428 31754 2468
rect 43990 2456 43996 2468
rect 44048 2456 44054 2508
rect 32950 2428 32956 2440
rect 27764 2400 31754 2428
rect 32911 2400 32956 2428
rect 27764 2388 27770 2400
rect 32950 2388 32956 2400
rect 33008 2388 33014 2440
rect 37090 2388 37096 2440
rect 37148 2428 37154 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37148 2400 38117 2428
rect 37148 2388 37154 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 43441 2431 43499 2437
rect 43441 2397 43453 2431
rect 43487 2428 43499 2431
rect 43806 2428 43812 2440
rect 43487 2400 43812 2428
rect 43487 2397 43499 2400
rect 43441 2391 43499 2397
rect 43806 2388 43812 2400
rect 43864 2428 43870 2440
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 43864 2400 43913 2428
rect 43864 2388 43870 2400
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 48286 2428 48314 2536
rect 51046 2496 51074 2604
rect 57425 2499 57483 2505
rect 57425 2496 57437 2499
rect 51046 2468 57437 2496
rect 57425 2465 57437 2468
rect 57471 2465 57483 2499
rect 57425 2459 57483 2465
rect 48501 2431 48559 2437
rect 48501 2428 48513 2431
rect 48286 2400 48513 2428
rect 43901 2391 43959 2397
rect 48501 2397 48513 2400
rect 48547 2428 48559 2431
rect 49053 2431 49111 2437
rect 49053 2428 49065 2431
rect 48547 2400 49065 2428
rect 48547 2397 48559 2400
rect 48501 2391 48559 2397
rect 49053 2397 49065 2400
rect 49099 2397 49111 2431
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 49053 2391 49111 2397
rect 55186 2400 55505 2428
rect 54849 2363 54907 2369
rect 54849 2360 54861 2363
rect 31726 2332 54861 2360
rect 31726 2292 31754 2332
rect 54849 2329 54861 2332
rect 54895 2360 54907 2363
rect 55186 2360 55214 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 57440 2428 57468 2459
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 57440 2400 58081 2428
rect 55493 2391 55551 2397
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 54895 2332 55214 2360
rect 54895 2329 54907 2332
rect 54849 2323 54907 2329
rect 27356 2264 31754 2292
rect 27249 2255 27307 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 33137 2295 33195 2301
rect 33137 2292 33149 2295
rect 32916 2264 33149 2292
rect 32916 2252 32922 2264
rect 33137 2261 33149 2264
rect 33183 2261 33195 2295
rect 33137 2255 33195 2261
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 38068 2264 38301 2292
rect 38068 2252 38074 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 48958 2252 48964 2304
rect 49016 2292 49022 2304
rect 49237 2295 49295 2301
rect 49237 2292 49249 2295
rect 49016 2264 49249 2292
rect 49016 2252 49022 2264
rect 49237 2261 49249 2264
rect 49283 2261 49295 2295
rect 49237 2255 49295 2261
rect 55122 2252 55128 2304
rect 55180 2292 55186 2304
rect 55677 2295 55735 2301
rect 55677 2292 55689 2295
rect 55180 2264 55689 2292
rect 55180 2252 55186 2264
rect 55677 2261 55689 2264
rect 55723 2261 55735 2295
rect 55677 2255 55735 2261
rect 58253 2295 58311 2301
rect 58253 2261 58265 2295
rect 58299 2292 58311 2295
rect 59906 2292 59912 2304
rect 58299 2264 59912 2292
rect 58299 2261 58311 2264
rect 58253 2255 58311 2261
rect 59906 2252 59912 2264
rect 59964 2252 59970 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1676 57579 1728 57588
rect 1676 57545 1685 57579
rect 1685 57545 1719 57579
rect 1719 57545 1728 57579
rect 1676 57536 1728 57545
rect 8392 57536 8444 57588
rect 13544 57536 13596 57588
rect 19340 57536 19392 57588
rect 24492 57536 24544 57588
rect 35440 57536 35492 57588
rect 41420 57536 41472 57588
rect 46388 57536 46440 57588
rect 52184 57536 52236 57588
rect 57336 57536 57388 57588
rect 2596 57468 2648 57520
rect 30288 57468 30340 57520
rect 1860 57443 1912 57452
rect 1860 57409 1869 57443
rect 1869 57409 1903 57443
rect 1903 57409 1912 57443
rect 1860 57400 1912 57409
rect 9864 57400 9916 57452
rect 14280 57443 14332 57452
rect 14280 57409 14289 57443
rect 14289 57409 14323 57443
rect 14323 57409 14332 57443
rect 14280 57400 14332 57409
rect 25320 57400 25372 57452
rect 35532 57443 35584 57452
rect 35532 57409 35541 57443
rect 35541 57409 35575 57443
rect 35575 57409 35584 57443
rect 35532 57400 35584 57409
rect 41328 57443 41380 57452
rect 41328 57409 41337 57443
rect 41337 57409 41371 57443
rect 41371 57409 41380 57443
rect 41328 57400 41380 57409
rect 46480 57443 46532 57452
rect 46480 57409 46489 57443
rect 46489 57409 46523 57443
rect 46523 57409 46532 57443
rect 46480 57400 46532 57409
rect 52276 57400 52328 57452
rect 32404 57332 32456 57384
rect 2872 57239 2924 57248
rect 2872 57205 2881 57239
rect 2881 57205 2915 57239
rect 2915 57205 2924 57239
rect 2872 57196 2924 57205
rect 9864 57239 9916 57248
rect 9864 57205 9873 57239
rect 9873 57205 9907 57239
rect 9907 57205 9916 57239
rect 9864 57196 9916 57205
rect 25320 57239 25372 57248
rect 25320 57205 25329 57239
rect 25329 57205 25363 57239
rect 25363 57205 25372 57239
rect 25320 57196 25372 57205
rect 30564 57239 30616 57248
rect 30564 57205 30573 57239
rect 30573 57205 30607 57239
rect 30607 57205 30616 57239
rect 30564 57196 30616 57205
rect 52276 57239 52328 57248
rect 52276 57205 52285 57239
rect 52285 57205 52319 57239
rect 52319 57205 52328 57239
rect 52276 57196 52328 57205
rect 57152 57196 57204 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 2596 57035 2648 57044
rect 2596 57001 2605 57035
rect 2605 57001 2639 57035
rect 2639 57001 2648 57035
rect 2596 56992 2648 57001
rect 35532 56992 35584 57044
rect 58256 57035 58308 57044
rect 58256 57001 58265 57035
rect 58265 57001 58299 57035
rect 58299 57001 58308 57035
rect 58256 56992 58308 57001
rect 1860 56652 1912 56704
rect 35624 56652 35676 56704
rect 57612 56695 57664 56704
rect 57612 56661 57621 56695
rect 57621 56661 57655 56695
rect 57655 56661 57664 56695
rect 57612 56652 57664 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 2136 51960 2188 52012
rect 1676 51799 1728 51808
rect 1676 51765 1685 51799
rect 1685 51765 1719 51799
rect 1719 51765 1728 51799
rect 1676 51756 1728 51765
rect 2136 51756 2188 51808
rect 57244 51756 57296 51808
rect 58256 51799 58308 51808
rect 58256 51765 58265 51799
rect 58265 51765 58299 51799
rect 58299 51765 58308 51799
rect 58256 51756 58308 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 29736 47991 29788 48000
rect 29736 47957 29745 47991
rect 29745 47957 29779 47991
rect 29779 47957 29788 47991
rect 29736 47948 29788 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 25964 47744 26016 47796
rect 27252 47676 27304 47728
rect 28264 47651 28316 47660
rect 28264 47617 28273 47651
rect 28273 47617 28307 47651
rect 28307 47617 28316 47651
rect 28264 47608 28316 47617
rect 28448 47651 28500 47660
rect 28448 47617 28457 47651
rect 28457 47617 28491 47651
rect 28491 47617 28500 47651
rect 28448 47608 28500 47617
rect 31760 47676 31812 47728
rect 32588 47608 32640 47660
rect 22376 47447 22428 47456
rect 22376 47413 22385 47447
rect 22385 47413 22419 47447
rect 22419 47413 22428 47447
rect 22376 47404 22428 47413
rect 23204 47404 23256 47456
rect 25780 47540 25832 47592
rect 29368 47540 29420 47592
rect 33232 47583 33284 47592
rect 33232 47549 33241 47583
rect 33241 47549 33275 47583
rect 33275 47549 33284 47583
rect 33232 47540 33284 47549
rect 24676 47404 24728 47456
rect 31024 47472 31076 47524
rect 29736 47404 29788 47456
rect 31300 47447 31352 47456
rect 31300 47413 31309 47447
rect 31309 47413 31343 47447
rect 31343 47413 31352 47447
rect 31300 47404 31352 47413
rect 34428 47404 34480 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 32588 47243 32640 47252
rect 25228 47132 25280 47184
rect 26976 47132 27028 47184
rect 28632 47132 28684 47184
rect 21272 47064 21324 47116
rect 23020 47039 23072 47048
rect 22100 46971 22152 46980
rect 22100 46937 22109 46971
rect 22109 46937 22143 46971
rect 22143 46937 22152 46971
rect 23020 47005 23029 47039
rect 23029 47005 23063 47039
rect 23063 47005 23072 47039
rect 23020 46996 23072 47005
rect 25964 47064 26016 47116
rect 32588 47209 32597 47243
rect 32597 47209 32631 47243
rect 32631 47209 32640 47243
rect 32588 47200 32640 47209
rect 24768 46996 24820 47048
rect 25136 47039 25188 47048
rect 25136 47005 25145 47039
rect 25145 47005 25179 47039
rect 25179 47005 25188 47039
rect 25136 46996 25188 47005
rect 26516 47039 26568 47048
rect 26516 47005 26525 47039
rect 26525 47005 26559 47039
rect 26559 47005 26568 47039
rect 26516 46996 26568 47005
rect 26792 47039 26844 47048
rect 26792 47005 26801 47039
rect 26801 47005 26835 47039
rect 26835 47005 26844 47039
rect 28908 47064 28960 47116
rect 31760 47107 31812 47116
rect 31760 47073 31769 47107
rect 31769 47073 31803 47107
rect 31803 47073 31812 47107
rect 31760 47064 31812 47073
rect 26792 46996 26844 47005
rect 22100 46928 22152 46937
rect 24676 46928 24728 46980
rect 23296 46860 23348 46912
rect 25780 46928 25832 46980
rect 28540 46996 28592 47048
rect 30932 46996 30984 47048
rect 31024 47039 31076 47048
rect 31024 47005 31033 47039
rect 31033 47005 31067 47039
rect 31067 47005 31076 47039
rect 31024 46996 31076 47005
rect 30104 46928 30156 46980
rect 31300 46928 31352 46980
rect 33600 46928 33652 46980
rect 25320 46903 25372 46912
rect 25320 46869 25329 46903
rect 25329 46869 25363 46903
rect 25363 46869 25372 46903
rect 25320 46860 25372 46869
rect 26056 46860 26108 46912
rect 26332 46903 26384 46912
rect 26332 46869 26341 46903
rect 26341 46869 26375 46903
rect 26375 46869 26384 46903
rect 26332 46860 26384 46869
rect 27620 46860 27672 46912
rect 28724 46903 28776 46912
rect 28724 46869 28733 46903
rect 28733 46869 28767 46903
rect 28767 46869 28776 46903
rect 28724 46860 28776 46869
rect 28908 46860 28960 46912
rect 32312 46860 32364 46912
rect 33324 46903 33376 46912
rect 33324 46869 33333 46903
rect 33333 46869 33367 46903
rect 33367 46869 33376 46903
rect 33324 46860 33376 46869
rect 33968 46903 34020 46912
rect 33968 46869 33977 46903
rect 33977 46869 34011 46903
rect 34011 46869 34020 46903
rect 33968 46860 34020 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 27712 46656 27764 46708
rect 28724 46656 28776 46708
rect 33324 46656 33376 46708
rect 2320 46520 2372 46572
rect 21272 46563 21324 46572
rect 21272 46529 21281 46563
rect 21281 46529 21315 46563
rect 21315 46529 21324 46563
rect 21272 46520 21324 46529
rect 21548 46520 21600 46572
rect 22376 46520 22428 46572
rect 23020 46520 23072 46572
rect 25136 46588 25188 46640
rect 24032 46427 24084 46436
rect 24032 46393 24041 46427
rect 24041 46393 24075 46427
rect 24075 46393 24084 46427
rect 24676 46520 24728 46572
rect 25228 46563 25280 46572
rect 25228 46529 25237 46563
rect 25237 46529 25271 46563
rect 25271 46529 25280 46563
rect 25228 46520 25280 46529
rect 26056 46520 26108 46572
rect 26516 46588 26568 46640
rect 27896 46588 27948 46640
rect 26700 46520 26752 46572
rect 27712 46520 27764 46572
rect 24308 46495 24360 46504
rect 24308 46461 24317 46495
rect 24317 46461 24351 46495
rect 24351 46461 24360 46495
rect 24308 46452 24360 46461
rect 24768 46452 24820 46504
rect 28540 46520 28592 46572
rect 30656 46588 30708 46640
rect 32312 46588 32364 46640
rect 33140 46588 33192 46640
rect 29184 46520 29236 46572
rect 29736 46520 29788 46572
rect 31300 46520 31352 46572
rect 25136 46427 25188 46436
rect 24032 46384 24084 46393
rect 25136 46393 25145 46427
rect 25145 46393 25179 46427
rect 25179 46393 25188 46427
rect 25136 46384 25188 46393
rect 1676 46359 1728 46368
rect 1676 46325 1685 46359
rect 1685 46325 1719 46359
rect 1719 46325 1728 46359
rect 1676 46316 1728 46325
rect 2320 46359 2372 46368
rect 2320 46325 2329 46359
rect 2329 46325 2363 46359
rect 2363 46325 2372 46359
rect 2320 46316 2372 46325
rect 20812 46316 20864 46368
rect 22100 46316 22152 46368
rect 23664 46316 23716 46368
rect 23848 46359 23900 46368
rect 23848 46325 23857 46359
rect 23857 46325 23891 46359
rect 23891 46325 23900 46359
rect 23848 46316 23900 46325
rect 24768 46316 24820 46368
rect 25872 46359 25924 46368
rect 25872 46325 25881 46359
rect 25881 46325 25915 46359
rect 25915 46325 25924 46359
rect 25872 46316 25924 46325
rect 26792 46384 26844 46436
rect 28264 46384 28316 46436
rect 28908 46384 28960 46436
rect 30288 46384 30340 46436
rect 32312 46452 32364 46504
rect 32496 46520 32548 46572
rect 32588 46452 32640 46504
rect 27436 46316 27488 46368
rect 28448 46359 28500 46368
rect 28448 46325 28457 46359
rect 28457 46325 28491 46359
rect 28491 46325 28500 46359
rect 28448 46316 28500 46325
rect 28540 46316 28592 46368
rect 29276 46359 29328 46368
rect 29276 46325 29285 46359
rect 29285 46325 29319 46359
rect 29319 46325 29328 46359
rect 29276 46316 29328 46325
rect 29736 46359 29788 46368
rect 29736 46325 29745 46359
rect 29745 46325 29779 46359
rect 29779 46325 29788 46359
rect 29736 46316 29788 46325
rect 30656 46316 30708 46368
rect 31852 46316 31904 46368
rect 33784 46316 33836 46368
rect 34152 46359 34204 46368
rect 34152 46325 34161 46359
rect 34161 46325 34195 46359
rect 34195 46325 34204 46359
rect 34152 46316 34204 46325
rect 34704 46359 34756 46368
rect 34704 46325 34713 46359
rect 34713 46325 34747 46359
rect 34747 46325 34756 46359
rect 34704 46316 34756 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 29276 46112 29328 46164
rect 31208 46112 31260 46164
rect 22376 46044 22428 46096
rect 27344 46044 27396 46096
rect 27988 46044 28040 46096
rect 30748 46087 30800 46096
rect 22560 45951 22612 45960
rect 22560 45917 22569 45951
rect 22569 45917 22603 45951
rect 22603 45917 22612 45951
rect 22560 45908 22612 45917
rect 23204 45908 23256 45960
rect 24032 45976 24084 46028
rect 24584 45976 24636 46028
rect 27436 45976 27488 46028
rect 24308 45908 24360 45960
rect 24952 45951 25004 45960
rect 22284 45840 22336 45892
rect 23572 45840 23624 45892
rect 24952 45917 24961 45951
rect 24961 45917 24995 45951
rect 24995 45917 25004 45951
rect 24952 45908 25004 45917
rect 26148 45908 26200 45960
rect 26700 45908 26752 45960
rect 26976 45951 27028 45960
rect 26976 45917 26985 45951
rect 26985 45917 27019 45951
rect 27019 45917 27028 45951
rect 27804 45976 27856 46028
rect 28264 45976 28316 46028
rect 30748 46053 30757 46087
rect 30757 46053 30791 46087
rect 30791 46053 30800 46087
rect 30748 46044 30800 46053
rect 26976 45908 27028 45917
rect 26608 45840 26660 45892
rect 27712 45951 27764 45960
rect 27712 45917 27721 45951
rect 27721 45917 27755 45951
rect 27755 45917 27764 45951
rect 27896 45951 27948 45960
rect 27712 45908 27764 45917
rect 27896 45917 27905 45951
rect 27905 45917 27939 45951
rect 27939 45917 27948 45951
rect 27896 45908 27948 45917
rect 28908 45908 28960 45960
rect 29736 45908 29788 45960
rect 29184 45883 29236 45892
rect 29184 45849 29193 45883
rect 29193 45849 29227 45883
rect 29227 45849 29236 45883
rect 29184 45840 29236 45849
rect 29368 45840 29420 45892
rect 30288 45908 30340 45960
rect 30656 46019 30708 46028
rect 30656 45985 30665 46019
rect 30665 45985 30699 46019
rect 30699 45985 30708 46019
rect 31852 46019 31904 46028
rect 30656 45976 30708 45985
rect 31852 45985 31861 46019
rect 31861 45985 31895 46019
rect 31895 45985 31904 46019
rect 31852 45976 31904 45985
rect 33324 45976 33376 46028
rect 32496 45908 32548 45960
rect 33600 45908 33652 45960
rect 33784 45908 33836 45960
rect 1860 45772 1912 45824
rect 20444 45815 20496 45824
rect 20444 45781 20453 45815
rect 20453 45781 20487 45815
rect 20487 45781 20496 45815
rect 20444 45772 20496 45781
rect 21088 45772 21140 45824
rect 22376 45815 22428 45824
rect 22376 45781 22385 45815
rect 22385 45781 22419 45815
rect 22419 45781 22428 45815
rect 22376 45772 22428 45781
rect 22744 45815 22796 45824
rect 22744 45781 22753 45815
rect 22753 45781 22787 45815
rect 22787 45781 22796 45815
rect 22744 45772 22796 45781
rect 23480 45772 23532 45824
rect 24032 45772 24084 45824
rect 27344 45772 27396 45824
rect 31300 45772 31352 45824
rect 33876 45815 33928 45824
rect 33876 45781 33885 45815
rect 33885 45781 33919 45815
rect 33919 45781 33928 45815
rect 33876 45772 33928 45781
rect 33968 45772 34020 45824
rect 34704 45772 34756 45824
rect 57336 45772 57388 45824
rect 58256 45815 58308 45824
rect 58256 45781 58265 45815
rect 58265 45781 58299 45815
rect 58299 45781 58308 45815
rect 58256 45772 58308 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 22376 45568 22428 45620
rect 22560 45568 22612 45620
rect 25136 45568 25188 45620
rect 30932 45611 30984 45620
rect 20720 45432 20772 45484
rect 20904 45432 20956 45484
rect 21456 45500 21508 45552
rect 24860 45500 24912 45552
rect 27252 45543 27304 45552
rect 27252 45509 27261 45543
rect 27261 45509 27295 45543
rect 27295 45509 27304 45543
rect 27252 45500 27304 45509
rect 21364 45432 21416 45484
rect 22192 45475 22244 45484
rect 22192 45441 22201 45475
rect 22201 45441 22235 45475
rect 22235 45441 22244 45475
rect 22192 45432 22244 45441
rect 22376 45432 22428 45484
rect 23296 45475 23348 45484
rect 23296 45441 23305 45475
rect 23305 45441 23339 45475
rect 23339 45441 23348 45475
rect 23296 45432 23348 45441
rect 21088 45407 21140 45416
rect 21088 45373 21097 45407
rect 21097 45373 21131 45407
rect 21131 45373 21140 45407
rect 21088 45364 21140 45373
rect 23480 45364 23532 45416
rect 24308 45364 24360 45416
rect 25504 45475 25556 45484
rect 25504 45441 25513 45475
rect 25513 45441 25547 45475
rect 25547 45441 25556 45475
rect 25504 45432 25556 45441
rect 26148 45432 26200 45484
rect 26424 45475 26476 45484
rect 26424 45441 26433 45475
rect 26433 45441 26467 45475
rect 26467 45441 26476 45475
rect 26424 45432 26476 45441
rect 26608 45475 26660 45484
rect 26608 45441 26617 45475
rect 26617 45441 26651 45475
rect 26651 45441 26660 45475
rect 26608 45432 26660 45441
rect 29092 45500 29144 45552
rect 29736 45500 29788 45552
rect 24676 45339 24728 45348
rect 21180 45228 21232 45280
rect 22652 45271 22704 45280
rect 22652 45237 22661 45271
rect 22661 45237 22695 45271
rect 22695 45237 22704 45271
rect 22652 45228 22704 45237
rect 23112 45271 23164 45280
rect 23112 45237 23121 45271
rect 23121 45237 23155 45271
rect 23155 45237 23164 45271
rect 23112 45228 23164 45237
rect 23204 45228 23256 45280
rect 24676 45305 24685 45339
rect 24685 45305 24719 45339
rect 24719 45305 24728 45339
rect 24676 45296 24728 45305
rect 24952 45364 25004 45416
rect 25228 45296 25280 45348
rect 25688 45296 25740 45348
rect 27436 45364 27488 45416
rect 28908 45432 28960 45484
rect 30932 45577 30941 45611
rect 30941 45577 30975 45611
rect 30975 45577 30984 45611
rect 30932 45568 30984 45577
rect 31024 45611 31076 45620
rect 31024 45577 31033 45611
rect 31033 45577 31067 45611
rect 31067 45577 31076 45611
rect 31024 45568 31076 45577
rect 31208 45568 31260 45620
rect 33416 45568 33468 45620
rect 34520 45500 34572 45552
rect 30656 45432 30708 45484
rect 31024 45432 31076 45484
rect 31300 45432 31352 45484
rect 33324 45432 33376 45484
rect 33600 45475 33652 45484
rect 33600 45441 33609 45475
rect 33609 45441 33643 45475
rect 33643 45441 33652 45475
rect 33600 45432 33652 45441
rect 26884 45296 26936 45348
rect 27804 45296 27856 45348
rect 28080 45296 28132 45348
rect 30840 45296 30892 45348
rect 33968 45432 34020 45484
rect 34428 45475 34480 45484
rect 34428 45441 34437 45475
rect 34437 45441 34471 45475
rect 34471 45441 34480 45475
rect 34428 45432 34480 45441
rect 32312 45296 32364 45348
rect 32588 45296 32640 45348
rect 24400 45271 24452 45280
rect 24400 45237 24409 45271
rect 24409 45237 24443 45271
rect 24443 45237 24452 45271
rect 24400 45228 24452 45237
rect 25780 45271 25832 45280
rect 25780 45237 25789 45271
rect 25789 45237 25823 45271
rect 25823 45237 25832 45271
rect 25780 45228 25832 45237
rect 26516 45271 26568 45280
rect 26516 45237 26525 45271
rect 26525 45237 26559 45271
rect 26559 45237 26568 45271
rect 26516 45228 26568 45237
rect 27528 45228 27580 45280
rect 28356 45271 28408 45280
rect 28356 45237 28365 45271
rect 28365 45237 28399 45271
rect 28399 45237 28408 45271
rect 28356 45228 28408 45237
rect 29736 45271 29788 45280
rect 29736 45237 29745 45271
rect 29745 45237 29779 45271
rect 29779 45237 29788 45271
rect 29736 45228 29788 45237
rect 30104 45271 30156 45280
rect 30104 45237 30113 45271
rect 30113 45237 30147 45271
rect 30147 45237 30156 45271
rect 30104 45228 30156 45237
rect 31300 45228 31352 45280
rect 34428 45228 34480 45280
rect 35900 45271 35952 45280
rect 35900 45237 35909 45271
rect 35909 45237 35943 45271
rect 35943 45237 35952 45271
rect 35900 45228 35952 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 21088 44888 21140 44940
rect 22192 45024 22244 45076
rect 26884 45024 26936 45076
rect 34152 45067 34204 45076
rect 22376 44956 22428 45008
rect 20996 44820 21048 44872
rect 21456 44863 21508 44872
rect 21456 44829 21465 44863
rect 21465 44829 21499 44863
rect 21499 44829 21508 44863
rect 22192 44888 22244 44940
rect 22468 44863 22520 44872
rect 21456 44820 21508 44829
rect 22468 44829 22477 44863
rect 22477 44829 22511 44863
rect 22511 44829 22520 44863
rect 22468 44820 22520 44829
rect 23388 44888 23440 44940
rect 22008 44752 22060 44804
rect 22100 44752 22152 44804
rect 20536 44684 20588 44736
rect 20628 44684 20680 44736
rect 22468 44684 22520 44736
rect 22836 44863 22888 44872
rect 22836 44829 22845 44863
rect 22845 44829 22879 44863
rect 22879 44829 22888 44863
rect 23480 44863 23532 44872
rect 22836 44820 22888 44829
rect 23480 44829 23489 44863
rect 23489 44829 23523 44863
rect 23523 44829 23532 44863
rect 23480 44820 23532 44829
rect 23940 44820 23992 44872
rect 24860 44888 24912 44940
rect 25228 44888 25280 44940
rect 26148 44956 26200 45008
rect 28724 44956 28776 45008
rect 25596 44863 25648 44872
rect 25596 44829 25605 44863
rect 25605 44829 25639 44863
rect 25639 44829 25648 44863
rect 25596 44820 25648 44829
rect 25780 44863 25832 44872
rect 25780 44829 25789 44863
rect 25789 44829 25823 44863
rect 25823 44829 25832 44863
rect 26424 44888 26476 44940
rect 27804 44888 27856 44940
rect 34152 45033 34161 45067
rect 34161 45033 34195 45067
rect 34195 45033 34204 45067
rect 34152 45024 34204 45033
rect 32128 44999 32180 45008
rect 32128 44965 32137 44999
rect 32137 44965 32171 44999
rect 32171 44965 32180 44999
rect 32128 44956 32180 44965
rect 25780 44820 25832 44829
rect 25504 44752 25556 44804
rect 27528 44820 27580 44872
rect 27896 44820 27948 44872
rect 28080 44863 28132 44872
rect 28080 44829 28089 44863
rect 28089 44829 28123 44863
rect 28123 44829 28132 44863
rect 28080 44820 28132 44829
rect 29092 44820 29144 44872
rect 29368 44820 29420 44872
rect 27436 44795 27488 44804
rect 27436 44761 27445 44795
rect 27445 44761 27479 44795
rect 27479 44761 27488 44795
rect 27436 44752 27488 44761
rect 29828 44820 29880 44872
rect 30564 44888 30616 44940
rect 32496 44888 32548 44940
rect 30288 44820 30340 44872
rect 30932 44820 30984 44872
rect 29644 44752 29696 44804
rect 30656 44752 30708 44804
rect 33140 44820 33192 44872
rect 33508 44820 33560 44872
rect 33600 44863 33652 44872
rect 33600 44829 33609 44863
rect 33609 44829 33643 44863
rect 33643 44829 33652 44863
rect 33600 44820 33652 44829
rect 33232 44752 33284 44804
rect 22744 44684 22796 44736
rect 23020 44684 23072 44736
rect 25320 44727 25372 44736
rect 25320 44693 25329 44727
rect 25329 44693 25363 44727
rect 25363 44693 25372 44727
rect 25320 44684 25372 44693
rect 25688 44684 25740 44736
rect 28908 44684 28960 44736
rect 30012 44684 30064 44736
rect 31300 44727 31352 44736
rect 31300 44693 31309 44727
rect 31309 44693 31343 44727
rect 31343 44693 31352 44727
rect 31300 44684 31352 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 21456 44480 21508 44532
rect 22836 44480 22888 44532
rect 23480 44480 23532 44532
rect 24308 44480 24360 44532
rect 25688 44480 25740 44532
rect 20444 44455 20496 44464
rect 20444 44421 20453 44455
rect 20453 44421 20487 44455
rect 20487 44421 20496 44455
rect 20444 44412 20496 44421
rect 18696 44344 18748 44396
rect 21088 44412 21140 44464
rect 19432 44319 19484 44328
rect 19432 44285 19441 44319
rect 19441 44285 19475 44319
rect 19475 44285 19484 44319
rect 19432 44276 19484 44285
rect 19156 44140 19208 44192
rect 22008 44387 22060 44396
rect 20536 44276 20588 44328
rect 22008 44353 22017 44387
rect 22017 44353 22051 44387
rect 22051 44353 22060 44387
rect 22008 44344 22060 44353
rect 22192 44387 22244 44396
rect 22192 44353 22201 44387
rect 22201 44353 22235 44387
rect 22235 44353 22244 44387
rect 22192 44344 22244 44353
rect 22836 44344 22888 44396
rect 21732 44276 21784 44328
rect 22284 44276 22336 44328
rect 23756 44344 23808 44396
rect 24216 44344 24268 44396
rect 23664 44276 23716 44328
rect 24584 44344 24636 44396
rect 25136 44387 25188 44396
rect 25136 44353 25145 44387
rect 25145 44353 25179 44387
rect 25179 44353 25188 44387
rect 25136 44344 25188 44353
rect 25964 44344 26016 44396
rect 26700 44344 26752 44396
rect 27896 44387 27948 44396
rect 27160 44276 27212 44328
rect 27896 44353 27905 44387
rect 27905 44353 27939 44387
rect 27939 44353 27948 44387
rect 27896 44344 27948 44353
rect 28908 44387 28960 44396
rect 28908 44353 28917 44387
rect 28917 44353 28951 44387
rect 28951 44353 28960 44387
rect 28908 44344 28960 44353
rect 29644 44412 29696 44464
rect 29828 44480 29880 44532
rect 32312 44480 32364 44532
rect 34152 44480 34204 44532
rect 29552 44387 29604 44396
rect 29552 44353 29561 44387
rect 29561 44353 29595 44387
rect 29595 44353 29604 44387
rect 29552 44344 29604 44353
rect 31852 44412 31904 44464
rect 30288 44387 30340 44396
rect 30288 44353 30297 44387
rect 30297 44353 30331 44387
rect 30331 44353 30340 44387
rect 30288 44344 30340 44353
rect 31116 44344 31168 44396
rect 31392 44344 31444 44396
rect 34428 44412 34480 44464
rect 33324 44344 33376 44396
rect 27528 44276 27580 44328
rect 30380 44319 30432 44328
rect 30380 44285 30389 44319
rect 30389 44285 30423 44319
rect 30423 44285 30432 44319
rect 30380 44276 30432 44285
rect 33232 44319 33284 44328
rect 33232 44285 33241 44319
rect 33241 44285 33275 44319
rect 33275 44285 33284 44319
rect 33232 44276 33284 44285
rect 33508 44344 33560 44396
rect 34428 44276 34480 44328
rect 22008 44208 22060 44260
rect 22192 44183 22244 44192
rect 22192 44149 22201 44183
rect 22201 44149 22235 44183
rect 22235 44149 22244 44183
rect 22192 44140 22244 44149
rect 23664 44140 23716 44192
rect 23940 44208 23992 44260
rect 29736 44208 29788 44260
rect 24124 44140 24176 44192
rect 24952 44183 25004 44192
rect 24952 44149 24961 44183
rect 24961 44149 24995 44183
rect 24995 44149 25004 44183
rect 24952 44140 25004 44149
rect 25228 44140 25280 44192
rect 26424 44183 26476 44192
rect 26424 44149 26433 44183
rect 26433 44149 26467 44183
rect 26467 44149 26476 44183
rect 26424 44140 26476 44149
rect 27160 44140 27212 44192
rect 28080 44183 28132 44192
rect 28080 44149 28089 44183
rect 28089 44149 28123 44183
rect 28123 44149 28132 44183
rect 28080 44140 28132 44149
rect 29092 44183 29144 44192
rect 29092 44149 29101 44183
rect 29101 44149 29135 44183
rect 29135 44149 29144 44183
rect 29092 44140 29144 44149
rect 29368 44140 29420 44192
rect 31024 44183 31076 44192
rect 31024 44149 31033 44183
rect 31033 44149 31067 44183
rect 31067 44149 31076 44183
rect 31024 44140 31076 44149
rect 32404 44183 32456 44192
rect 32404 44149 32413 44183
rect 32413 44149 32447 44183
rect 32447 44149 32456 44183
rect 32404 44140 32456 44149
rect 33876 44251 33928 44260
rect 33876 44217 33885 44251
rect 33885 44217 33919 44251
rect 33919 44217 33928 44251
rect 33876 44208 33928 44217
rect 35348 44140 35400 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 20536 43936 20588 43988
rect 22192 43936 22244 43988
rect 23848 43979 23900 43988
rect 23848 43945 23857 43979
rect 23857 43945 23891 43979
rect 23891 43945 23900 43979
rect 23848 43936 23900 43945
rect 24308 43936 24360 43988
rect 18696 43775 18748 43784
rect 18696 43741 18705 43775
rect 18705 43741 18739 43775
rect 18739 43741 18748 43775
rect 18696 43732 18748 43741
rect 19432 43800 19484 43852
rect 20628 43800 20680 43852
rect 26240 43936 26292 43988
rect 29920 43936 29972 43988
rect 30564 43936 30616 43988
rect 31208 43936 31260 43988
rect 33416 43936 33468 43988
rect 33876 43936 33928 43988
rect 21916 43800 21968 43852
rect 20352 43775 20404 43784
rect 20352 43741 20361 43775
rect 20361 43741 20395 43775
rect 20395 43741 20404 43775
rect 20352 43732 20404 43741
rect 18604 43639 18656 43648
rect 18604 43605 18613 43639
rect 18613 43605 18647 43639
rect 18647 43605 18656 43639
rect 18604 43596 18656 43605
rect 19340 43596 19392 43648
rect 20444 43664 20496 43716
rect 20628 43664 20680 43716
rect 21364 43732 21416 43784
rect 23296 43732 23348 43784
rect 21824 43664 21876 43716
rect 22376 43664 22428 43716
rect 24308 43732 24360 43784
rect 25596 43775 25648 43784
rect 25596 43741 25605 43775
rect 25605 43741 25639 43775
rect 25639 43741 25648 43775
rect 25596 43732 25648 43741
rect 25780 43732 25832 43784
rect 25964 43732 26016 43784
rect 29092 43868 29144 43920
rect 26240 43732 26292 43784
rect 26516 43732 26568 43784
rect 27160 43775 27212 43784
rect 27160 43741 27169 43775
rect 27169 43741 27203 43775
rect 27203 43741 27212 43775
rect 27160 43732 27212 43741
rect 24124 43664 24176 43716
rect 27988 43732 28040 43784
rect 29184 43800 29236 43852
rect 31116 43868 31168 43920
rect 31852 43911 31904 43920
rect 31852 43877 31861 43911
rect 31861 43877 31895 43911
rect 31895 43877 31904 43911
rect 31852 43868 31904 43877
rect 28264 43732 28316 43784
rect 28632 43732 28684 43784
rect 34980 43843 35032 43852
rect 34980 43809 34989 43843
rect 34989 43809 35023 43843
rect 35023 43809 35032 43843
rect 34980 43800 35032 43809
rect 29828 43732 29880 43784
rect 30012 43775 30064 43784
rect 30012 43741 30021 43775
rect 30021 43741 30055 43775
rect 30055 43741 30064 43775
rect 30012 43732 30064 43741
rect 30656 43732 30708 43784
rect 31024 43775 31076 43784
rect 31024 43741 31033 43775
rect 31033 43741 31067 43775
rect 31067 43741 31076 43775
rect 31024 43732 31076 43741
rect 31116 43732 31168 43784
rect 31300 43732 31352 43784
rect 32404 43732 32456 43784
rect 35348 43732 35400 43784
rect 29460 43664 29512 43716
rect 30472 43664 30524 43716
rect 32588 43707 32640 43716
rect 32588 43673 32597 43707
rect 32597 43673 32631 43707
rect 32631 43673 32640 43707
rect 32588 43664 32640 43673
rect 33324 43664 33376 43716
rect 22560 43596 22612 43648
rect 23480 43639 23532 43648
rect 23480 43605 23489 43639
rect 23489 43605 23523 43639
rect 23523 43605 23532 43639
rect 23480 43596 23532 43605
rect 24032 43596 24084 43648
rect 25044 43596 25096 43648
rect 28264 43639 28316 43648
rect 28264 43605 28273 43639
rect 28273 43605 28307 43639
rect 28307 43605 28316 43639
rect 28264 43596 28316 43605
rect 28908 43639 28960 43648
rect 28908 43605 28917 43639
rect 28917 43605 28951 43639
rect 28951 43605 28960 43639
rect 28908 43596 28960 43605
rect 29736 43639 29788 43648
rect 29736 43605 29745 43639
rect 29745 43605 29779 43639
rect 29779 43605 29788 43639
rect 29736 43596 29788 43605
rect 31484 43596 31536 43648
rect 35808 43596 35860 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 18604 43324 18656 43376
rect 19984 43256 20036 43308
rect 19156 43188 19208 43240
rect 20260 43299 20312 43308
rect 20260 43265 20269 43299
rect 20269 43265 20303 43299
rect 20303 43265 20312 43299
rect 22100 43324 22152 43376
rect 22284 43324 22336 43376
rect 24124 43392 24176 43444
rect 25596 43392 25648 43444
rect 26516 43392 26568 43444
rect 20260 43256 20312 43265
rect 20996 43256 21048 43308
rect 21180 43299 21232 43308
rect 21180 43265 21189 43299
rect 21189 43265 21223 43299
rect 21223 43265 21232 43299
rect 22468 43299 22520 43308
rect 21180 43256 21232 43265
rect 22468 43265 22477 43299
rect 22477 43265 22511 43299
rect 22511 43265 22520 43299
rect 22468 43256 22520 43265
rect 24768 43324 24820 43376
rect 26332 43324 26384 43376
rect 27528 43367 27580 43376
rect 27528 43333 27537 43367
rect 27537 43333 27571 43367
rect 27571 43333 27580 43367
rect 27528 43324 27580 43333
rect 29184 43392 29236 43444
rect 32128 43392 32180 43444
rect 20352 43120 20404 43172
rect 22192 43120 22244 43172
rect 23480 43256 23532 43308
rect 23756 43299 23808 43308
rect 23756 43265 23765 43299
rect 23765 43265 23799 43299
rect 23799 43265 23808 43299
rect 23756 43256 23808 43265
rect 23940 43299 23992 43308
rect 23940 43265 23948 43299
rect 23948 43265 23982 43299
rect 23982 43265 23992 43299
rect 23940 43256 23992 43265
rect 24124 43256 24176 43308
rect 24216 43256 24268 43308
rect 24676 43299 24728 43308
rect 24676 43265 24685 43299
rect 24685 43265 24719 43299
rect 24719 43265 24728 43299
rect 24676 43256 24728 43265
rect 25504 43256 25556 43308
rect 25780 43256 25832 43308
rect 25964 43256 26016 43308
rect 28264 43299 28316 43308
rect 28264 43265 28273 43299
rect 28273 43265 28307 43299
rect 28307 43265 28316 43299
rect 28264 43256 28316 43265
rect 23572 43120 23624 43172
rect 25596 43120 25648 43172
rect 27068 43188 27120 43240
rect 28448 43188 28500 43240
rect 26608 43120 26660 43172
rect 27160 43163 27212 43172
rect 27160 43129 27169 43163
rect 27169 43129 27203 43163
rect 27203 43129 27212 43163
rect 27160 43120 27212 43129
rect 27252 43120 27304 43172
rect 28264 43120 28316 43172
rect 19248 43095 19300 43104
rect 19248 43061 19257 43095
rect 19257 43061 19291 43095
rect 19291 43061 19300 43095
rect 19248 43052 19300 43061
rect 19432 43052 19484 43104
rect 22560 43052 22612 43104
rect 24768 43052 24820 43104
rect 26056 43052 26108 43104
rect 27896 43052 27948 43104
rect 29368 43299 29420 43308
rect 29368 43265 29377 43299
rect 29377 43265 29411 43299
rect 29411 43265 29420 43299
rect 29368 43256 29420 43265
rect 29460 43256 29512 43308
rect 29828 43120 29880 43172
rect 30196 43120 30248 43172
rect 30012 43052 30064 43104
rect 32404 43367 32456 43376
rect 32404 43333 32413 43367
rect 32413 43333 32447 43367
rect 32447 43333 32456 43367
rect 32404 43324 32456 43333
rect 33692 43299 33744 43308
rect 33692 43265 33701 43299
rect 33701 43265 33735 43299
rect 33735 43265 33744 43299
rect 33692 43256 33744 43265
rect 35440 43256 35492 43308
rect 31668 43188 31720 43240
rect 33508 43188 33560 43240
rect 35992 43120 36044 43172
rect 31300 43095 31352 43104
rect 31300 43061 31309 43095
rect 31309 43061 31343 43095
rect 31343 43061 31352 43095
rect 31300 43052 31352 43061
rect 32680 43095 32732 43104
rect 32680 43061 32689 43095
rect 32689 43061 32723 43095
rect 32723 43061 32732 43095
rect 32680 43052 32732 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 20260 42848 20312 42900
rect 24676 42848 24728 42900
rect 25504 42848 25556 42900
rect 29920 42848 29972 42900
rect 30288 42848 30340 42900
rect 30656 42848 30708 42900
rect 21824 42780 21876 42832
rect 25596 42780 25648 42832
rect 20628 42712 20680 42764
rect 20904 42712 20956 42764
rect 21916 42712 21968 42764
rect 20720 42687 20772 42696
rect 20352 42576 20404 42628
rect 20720 42653 20729 42687
rect 20729 42653 20763 42687
rect 20763 42653 20772 42687
rect 20720 42644 20772 42653
rect 21088 42644 21140 42696
rect 21456 42687 21508 42696
rect 21456 42653 21465 42687
rect 21465 42653 21499 42687
rect 21499 42653 21508 42687
rect 21456 42644 21508 42653
rect 21732 42687 21784 42696
rect 21732 42653 21741 42687
rect 21741 42653 21775 42687
rect 21775 42653 21784 42687
rect 21732 42644 21784 42653
rect 22652 42712 22704 42764
rect 23204 42712 23256 42764
rect 20996 42576 21048 42628
rect 22744 42644 22796 42696
rect 23388 42644 23440 42696
rect 23664 42644 23716 42696
rect 23756 42644 23808 42696
rect 24676 42712 24728 42764
rect 26332 42780 26384 42832
rect 26976 42780 27028 42832
rect 26424 42712 26476 42764
rect 26792 42712 26844 42764
rect 27436 42712 27488 42764
rect 28172 42712 28224 42764
rect 29092 42780 29144 42832
rect 29460 42712 29512 42764
rect 24124 42576 24176 42628
rect 25044 42644 25096 42696
rect 25780 42687 25832 42696
rect 25780 42653 25789 42687
rect 25789 42653 25823 42687
rect 25823 42653 25832 42687
rect 25780 42644 25832 42653
rect 26056 42644 26108 42696
rect 27252 42687 27304 42696
rect 27252 42653 27261 42687
rect 27261 42653 27295 42687
rect 27295 42653 27304 42687
rect 27252 42644 27304 42653
rect 27344 42687 27396 42696
rect 27344 42653 27353 42687
rect 27353 42653 27387 42687
rect 27387 42653 27396 42687
rect 27344 42644 27396 42653
rect 29276 42644 29328 42696
rect 29736 42644 29788 42696
rect 30012 42644 30064 42696
rect 31944 42780 31996 42832
rect 32956 42780 33008 42832
rect 32404 42712 32456 42764
rect 32588 42712 32640 42764
rect 31760 42644 31812 42696
rect 35808 42712 35860 42764
rect 20260 42551 20312 42560
rect 20260 42517 20269 42551
rect 20269 42517 20303 42551
rect 20303 42517 20312 42551
rect 20260 42508 20312 42517
rect 21640 42508 21692 42560
rect 22192 42508 22244 42560
rect 22836 42508 22888 42560
rect 26148 42508 26200 42560
rect 27160 42508 27212 42560
rect 27528 42551 27580 42560
rect 27528 42517 27537 42551
rect 27537 42517 27571 42551
rect 27571 42517 27580 42551
rect 27528 42508 27580 42517
rect 28264 42551 28316 42560
rect 28264 42517 28273 42551
rect 28273 42517 28307 42551
rect 28307 42517 28316 42551
rect 28264 42508 28316 42517
rect 28448 42508 28500 42560
rect 31852 42576 31904 42628
rect 33784 42644 33836 42696
rect 33048 42576 33100 42628
rect 33508 42576 33560 42628
rect 29828 42508 29880 42560
rect 33416 42508 33468 42560
rect 33692 42508 33744 42560
rect 35808 42551 35860 42560
rect 35808 42517 35817 42551
rect 35817 42517 35851 42551
rect 35851 42517 35860 42551
rect 35808 42508 35860 42517
rect 37096 42508 37148 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 20628 42304 20680 42356
rect 21732 42304 21784 42356
rect 20168 42236 20220 42288
rect 20444 42168 20496 42220
rect 20904 42236 20956 42288
rect 21824 42236 21876 42288
rect 23664 42304 23716 42356
rect 26056 42304 26108 42356
rect 27988 42304 28040 42356
rect 28816 42304 28868 42356
rect 20720 42168 20772 42220
rect 22008 42168 22060 42220
rect 23480 42236 23532 42288
rect 23848 42236 23900 42288
rect 22744 42168 22796 42220
rect 23664 42211 23716 42220
rect 23664 42177 23673 42211
rect 23673 42177 23707 42211
rect 23707 42177 23716 42211
rect 23664 42168 23716 42177
rect 21916 42032 21968 42084
rect 22376 42032 22428 42084
rect 23020 42032 23072 42084
rect 24216 42100 24268 42152
rect 23940 42032 23992 42084
rect 24676 42168 24728 42220
rect 25044 42211 25096 42220
rect 25044 42177 25053 42211
rect 25053 42177 25087 42211
rect 25087 42177 25096 42211
rect 27804 42236 27856 42288
rect 28632 42279 28684 42288
rect 28632 42245 28641 42279
rect 28641 42245 28675 42279
rect 28675 42245 28684 42279
rect 28632 42236 28684 42245
rect 29644 42304 29696 42356
rect 25044 42168 25096 42177
rect 25688 42168 25740 42220
rect 25872 42211 25924 42220
rect 25872 42177 25881 42211
rect 25881 42177 25915 42211
rect 25915 42177 25924 42211
rect 25872 42168 25924 42177
rect 26240 42168 26292 42220
rect 28080 42168 28132 42220
rect 26332 42100 26384 42152
rect 28816 42168 28868 42220
rect 30012 42236 30064 42288
rect 30748 42236 30800 42288
rect 31852 42304 31904 42356
rect 33140 42304 33192 42356
rect 29092 42211 29144 42220
rect 29092 42177 29101 42211
rect 29101 42177 29135 42211
rect 29135 42177 29144 42211
rect 29092 42168 29144 42177
rect 29460 42168 29512 42220
rect 30288 42168 30340 42220
rect 30472 42211 30524 42220
rect 30472 42177 30481 42211
rect 30481 42177 30515 42211
rect 30515 42177 30524 42211
rect 30656 42211 30708 42220
rect 30472 42168 30524 42177
rect 30656 42177 30665 42211
rect 30665 42177 30699 42211
rect 30699 42177 30708 42211
rect 30656 42168 30708 42177
rect 31576 42211 31628 42220
rect 31576 42177 31600 42211
rect 31600 42177 31628 42211
rect 31576 42168 31628 42177
rect 32312 42236 32364 42288
rect 31944 42168 31996 42220
rect 32680 42168 32732 42220
rect 33692 42236 33744 42288
rect 33048 42168 33100 42220
rect 34796 42168 34848 42220
rect 34704 42100 34756 42152
rect 24492 42032 24544 42084
rect 25044 42032 25096 42084
rect 20076 41964 20128 42016
rect 21272 41964 21324 42016
rect 21824 41964 21876 42016
rect 24584 42007 24636 42016
rect 24584 41973 24593 42007
rect 24593 41973 24627 42007
rect 24627 41973 24636 42007
rect 24584 41964 24636 41973
rect 25320 41964 25372 42016
rect 25688 42007 25740 42016
rect 25688 41973 25697 42007
rect 25697 41973 25731 42007
rect 25731 41973 25740 42007
rect 25688 41964 25740 41973
rect 26976 42032 27028 42084
rect 29460 42032 29512 42084
rect 26608 42007 26660 42016
rect 26608 41973 26617 42007
rect 26617 41973 26651 42007
rect 26651 41973 26660 42007
rect 26608 41964 26660 41973
rect 26884 41964 26936 42016
rect 27988 41964 28040 42016
rect 30748 41964 30800 42016
rect 32036 41964 32088 42016
rect 32588 41964 32640 42016
rect 33968 41964 34020 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 21456 41760 21508 41812
rect 23664 41803 23716 41812
rect 21548 41692 21600 41744
rect 22192 41692 22244 41744
rect 20352 41624 20404 41676
rect 21916 41599 21968 41608
rect 21916 41565 21925 41599
rect 21925 41565 21959 41599
rect 21959 41565 21968 41599
rect 23664 41769 23673 41803
rect 23673 41769 23707 41803
rect 23707 41769 23716 41803
rect 23664 41760 23716 41769
rect 23756 41760 23808 41812
rect 26976 41760 27028 41812
rect 30656 41803 30708 41812
rect 30656 41769 30665 41803
rect 30665 41769 30699 41803
rect 30699 41769 30708 41803
rect 30656 41760 30708 41769
rect 31208 41760 31260 41812
rect 33600 41760 33652 41812
rect 34704 41760 34756 41812
rect 31300 41692 31352 41744
rect 31944 41692 31996 41744
rect 32588 41692 32640 41744
rect 21916 41556 21968 41565
rect 22468 41556 22520 41608
rect 24584 41624 24636 41676
rect 22744 41488 22796 41540
rect 25044 41556 25096 41608
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 25596 41599 25648 41608
rect 25596 41565 25605 41599
rect 25605 41565 25639 41599
rect 25639 41565 25648 41599
rect 25596 41556 25648 41565
rect 25872 41556 25924 41608
rect 27068 41599 27120 41608
rect 20444 41420 20496 41472
rect 20904 41420 20956 41472
rect 21916 41463 21968 41472
rect 21916 41429 21925 41463
rect 21925 41429 21959 41463
rect 21959 41429 21968 41463
rect 21916 41420 21968 41429
rect 24308 41488 24360 41540
rect 26148 41488 26200 41540
rect 27068 41565 27077 41599
rect 27077 41565 27111 41599
rect 27111 41565 27120 41599
rect 27068 41556 27120 41565
rect 27896 41624 27948 41676
rect 27344 41556 27396 41608
rect 27436 41599 27488 41608
rect 27436 41565 27445 41599
rect 27445 41565 27479 41599
rect 27479 41565 27488 41599
rect 27436 41556 27488 41565
rect 27620 41556 27672 41608
rect 29276 41624 29328 41676
rect 29552 41556 29604 41608
rect 29736 41599 29788 41608
rect 29736 41565 29745 41599
rect 29745 41565 29779 41599
rect 29779 41565 29788 41599
rect 29736 41556 29788 41565
rect 29920 41599 29972 41608
rect 29920 41565 29929 41599
rect 29929 41565 29963 41599
rect 29963 41565 29972 41599
rect 29920 41556 29972 41565
rect 30748 41599 30800 41608
rect 30748 41565 30757 41599
rect 30757 41565 30791 41599
rect 30791 41565 30800 41599
rect 30748 41556 30800 41565
rect 30932 41556 30984 41608
rect 31392 41556 31444 41608
rect 31576 41599 31628 41608
rect 31576 41565 31585 41599
rect 31585 41565 31619 41599
rect 31619 41565 31628 41599
rect 31576 41556 31628 41565
rect 35348 41692 35400 41744
rect 33048 41624 33100 41676
rect 33600 41599 33652 41608
rect 28816 41531 28868 41540
rect 28816 41497 28825 41531
rect 28825 41497 28859 41531
rect 28859 41497 28868 41531
rect 28816 41488 28868 41497
rect 25136 41463 25188 41472
rect 25136 41429 25145 41463
rect 25145 41429 25179 41463
rect 25179 41429 25188 41463
rect 25136 41420 25188 41429
rect 26516 41420 26568 41472
rect 26608 41420 26660 41472
rect 28080 41420 28132 41472
rect 28724 41420 28776 41472
rect 33600 41565 33609 41599
rect 33609 41565 33643 41599
rect 33643 41565 33652 41599
rect 33600 41556 33652 41565
rect 34796 41556 34848 41608
rect 35900 41556 35952 41608
rect 33784 41531 33836 41540
rect 30012 41420 30064 41472
rect 32772 41420 32824 41472
rect 33784 41497 33793 41531
rect 33793 41497 33827 41531
rect 33827 41497 33836 41531
rect 33784 41488 33836 41497
rect 33692 41420 33744 41472
rect 35164 41463 35216 41472
rect 35164 41429 35173 41463
rect 35173 41429 35207 41463
rect 35207 41429 35216 41463
rect 35164 41420 35216 41429
rect 35716 41463 35768 41472
rect 35716 41429 35725 41463
rect 35725 41429 35759 41463
rect 35759 41429 35768 41463
rect 35716 41420 35768 41429
rect 37464 41420 37516 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 21180 41216 21232 41268
rect 24768 41216 24820 41268
rect 25596 41216 25648 41268
rect 26240 41259 26292 41268
rect 26240 41225 26249 41259
rect 26249 41225 26283 41259
rect 26283 41225 26292 41259
rect 26240 41216 26292 41225
rect 26976 41216 27028 41268
rect 19340 41123 19392 41132
rect 19340 41089 19349 41123
rect 19349 41089 19383 41123
rect 19383 41089 19392 41123
rect 20628 41148 20680 41200
rect 23388 41191 23440 41200
rect 23388 41157 23397 41191
rect 23397 41157 23431 41191
rect 23431 41157 23440 41191
rect 23388 41148 23440 41157
rect 24492 41148 24544 41200
rect 20076 41123 20128 41132
rect 19340 41080 19392 41089
rect 20076 41089 20085 41123
rect 20085 41089 20119 41123
rect 20119 41089 20128 41123
rect 20076 41080 20128 41089
rect 21088 41123 21140 41132
rect 21088 41089 21097 41123
rect 21097 41089 21131 41123
rect 21131 41089 21140 41123
rect 21088 41080 21140 41089
rect 21456 41080 21508 41132
rect 22192 41123 22244 41132
rect 22192 41089 22201 41123
rect 22201 41089 22235 41123
rect 22235 41089 22244 41123
rect 22192 41080 22244 41089
rect 22468 41123 22520 41132
rect 22468 41089 22477 41123
rect 22477 41089 22511 41123
rect 22511 41089 22520 41123
rect 22468 41080 22520 41089
rect 23296 41080 23348 41132
rect 24860 41080 24912 41132
rect 25136 41123 25188 41132
rect 20720 41012 20772 41064
rect 21824 41012 21876 41064
rect 18696 40919 18748 40928
rect 18696 40885 18705 40919
rect 18705 40885 18739 40919
rect 18739 40885 18748 40919
rect 18696 40876 18748 40885
rect 20628 40876 20680 40928
rect 21364 40944 21416 40996
rect 21548 40944 21600 40996
rect 22928 41012 22980 41064
rect 23112 41012 23164 41064
rect 23940 41012 23992 41064
rect 24308 41055 24360 41064
rect 24308 41021 24317 41055
rect 24317 41021 24351 41055
rect 24351 41021 24360 41055
rect 24308 41012 24360 41021
rect 25136 41089 25145 41123
rect 25145 41089 25179 41123
rect 25179 41089 25188 41123
rect 25136 41080 25188 41089
rect 26148 41148 26200 41200
rect 25688 41123 25740 41132
rect 25688 41089 25697 41123
rect 25697 41089 25731 41123
rect 25731 41089 25740 41123
rect 25688 41080 25740 41089
rect 26516 41148 26568 41200
rect 27344 41148 27396 41200
rect 27804 41216 27856 41268
rect 28816 41216 28868 41268
rect 31024 41216 31076 41268
rect 31484 41259 31536 41268
rect 31484 41225 31493 41259
rect 31493 41225 31527 41259
rect 31527 41225 31536 41259
rect 31484 41216 31536 41225
rect 31760 41216 31812 41268
rect 32128 41216 32180 41268
rect 33784 41216 33836 41268
rect 27620 41080 27672 41132
rect 29276 41080 29328 41132
rect 29920 41148 29972 41200
rect 32680 41148 32732 41200
rect 30104 41080 30156 41132
rect 32220 41080 32272 41132
rect 33600 41148 33652 41200
rect 33140 41080 33192 41132
rect 33692 41123 33744 41132
rect 33692 41089 33701 41123
rect 33701 41089 33735 41123
rect 33735 41089 33744 41123
rect 33692 41080 33744 41089
rect 33968 41123 34020 41132
rect 27160 41012 27212 41064
rect 27344 41012 27396 41064
rect 32588 41012 32640 41064
rect 33968 41089 33977 41123
rect 33977 41089 34011 41123
rect 34011 41089 34020 41123
rect 33968 41080 34020 41089
rect 25320 40987 25372 40996
rect 25320 40953 25329 40987
rect 25329 40953 25363 40987
rect 25363 40953 25372 40987
rect 25320 40944 25372 40953
rect 28080 40944 28132 40996
rect 29920 40944 29972 40996
rect 30932 40944 30984 40996
rect 32128 40944 32180 40996
rect 33048 40944 33100 40996
rect 35164 41012 35216 41064
rect 33784 40944 33836 40996
rect 22928 40876 22980 40928
rect 23480 40876 23532 40928
rect 26424 40919 26476 40928
rect 26424 40885 26433 40919
rect 26433 40885 26467 40919
rect 26467 40885 26476 40919
rect 26424 40876 26476 40885
rect 27068 40876 27120 40928
rect 27804 40876 27856 40928
rect 28816 40876 28868 40928
rect 30288 40876 30340 40928
rect 30380 40876 30432 40928
rect 32312 40876 32364 40928
rect 32680 40919 32732 40928
rect 32680 40885 32689 40919
rect 32689 40885 32723 40919
rect 32723 40885 32732 40919
rect 32680 40876 32732 40885
rect 33232 40876 33284 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 20260 40672 20312 40724
rect 21640 40672 21692 40724
rect 23940 40672 23992 40724
rect 24308 40672 24360 40724
rect 26240 40672 26292 40724
rect 26608 40672 26660 40724
rect 27252 40672 27304 40724
rect 28172 40672 28224 40724
rect 31944 40672 31996 40724
rect 32312 40672 32364 40724
rect 25688 40604 25740 40656
rect 26516 40604 26568 40656
rect 19432 40536 19484 40588
rect 21180 40536 21232 40588
rect 1952 40468 2004 40520
rect 18328 40511 18380 40520
rect 18328 40477 18337 40511
rect 18337 40477 18371 40511
rect 18371 40477 18380 40511
rect 18328 40468 18380 40477
rect 21732 40511 21784 40520
rect 18880 40400 18932 40452
rect 21732 40477 21741 40511
rect 21741 40477 21775 40511
rect 21775 40477 21784 40511
rect 21732 40468 21784 40477
rect 22284 40468 22336 40520
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 27068 40579 27120 40588
rect 27068 40545 27077 40579
rect 27077 40545 27111 40579
rect 27111 40545 27120 40579
rect 27068 40536 27120 40545
rect 30564 40604 30616 40656
rect 27344 40579 27396 40588
rect 27344 40545 27353 40579
rect 27353 40545 27387 40579
rect 27387 40545 27396 40579
rect 33692 40604 33744 40656
rect 27344 40536 27396 40545
rect 22836 40400 22888 40452
rect 23664 40468 23716 40520
rect 24032 40468 24084 40520
rect 24216 40468 24268 40520
rect 24768 40511 24820 40520
rect 1676 40375 1728 40384
rect 1676 40341 1685 40375
rect 1685 40341 1719 40375
rect 1719 40341 1728 40375
rect 1676 40332 1728 40341
rect 18512 40375 18564 40384
rect 18512 40341 18521 40375
rect 18521 40341 18555 40375
rect 18555 40341 18564 40375
rect 18512 40332 18564 40341
rect 18788 40332 18840 40384
rect 19984 40332 20036 40384
rect 21088 40375 21140 40384
rect 21088 40341 21097 40375
rect 21097 40341 21131 40375
rect 21131 40341 21140 40375
rect 21088 40332 21140 40341
rect 21180 40332 21232 40384
rect 21732 40332 21784 40384
rect 23020 40332 23072 40384
rect 23388 40400 23440 40452
rect 24768 40477 24777 40511
rect 24777 40477 24811 40511
rect 24811 40477 24820 40511
rect 24768 40468 24820 40477
rect 27160 40511 27212 40520
rect 27160 40477 27169 40511
rect 27169 40477 27203 40511
rect 27203 40477 27212 40511
rect 27160 40468 27212 40477
rect 24584 40332 24636 40384
rect 25780 40400 25832 40452
rect 25964 40400 26016 40452
rect 27712 40468 27764 40520
rect 28540 40443 28592 40452
rect 28540 40409 28549 40443
rect 28549 40409 28583 40443
rect 28583 40409 28592 40443
rect 28540 40400 28592 40409
rect 28724 40468 28776 40520
rect 29920 40468 29972 40520
rect 31024 40536 31076 40588
rect 31944 40536 31996 40588
rect 32036 40511 32088 40520
rect 32036 40477 32045 40511
rect 32045 40477 32079 40511
rect 32079 40477 32088 40511
rect 32036 40468 32088 40477
rect 32404 40468 32456 40520
rect 32496 40468 32548 40520
rect 33416 40511 33468 40520
rect 25504 40332 25556 40384
rect 27160 40332 27212 40384
rect 27436 40332 27488 40384
rect 29184 40332 29236 40384
rect 30288 40375 30340 40384
rect 30288 40341 30297 40375
rect 30297 40341 30331 40375
rect 30331 40341 30340 40375
rect 30288 40332 30340 40341
rect 30564 40332 30616 40384
rect 31300 40332 31352 40384
rect 32496 40332 32548 40384
rect 33416 40477 33425 40511
rect 33425 40477 33459 40511
rect 33459 40477 33468 40511
rect 33416 40468 33468 40477
rect 35348 40468 35400 40520
rect 33324 40375 33376 40384
rect 33324 40341 33333 40375
rect 33333 40341 33367 40375
rect 33367 40341 33376 40375
rect 33324 40332 33376 40341
rect 35808 40332 35860 40384
rect 35900 40332 35952 40384
rect 57704 40332 57756 40384
rect 58256 40375 58308 40384
rect 58256 40341 58265 40375
rect 58265 40341 58299 40375
rect 58299 40341 58308 40375
rect 58256 40332 58308 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 19892 40171 19944 40180
rect 19892 40137 19894 40171
rect 19894 40137 19928 40171
rect 19928 40137 19944 40171
rect 19892 40128 19944 40137
rect 22100 40128 22152 40180
rect 17776 40035 17828 40044
rect 17776 40001 17785 40035
rect 17785 40001 17819 40035
rect 17819 40001 17828 40035
rect 17776 39992 17828 40001
rect 17960 40035 18012 40044
rect 17960 40001 17969 40035
rect 17969 40001 18003 40035
rect 18003 40001 18012 40035
rect 17960 39992 18012 40001
rect 18328 39992 18380 40044
rect 18880 39992 18932 40044
rect 19340 39992 19392 40044
rect 20168 40060 20220 40112
rect 20904 40035 20956 40044
rect 20904 40001 20913 40035
rect 20913 40001 20947 40035
rect 20947 40001 20956 40035
rect 20904 39992 20956 40001
rect 22100 39992 22152 40044
rect 22284 39992 22336 40044
rect 23388 40103 23440 40112
rect 23388 40069 23397 40103
rect 23397 40069 23431 40103
rect 23431 40069 23440 40103
rect 23388 40060 23440 40069
rect 22928 39992 22980 40044
rect 23480 40035 23532 40044
rect 23480 40001 23489 40035
rect 23489 40001 23523 40035
rect 23523 40001 23532 40035
rect 27160 40060 27212 40112
rect 27344 40128 27396 40180
rect 27620 40060 27672 40112
rect 27988 40060 28040 40112
rect 28540 40060 28592 40112
rect 28724 40060 28776 40112
rect 30288 40128 30340 40180
rect 32220 40128 32272 40180
rect 32496 40128 32548 40180
rect 24124 40035 24176 40044
rect 23480 39992 23532 40001
rect 24124 40001 24133 40035
rect 24133 40001 24167 40035
rect 24167 40001 24176 40035
rect 24124 39992 24176 40001
rect 24768 39992 24820 40044
rect 25872 39992 25924 40044
rect 26240 39992 26292 40044
rect 27068 39992 27120 40044
rect 23388 39924 23440 39976
rect 24400 39967 24452 39976
rect 24400 39933 24409 39967
rect 24409 39933 24443 39967
rect 24443 39933 24452 39967
rect 24400 39924 24452 39933
rect 25136 39967 25188 39976
rect 25136 39933 25145 39967
rect 25145 39933 25179 39967
rect 25179 39933 25188 39967
rect 25136 39924 25188 39933
rect 19432 39856 19484 39908
rect 22100 39856 22152 39908
rect 23480 39856 23532 39908
rect 25044 39856 25096 39908
rect 25688 39924 25740 39976
rect 26976 39924 27028 39976
rect 28816 40035 28868 40044
rect 28816 40001 28825 40035
rect 28825 40001 28859 40035
rect 28859 40001 28868 40035
rect 28816 39992 28868 40001
rect 27344 39967 27396 39976
rect 27344 39933 27353 39967
rect 27353 39933 27387 39967
rect 27387 39933 27396 39967
rect 27344 39924 27396 39933
rect 27436 39967 27488 39976
rect 27436 39933 27445 39967
rect 27445 39933 27479 39967
rect 27479 39933 27488 39967
rect 27436 39924 27488 39933
rect 27620 39967 27672 39976
rect 27620 39933 27629 39967
rect 27629 39933 27663 39967
rect 27663 39933 27672 39967
rect 27620 39924 27672 39933
rect 27804 39924 27856 39976
rect 27988 39924 28040 39976
rect 32128 40060 32180 40112
rect 29000 40035 29052 40044
rect 29000 40001 29009 40035
rect 29009 40001 29043 40035
rect 29043 40001 29052 40035
rect 29184 40035 29236 40044
rect 29000 39992 29052 40001
rect 29184 40001 29193 40035
rect 29193 40001 29227 40035
rect 29227 40001 29236 40035
rect 29184 39992 29236 40001
rect 29736 39924 29788 39976
rect 31484 39992 31536 40044
rect 31760 39992 31812 40044
rect 33324 40060 33376 40112
rect 35440 40128 35492 40180
rect 35716 40060 35768 40112
rect 18604 39788 18656 39840
rect 20996 39788 21048 39840
rect 21824 39788 21876 39840
rect 22376 39831 22428 39840
rect 22376 39797 22385 39831
rect 22385 39797 22419 39831
rect 22419 39797 22428 39831
rect 22376 39788 22428 39797
rect 22468 39788 22520 39840
rect 23940 39831 23992 39840
rect 23940 39797 23949 39831
rect 23949 39797 23983 39831
rect 23983 39797 23992 39831
rect 23940 39788 23992 39797
rect 24952 39788 25004 39840
rect 27436 39788 27488 39840
rect 27528 39788 27580 39840
rect 28632 39831 28684 39840
rect 28632 39797 28641 39831
rect 28641 39797 28675 39831
rect 28675 39797 28684 39831
rect 32128 39924 32180 39976
rect 35808 39992 35860 40044
rect 33876 39967 33928 39976
rect 33508 39856 33560 39908
rect 28632 39788 28684 39797
rect 29552 39788 29604 39840
rect 30012 39831 30064 39840
rect 30012 39797 30021 39831
rect 30021 39797 30055 39831
rect 30055 39797 30064 39831
rect 30012 39788 30064 39797
rect 30104 39788 30156 39840
rect 31576 39788 31628 39840
rect 32220 39788 32272 39840
rect 33876 39933 33885 39967
rect 33885 39933 33919 39967
rect 33919 39933 33928 39967
rect 33876 39924 33928 39933
rect 35900 39967 35952 39976
rect 35900 39933 35909 39967
rect 35909 39933 35943 39967
rect 35943 39933 35952 39967
rect 35900 39924 35952 39933
rect 35716 39788 35768 39840
rect 36084 39788 36136 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 18512 39627 18564 39636
rect 18512 39593 18521 39627
rect 18521 39593 18555 39627
rect 18555 39593 18564 39627
rect 18512 39584 18564 39593
rect 18696 39584 18748 39636
rect 23388 39584 23440 39636
rect 26056 39584 26108 39636
rect 27344 39584 27396 39636
rect 27620 39584 27672 39636
rect 20904 39516 20956 39568
rect 20352 39448 20404 39500
rect 21640 39516 21692 39568
rect 21824 39516 21876 39568
rect 25136 39559 25188 39568
rect 20168 39423 20220 39432
rect 18604 39312 18656 39364
rect 20168 39389 20177 39423
rect 20177 39389 20211 39423
rect 20211 39389 20220 39423
rect 20168 39380 20220 39389
rect 20260 39423 20312 39432
rect 20260 39389 20269 39423
rect 20269 39389 20303 39423
rect 20303 39389 20312 39423
rect 22100 39448 22152 39500
rect 20260 39380 20312 39389
rect 21180 39380 21232 39432
rect 21364 39423 21416 39432
rect 21364 39389 21373 39423
rect 21373 39389 21407 39423
rect 21407 39389 21416 39423
rect 21364 39380 21416 39389
rect 21548 39380 21600 39432
rect 16580 39244 16632 39296
rect 17316 39287 17368 39296
rect 17316 39253 17325 39287
rect 17325 39253 17359 39287
rect 17359 39253 17368 39287
rect 17316 39244 17368 39253
rect 18052 39244 18104 39296
rect 20720 39244 20772 39296
rect 21456 39244 21508 39296
rect 22744 39423 22796 39432
rect 22744 39389 22753 39423
rect 22753 39389 22787 39423
rect 22787 39389 22796 39423
rect 22744 39380 22796 39389
rect 22928 39423 22980 39432
rect 22928 39389 22937 39423
rect 22937 39389 22971 39423
rect 22971 39389 22980 39423
rect 22928 39380 22980 39389
rect 23388 39380 23440 39432
rect 24860 39423 24912 39432
rect 24860 39389 24869 39423
rect 24869 39389 24903 39423
rect 24903 39389 24912 39423
rect 24860 39380 24912 39389
rect 25136 39525 25145 39559
rect 25145 39525 25179 39559
rect 25179 39525 25188 39559
rect 25136 39516 25188 39525
rect 28356 39584 28408 39636
rect 28816 39584 28868 39636
rect 30564 39584 30616 39636
rect 30932 39584 30984 39636
rect 32128 39584 32180 39636
rect 28172 39516 28224 39568
rect 29828 39516 29880 39568
rect 32496 39516 32548 39568
rect 27068 39448 27120 39500
rect 23848 39312 23900 39364
rect 25228 39380 25280 39432
rect 26148 39423 26200 39432
rect 26148 39389 26157 39423
rect 26157 39389 26191 39423
rect 26191 39389 26200 39423
rect 26148 39380 26200 39389
rect 25412 39312 25464 39364
rect 25688 39312 25740 39364
rect 22836 39244 22888 39296
rect 23388 39287 23440 39296
rect 23388 39253 23397 39287
rect 23397 39253 23431 39287
rect 23431 39253 23440 39287
rect 23388 39244 23440 39253
rect 23756 39244 23808 39296
rect 24032 39244 24084 39296
rect 26516 39312 26568 39364
rect 27620 39380 27672 39432
rect 28172 39380 28224 39432
rect 30288 39448 30340 39500
rect 30932 39448 30984 39500
rect 32772 39491 32824 39500
rect 32772 39457 32781 39491
rect 32781 39457 32815 39491
rect 32815 39457 32824 39491
rect 32772 39448 32824 39457
rect 32956 39516 33008 39568
rect 35440 39448 35492 39500
rect 35716 39491 35768 39500
rect 35716 39457 35725 39491
rect 35725 39457 35759 39491
rect 35759 39457 35768 39491
rect 35716 39448 35768 39457
rect 35900 39448 35952 39500
rect 36084 39491 36136 39500
rect 36084 39457 36093 39491
rect 36093 39457 36127 39491
rect 36127 39457 36136 39491
rect 36084 39448 36136 39457
rect 37464 39491 37516 39500
rect 37464 39457 37473 39491
rect 37473 39457 37507 39491
rect 37507 39457 37516 39491
rect 37464 39448 37516 39457
rect 29092 39423 29144 39432
rect 29092 39389 29100 39423
rect 29100 39389 29134 39423
rect 29134 39389 29144 39423
rect 29092 39380 29144 39389
rect 29276 39380 29328 39432
rect 29736 39423 29788 39432
rect 29736 39389 29745 39423
rect 29745 39389 29779 39423
rect 29779 39389 29788 39423
rect 29736 39380 29788 39389
rect 29828 39380 29880 39432
rect 30380 39380 30432 39432
rect 30104 39355 30156 39364
rect 30104 39321 30113 39355
rect 30113 39321 30147 39355
rect 30147 39321 30156 39355
rect 31208 39380 31260 39432
rect 32496 39380 32548 39432
rect 33508 39380 33560 39432
rect 34060 39380 34112 39432
rect 30104 39312 30156 39321
rect 26700 39287 26752 39296
rect 26700 39253 26709 39287
rect 26709 39253 26743 39287
rect 26743 39253 26752 39287
rect 26700 39244 26752 39253
rect 26792 39244 26844 39296
rect 26976 39244 27028 39296
rect 27712 39244 27764 39296
rect 27804 39244 27856 39296
rect 29092 39244 29144 39296
rect 32864 39312 32916 39364
rect 32128 39287 32180 39296
rect 32128 39253 32137 39287
rect 32137 39253 32171 39287
rect 32171 39253 32180 39287
rect 32128 39244 32180 39253
rect 32496 39244 32548 39296
rect 34520 39312 34572 39364
rect 33692 39287 33744 39296
rect 33692 39253 33701 39287
rect 33701 39253 33735 39287
rect 33735 39253 33744 39287
rect 33692 39244 33744 39253
rect 34244 39287 34296 39296
rect 34244 39253 34253 39287
rect 34253 39253 34287 39287
rect 34287 39253 34296 39287
rect 34244 39244 34296 39253
rect 35808 39244 35860 39296
rect 36176 39244 36228 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 17960 39040 18012 39092
rect 18512 39040 18564 39092
rect 18696 39083 18748 39092
rect 18696 39049 18705 39083
rect 18705 39049 18739 39083
rect 18739 39049 18748 39083
rect 18696 39040 18748 39049
rect 20168 39040 20220 39092
rect 16580 38904 16632 38956
rect 17040 38947 17092 38956
rect 17040 38913 17068 38947
rect 17068 38913 17092 38947
rect 17224 38947 17276 38956
rect 17040 38904 17092 38913
rect 17224 38913 17233 38947
rect 17233 38913 17267 38947
rect 17267 38913 17276 38947
rect 17224 38904 17276 38913
rect 20444 39040 20496 39092
rect 22100 39040 22152 39092
rect 20812 38972 20864 39024
rect 21180 38972 21232 39024
rect 21640 38972 21692 39024
rect 17132 38768 17184 38820
rect 16580 38700 16632 38752
rect 17040 38700 17092 38752
rect 22008 38904 22060 38956
rect 20720 38879 20772 38888
rect 20720 38845 20729 38879
rect 20729 38845 20763 38879
rect 20763 38845 20772 38879
rect 20720 38836 20772 38845
rect 22468 38904 22520 38956
rect 23296 38972 23348 39024
rect 23388 38972 23440 39024
rect 23480 38947 23532 38956
rect 23480 38913 23489 38947
rect 23489 38913 23523 38947
rect 23523 38913 23532 38947
rect 23480 38904 23532 38913
rect 23388 38836 23440 38888
rect 20444 38768 20496 38820
rect 17868 38700 17920 38752
rect 22008 38743 22060 38752
rect 22008 38709 22017 38743
rect 22017 38709 22051 38743
rect 22051 38709 22060 38743
rect 22008 38700 22060 38709
rect 22192 38768 22244 38820
rect 23664 38836 23716 38888
rect 23664 38700 23716 38752
rect 24032 38904 24084 38956
rect 24492 39040 24544 39092
rect 26332 39040 26384 39092
rect 26792 39040 26844 39092
rect 27436 39040 27488 39092
rect 27620 39040 27672 39092
rect 30196 39040 30248 39092
rect 30380 39040 30432 39092
rect 30472 39040 30524 39092
rect 26700 38972 26752 39024
rect 27344 38972 27396 39024
rect 27804 38972 27856 39024
rect 25136 38836 25188 38888
rect 26884 38904 26936 38956
rect 27436 38947 27488 38956
rect 27436 38913 27445 38947
rect 27445 38913 27479 38947
rect 27479 38913 27488 38947
rect 27436 38904 27488 38913
rect 29000 38972 29052 39024
rect 29736 38972 29788 39024
rect 32956 39040 33008 39092
rect 33876 39083 33928 39092
rect 33876 39049 33885 39083
rect 33885 39049 33919 39083
rect 33919 39049 33928 39083
rect 33876 39040 33928 39049
rect 34520 39040 34572 39092
rect 28448 38947 28500 38956
rect 28448 38913 28457 38947
rect 28457 38913 28491 38947
rect 28491 38913 28500 38947
rect 28448 38904 28500 38913
rect 27160 38836 27212 38888
rect 27252 38836 27304 38888
rect 26148 38768 26200 38820
rect 27804 38836 27856 38888
rect 28356 38836 28408 38888
rect 29184 38904 29236 38956
rect 29644 38904 29696 38956
rect 29920 38904 29972 38956
rect 30196 38947 30248 38956
rect 30196 38913 30205 38947
rect 30205 38913 30239 38947
rect 30239 38913 30248 38947
rect 30196 38904 30248 38913
rect 30288 38947 30340 38956
rect 30288 38913 30297 38947
rect 30297 38913 30331 38947
rect 30331 38913 30340 38947
rect 30288 38904 30340 38913
rect 31300 38947 31352 38956
rect 29828 38836 29880 38888
rect 27712 38768 27764 38820
rect 24124 38743 24176 38752
rect 24124 38709 24133 38743
rect 24133 38709 24167 38743
rect 24167 38709 24176 38743
rect 24124 38700 24176 38709
rect 26056 38743 26108 38752
rect 26056 38709 26065 38743
rect 26065 38709 26099 38743
rect 26099 38709 26108 38743
rect 26056 38700 26108 38709
rect 26608 38700 26660 38752
rect 27160 38743 27212 38752
rect 27160 38709 27169 38743
rect 27169 38709 27203 38743
rect 27203 38709 27212 38743
rect 27160 38700 27212 38709
rect 27344 38700 27396 38752
rect 27620 38700 27672 38752
rect 29736 38768 29788 38820
rect 31300 38913 31309 38947
rect 31309 38913 31343 38947
rect 31343 38913 31352 38947
rect 31300 38904 31352 38913
rect 32404 38972 32456 39024
rect 32128 38904 32180 38956
rect 32588 38947 32640 38956
rect 32588 38913 32597 38947
rect 32597 38913 32631 38947
rect 32631 38913 32640 38947
rect 32588 38904 32640 38913
rect 33140 38904 33192 38956
rect 27988 38700 28040 38752
rect 28632 38700 28684 38752
rect 29460 38743 29512 38752
rect 29460 38709 29469 38743
rect 29469 38709 29503 38743
rect 29503 38709 29512 38743
rect 29460 38700 29512 38709
rect 29644 38700 29696 38752
rect 30012 38700 30064 38752
rect 31944 38768 31996 38820
rect 36360 38972 36412 39024
rect 34520 38904 34572 38956
rect 34796 38904 34848 38956
rect 33600 38836 33652 38888
rect 34060 38879 34112 38888
rect 34060 38845 34069 38879
rect 34069 38845 34103 38879
rect 34103 38845 34112 38879
rect 34060 38836 34112 38845
rect 34244 38879 34296 38888
rect 34244 38845 34253 38879
rect 34253 38845 34287 38879
rect 34287 38845 34296 38879
rect 34244 38836 34296 38845
rect 34336 38879 34388 38888
rect 34336 38845 34345 38879
rect 34345 38845 34379 38879
rect 34379 38845 34388 38879
rect 34336 38836 34388 38845
rect 34612 38836 34664 38888
rect 35072 38836 35124 38888
rect 30656 38700 30708 38752
rect 31116 38743 31168 38752
rect 31116 38709 31125 38743
rect 31125 38709 31159 38743
rect 31159 38709 31168 38743
rect 31116 38700 31168 38709
rect 34428 38768 34480 38820
rect 35348 38836 35400 38888
rect 34520 38700 34572 38752
rect 34704 38700 34756 38752
rect 35072 38743 35124 38752
rect 35072 38709 35081 38743
rect 35081 38709 35115 38743
rect 35115 38709 35124 38743
rect 35072 38700 35124 38709
rect 36176 38700 36228 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 17132 38496 17184 38548
rect 18512 38539 18564 38548
rect 18512 38505 18521 38539
rect 18521 38505 18555 38539
rect 18555 38505 18564 38539
rect 18512 38496 18564 38505
rect 18604 38496 18656 38548
rect 17868 38428 17920 38480
rect 20812 38496 20864 38548
rect 22744 38496 22796 38548
rect 16580 38403 16632 38412
rect 16580 38369 16589 38403
rect 16589 38369 16623 38403
rect 16623 38369 16632 38403
rect 16580 38360 16632 38369
rect 19248 38360 19300 38412
rect 17224 38292 17276 38344
rect 17684 38292 17736 38344
rect 17868 38335 17920 38344
rect 17868 38301 17877 38335
rect 17877 38301 17911 38335
rect 17911 38301 17920 38335
rect 17868 38292 17920 38301
rect 19984 38403 20036 38412
rect 19984 38369 19993 38403
rect 19993 38369 20027 38403
rect 20027 38369 20036 38403
rect 19984 38360 20036 38369
rect 20536 38335 20588 38344
rect 17040 38224 17092 38276
rect 18696 38267 18748 38276
rect 18696 38233 18705 38267
rect 18705 38233 18739 38267
rect 18739 38233 18748 38267
rect 20536 38301 20545 38335
rect 20545 38301 20579 38335
rect 20579 38301 20588 38335
rect 20536 38292 20588 38301
rect 21180 38292 21232 38344
rect 21548 38360 21600 38412
rect 22468 38360 22520 38412
rect 18696 38224 18748 38233
rect 16304 38156 16356 38208
rect 16396 38156 16448 38208
rect 17776 38156 17828 38208
rect 20536 38156 20588 38208
rect 21916 38156 21968 38208
rect 22284 38335 22336 38344
rect 22284 38301 22293 38335
rect 22293 38301 22327 38335
rect 22327 38301 22336 38335
rect 23112 38360 23164 38412
rect 24124 38428 24176 38480
rect 25136 38428 25188 38480
rect 25964 38428 26016 38480
rect 26240 38360 26292 38412
rect 26608 38360 26660 38412
rect 22284 38292 22336 38301
rect 23572 38292 23624 38344
rect 24584 38335 24636 38344
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 26056 38335 26108 38344
rect 26056 38301 26065 38335
rect 26065 38301 26099 38335
rect 26099 38301 26108 38335
rect 26056 38292 26108 38301
rect 23296 38224 23348 38276
rect 26332 38292 26384 38344
rect 27068 38360 27120 38412
rect 27896 38428 27948 38480
rect 28908 38428 28960 38480
rect 28724 38360 28776 38412
rect 27436 38335 27488 38344
rect 22652 38156 22704 38208
rect 22928 38156 22980 38208
rect 23112 38156 23164 38208
rect 24032 38199 24084 38208
rect 24032 38165 24041 38199
rect 24041 38165 24075 38199
rect 24075 38165 24084 38199
rect 24032 38156 24084 38165
rect 25136 38156 25188 38208
rect 25596 38199 25648 38208
rect 25596 38165 25605 38199
rect 25605 38165 25639 38199
rect 25639 38165 25648 38199
rect 25596 38156 25648 38165
rect 26148 38156 26200 38208
rect 27436 38301 27445 38335
rect 27445 38301 27479 38335
rect 27479 38301 27488 38335
rect 27436 38292 27488 38301
rect 29092 38335 29144 38344
rect 29092 38301 29101 38335
rect 29101 38301 29135 38335
rect 29135 38301 29144 38335
rect 29092 38292 29144 38301
rect 30564 38496 30616 38548
rect 30196 38428 30248 38480
rect 32588 38496 32640 38548
rect 32864 38428 32916 38480
rect 32312 38403 32364 38412
rect 32312 38369 32321 38403
rect 32321 38369 32355 38403
rect 32355 38369 32364 38403
rect 32312 38360 32364 38369
rect 32588 38360 32640 38412
rect 34612 38496 34664 38548
rect 33324 38403 33376 38412
rect 33324 38369 33358 38403
rect 33358 38369 33376 38403
rect 33508 38403 33560 38412
rect 33324 38360 33376 38369
rect 33508 38369 33517 38403
rect 33517 38369 33551 38403
rect 33551 38369 33560 38403
rect 33508 38360 33560 38369
rect 35440 38360 35492 38412
rect 30380 38335 30432 38344
rect 30380 38301 30389 38335
rect 30389 38301 30423 38335
rect 30423 38301 30432 38335
rect 30380 38292 30432 38301
rect 30748 38292 30800 38344
rect 29000 38224 29052 38276
rect 29460 38224 29512 38276
rect 31300 38292 31352 38344
rect 31944 38292 31996 38344
rect 32496 38335 32548 38344
rect 32496 38301 32505 38335
rect 32505 38301 32539 38335
rect 32539 38301 32548 38335
rect 32496 38292 32548 38301
rect 35348 38224 35400 38276
rect 36176 38224 36228 38276
rect 37096 38224 37148 38276
rect 28816 38156 28868 38208
rect 29736 38199 29788 38208
rect 29736 38165 29745 38199
rect 29745 38165 29779 38199
rect 29779 38165 29788 38199
rect 29736 38156 29788 38165
rect 30012 38156 30064 38208
rect 31208 38156 31260 38208
rect 34152 38199 34204 38208
rect 34152 38165 34161 38199
rect 34161 38165 34195 38199
rect 34195 38165 34204 38199
rect 34152 38156 34204 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 17224 37952 17276 38004
rect 18696 37995 18748 38004
rect 18696 37961 18705 37995
rect 18705 37961 18739 37995
rect 18739 37961 18748 37995
rect 18696 37952 18748 37961
rect 20720 37952 20772 38004
rect 21088 37952 21140 38004
rect 17776 37884 17828 37936
rect 15568 37816 15620 37868
rect 16580 37816 16632 37868
rect 17960 37859 18012 37868
rect 17960 37825 17969 37859
rect 17969 37825 18003 37859
rect 18003 37825 18012 37859
rect 17960 37816 18012 37825
rect 18880 37816 18932 37868
rect 19800 37859 19852 37868
rect 19800 37825 19809 37859
rect 19809 37825 19843 37859
rect 19843 37825 19852 37859
rect 19800 37816 19852 37825
rect 22100 37884 22152 37936
rect 23480 37952 23532 38004
rect 31484 37995 31536 38004
rect 20904 37816 20956 37868
rect 21272 37816 21324 37868
rect 22560 37816 22612 37868
rect 24032 37884 24084 37936
rect 25412 37884 25464 37936
rect 26148 37927 26200 37936
rect 23756 37816 23808 37868
rect 24492 37816 24544 37868
rect 24676 37816 24728 37868
rect 26148 37893 26157 37927
rect 26157 37893 26191 37927
rect 26191 37893 26200 37927
rect 26148 37884 26200 37893
rect 27252 37816 27304 37868
rect 27804 37884 27856 37936
rect 28264 37884 28316 37936
rect 21732 37748 21784 37800
rect 21916 37748 21968 37800
rect 17684 37723 17736 37732
rect 17684 37689 17693 37723
rect 17693 37689 17727 37723
rect 17727 37689 17736 37723
rect 17684 37680 17736 37689
rect 16396 37612 16448 37664
rect 17224 37655 17276 37664
rect 17224 37621 17233 37655
rect 17233 37621 17267 37655
rect 17267 37621 17276 37655
rect 17224 37612 17276 37621
rect 22652 37748 22704 37800
rect 22284 37612 22336 37664
rect 22560 37655 22612 37664
rect 22560 37621 22569 37655
rect 22569 37621 22603 37655
rect 22603 37621 22612 37655
rect 22560 37612 22612 37621
rect 22652 37612 22704 37664
rect 23296 37680 23348 37732
rect 25228 37680 25280 37732
rect 25780 37680 25832 37732
rect 26148 37748 26200 37800
rect 27896 37748 27948 37800
rect 28448 37816 28500 37868
rect 28632 37816 28684 37868
rect 31484 37961 31493 37995
rect 31493 37961 31527 37995
rect 31527 37961 31536 37995
rect 31484 37952 31536 37961
rect 31944 37952 31996 38004
rect 34336 37952 34388 38004
rect 34704 37995 34756 38004
rect 34704 37961 34713 37995
rect 34713 37961 34747 37995
rect 34747 37961 34756 37995
rect 34704 37952 34756 37961
rect 35348 37995 35400 38004
rect 35348 37961 35357 37995
rect 35357 37961 35391 37995
rect 35391 37961 35400 37995
rect 35348 37952 35400 37961
rect 31668 37884 31720 37936
rect 29276 37816 29328 37868
rect 30472 37816 30524 37868
rect 31392 37816 31444 37868
rect 32496 37816 32548 37868
rect 33048 37816 33100 37868
rect 29460 37748 29512 37800
rect 28448 37680 28500 37732
rect 28724 37680 28776 37732
rect 29828 37723 29880 37732
rect 29828 37689 29837 37723
rect 29837 37689 29871 37723
rect 29871 37689 29880 37723
rect 29828 37680 29880 37689
rect 23664 37612 23716 37664
rect 24124 37612 24176 37664
rect 24216 37612 24268 37664
rect 25044 37612 25096 37664
rect 27804 37612 27856 37664
rect 28908 37655 28960 37664
rect 28908 37621 28917 37655
rect 28917 37621 28951 37655
rect 28951 37621 28960 37655
rect 28908 37612 28960 37621
rect 29184 37612 29236 37664
rect 33784 37748 33836 37800
rect 34704 37816 34756 37868
rect 32128 37680 32180 37732
rect 30380 37655 30432 37664
rect 30380 37621 30389 37655
rect 30389 37621 30423 37655
rect 30423 37621 30432 37655
rect 30380 37612 30432 37621
rect 31208 37612 31260 37664
rect 31392 37612 31444 37664
rect 31484 37612 31536 37664
rect 32036 37612 32088 37664
rect 33600 37612 33652 37664
rect 35992 37612 36044 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19800 37408 19852 37460
rect 20996 37408 21048 37460
rect 21088 37408 21140 37460
rect 23664 37408 23716 37460
rect 23848 37451 23900 37460
rect 23848 37417 23857 37451
rect 23857 37417 23891 37451
rect 23891 37417 23900 37451
rect 23848 37408 23900 37417
rect 24124 37408 24176 37460
rect 25504 37408 25556 37460
rect 25780 37408 25832 37460
rect 26148 37408 26200 37460
rect 26884 37408 26936 37460
rect 28356 37408 28408 37460
rect 30196 37408 30248 37460
rect 22100 37340 22152 37392
rect 23112 37340 23164 37392
rect 16580 37272 16632 37324
rect 17592 37272 17644 37324
rect 18880 37272 18932 37324
rect 21548 37272 21600 37324
rect 22192 37272 22244 37324
rect 15568 37247 15620 37256
rect 15568 37213 15577 37247
rect 15577 37213 15611 37247
rect 15611 37213 15620 37247
rect 15568 37204 15620 37213
rect 16396 37247 16448 37256
rect 15384 37179 15436 37188
rect 15384 37145 15393 37179
rect 15393 37145 15427 37179
rect 15427 37145 15436 37179
rect 16396 37213 16405 37247
rect 16405 37213 16439 37247
rect 16439 37213 16448 37247
rect 16396 37204 16448 37213
rect 17132 37204 17184 37256
rect 17224 37247 17276 37256
rect 17224 37213 17233 37247
rect 17233 37213 17267 37247
rect 17267 37213 17276 37247
rect 17224 37204 17276 37213
rect 15384 37136 15436 37145
rect 20168 37204 20220 37256
rect 21364 37204 21416 37256
rect 22008 37204 22060 37256
rect 22284 37204 22336 37256
rect 22468 37247 22520 37256
rect 22468 37213 22478 37247
rect 22478 37213 22512 37247
rect 22512 37213 22520 37247
rect 22468 37204 22520 37213
rect 21732 37136 21784 37188
rect 23388 37272 23440 37324
rect 23756 37315 23808 37324
rect 23756 37281 23765 37315
rect 23765 37281 23799 37315
rect 23799 37281 23808 37315
rect 23756 37272 23808 37281
rect 22836 37247 22888 37256
rect 22836 37213 22850 37247
rect 22850 37213 22884 37247
rect 22884 37213 22888 37247
rect 22836 37204 22888 37213
rect 23112 37204 23164 37256
rect 24768 37247 24820 37256
rect 16488 37111 16540 37120
rect 16488 37077 16497 37111
rect 16497 37077 16531 37111
rect 16531 37077 16540 37111
rect 16488 37068 16540 37077
rect 17500 37068 17552 37120
rect 17776 37111 17828 37120
rect 17776 37077 17785 37111
rect 17785 37077 17819 37111
rect 17819 37077 17828 37111
rect 17776 37068 17828 37077
rect 19432 37068 19484 37120
rect 20536 37068 20588 37120
rect 21548 37068 21600 37120
rect 22100 37068 22152 37120
rect 22468 37068 22520 37120
rect 23480 37136 23532 37188
rect 24768 37213 24777 37247
rect 24777 37213 24811 37247
rect 24811 37213 24820 37247
rect 24768 37204 24820 37213
rect 26240 37340 26292 37392
rect 25044 37247 25096 37256
rect 25044 37213 25053 37247
rect 25053 37213 25087 37247
rect 25087 37213 25096 37247
rect 25044 37204 25096 37213
rect 25964 37247 26016 37256
rect 24676 37136 24728 37188
rect 25964 37213 25973 37247
rect 25973 37213 26007 37247
rect 26007 37213 26016 37247
rect 25964 37204 26016 37213
rect 26240 37204 26292 37256
rect 26792 37204 26844 37256
rect 27804 37272 27856 37324
rect 28908 37340 28960 37392
rect 30288 37340 30340 37392
rect 30196 37272 30248 37324
rect 30932 37408 30984 37460
rect 32588 37408 32640 37460
rect 33876 37408 33928 37460
rect 34428 37408 34480 37460
rect 31668 37383 31720 37392
rect 31668 37349 31677 37383
rect 31677 37349 31711 37383
rect 31711 37349 31720 37383
rect 31668 37340 31720 37349
rect 33600 37340 33652 37392
rect 27712 37247 27764 37256
rect 27712 37213 27721 37247
rect 27721 37213 27755 37247
rect 27755 37213 27764 37247
rect 27712 37204 27764 37213
rect 28264 37204 28316 37256
rect 28448 37204 28500 37256
rect 26424 37136 26476 37188
rect 27252 37136 27304 37188
rect 22836 37068 22888 37120
rect 23664 37068 23716 37120
rect 24124 37068 24176 37120
rect 25872 37111 25924 37120
rect 25872 37077 25881 37111
rect 25881 37077 25915 37111
rect 25915 37077 25924 37111
rect 25872 37068 25924 37077
rect 26792 37068 26844 37120
rect 28816 37136 28868 37188
rect 30932 37204 30984 37256
rect 30104 37111 30156 37120
rect 30104 37077 30113 37111
rect 30113 37077 30147 37111
rect 30147 37077 30156 37111
rect 30104 37068 30156 37077
rect 30288 37068 30340 37120
rect 31024 37136 31076 37188
rect 31760 37247 31812 37256
rect 31760 37213 31769 37247
rect 31769 37213 31803 37247
rect 31803 37213 31812 37247
rect 31760 37204 31812 37213
rect 32588 37204 32640 37256
rect 33324 37272 33376 37324
rect 33140 37204 33192 37256
rect 33968 37204 34020 37256
rect 34060 37204 34112 37256
rect 33508 37136 33560 37188
rect 30932 37068 30984 37120
rect 31208 37068 31260 37120
rect 33600 37068 33652 37120
rect 34336 37136 34388 37188
rect 34980 37111 35032 37120
rect 34980 37077 34989 37111
rect 34989 37077 35023 37111
rect 35023 37077 35032 37111
rect 34980 37068 35032 37077
rect 36176 37111 36228 37120
rect 36176 37077 36185 37111
rect 36185 37077 36219 37111
rect 36219 37077 36228 37111
rect 36176 37068 36228 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 22468 36864 22520 36916
rect 22744 36864 22796 36916
rect 24124 36907 24176 36916
rect 24124 36873 24133 36907
rect 24133 36873 24167 36907
rect 24167 36873 24176 36907
rect 24124 36864 24176 36873
rect 25412 36864 25464 36916
rect 16304 36839 16356 36848
rect 16304 36805 16313 36839
rect 16313 36805 16347 36839
rect 16347 36805 16356 36839
rect 16304 36796 16356 36805
rect 22100 36839 22152 36848
rect 16120 36771 16172 36780
rect 16120 36737 16129 36771
rect 16129 36737 16163 36771
rect 16163 36737 16172 36771
rect 16120 36728 16172 36737
rect 17500 36771 17552 36780
rect 17500 36737 17509 36771
rect 17509 36737 17543 36771
rect 17543 36737 17552 36771
rect 17500 36728 17552 36737
rect 18788 36771 18840 36780
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 19616 36771 19668 36780
rect 19616 36737 19625 36771
rect 19625 36737 19659 36771
rect 19659 36737 19668 36771
rect 19616 36728 19668 36737
rect 20168 36728 20220 36780
rect 22100 36805 22109 36839
rect 22109 36805 22143 36839
rect 22143 36805 22152 36839
rect 22100 36796 22152 36805
rect 22192 36796 22244 36848
rect 15568 36660 15620 36712
rect 16856 36703 16908 36712
rect 16856 36669 16865 36703
rect 16865 36669 16899 36703
rect 16899 36669 16908 36703
rect 16856 36660 16908 36669
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 16120 36592 16172 36644
rect 17224 36592 17276 36644
rect 22468 36771 22520 36780
rect 22468 36737 22482 36771
rect 22482 36737 22516 36771
rect 22516 36737 22520 36771
rect 22468 36728 22520 36737
rect 23388 36728 23440 36780
rect 24400 36796 24452 36848
rect 24032 36728 24084 36780
rect 24216 36771 24268 36780
rect 24216 36737 24225 36771
rect 24225 36737 24259 36771
rect 24259 36737 24268 36771
rect 24216 36728 24268 36737
rect 25412 36728 25464 36780
rect 25872 36796 25924 36848
rect 29000 36864 29052 36916
rect 29920 36864 29972 36916
rect 31668 36907 31720 36916
rect 26608 36796 26660 36848
rect 26516 36728 26568 36780
rect 26976 36728 27028 36780
rect 28632 36796 28684 36848
rect 28724 36796 28776 36848
rect 22836 36660 22888 36712
rect 24768 36660 24820 36712
rect 28172 36728 28224 36780
rect 29000 36728 29052 36780
rect 29644 36728 29696 36780
rect 30012 36796 30064 36848
rect 20628 36592 20680 36644
rect 21824 36592 21876 36644
rect 28724 36660 28776 36712
rect 29736 36660 29788 36712
rect 30472 36728 30524 36780
rect 30748 36728 30800 36780
rect 31668 36873 31677 36907
rect 31677 36873 31711 36907
rect 31711 36873 31720 36907
rect 33876 36907 33928 36916
rect 31668 36864 31720 36873
rect 33876 36873 33885 36907
rect 33885 36873 33919 36907
rect 33919 36873 33928 36907
rect 33876 36864 33928 36873
rect 31116 36728 31168 36780
rect 31484 36771 31536 36780
rect 31484 36737 31493 36771
rect 31493 36737 31527 36771
rect 31527 36737 31536 36771
rect 31484 36728 31536 36737
rect 32496 36771 32548 36780
rect 32496 36737 32505 36771
rect 32505 36737 32539 36771
rect 32539 36737 32548 36771
rect 32496 36728 32548 36737
rect 32680 36771 32732 36780
rect 32680 36737 32689 36771
rect 32689 36737 32723 36771
rect 32723 36737 32732 36771
rect 32680 36728 32732 36737
rect 36176 36796 36228 36848
rect 33600 36728 33652 36780
rect 33784 36771 33836 36780
rect 33784 36737 33793 36771
rect 33793 36737 33827 36771
rect 33827 36737 33836 36771
rect 33784 36728 33836 36737
rect 33876 36728 33928 36780
rect 34980 36771 35032 36780
rect 34980 36737 34989 36771
rect 34989 36737 35023 36771
rect 35023 36737 35032 36771
rect 34980 36728 35032 36737
rect 30104 36703 30156 36712
rect 30104 36669 30113 36703
rect 30113 36669 30147 36703
rect 30147 36669 30156 36703
rect 31300 36703 31352 36712
rect 30104 36660 30156 36669
rect 31300 36669 31309 36703
rect 31309 36669 31343 36703
rect 31343 36669 31352 36703
rect 31300 36660 31352 36669
rect 34796 36660 34848 36712
rect 35440 36660 35492 36712
rect 36360 36703 36412 36712
rect 36360 36669 36369 36703
rect 36369 36669 36403 36703
rect 36403 36669 36412 36703
rect 36360 36660 36412 36669
rect 15568 36524 15620 36576
rect 20996 36524 21048 36576
rect 21548 36524 21600 36576
rect 25780 36524 25832 36576
rect 26148 36524 26200 36576
rect 26792 36524 26844 36576
rect 28080 36524 28132 36576
rect 28448 36567 28500 36576
rect 28448 36533 28457 36567
rect 28457 36533 28491 36567
rect 28491 36533 28500 36567
rect 28448 36524 28500 36533
rect 29644 36567 29696 36576
rect 29644 36533 29653 36567
rect 29653 36533 29687 36567
rect 29687 36533 29696 36567
rect 29644 36524 29696 36533
rect 30932 36524 30984 36576
rect 31116 36524 31168 36576
rect 31484 36524 31536 36576
rect 34060 36635 34112 36644
rect 34060 36601 34069 36635
rect 34069 36601 34103 36635
rect 34103 36601 34112 36635
rect 34060 36592 34112 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 17500 36363 17552 36372
rect 17500 36329 17509 36363
rect 17509 36329 17543 36363
rect 17543 36329 17552 36363
rect 17500 36320 17552 36329
rect 17592 36320 17644 36372
rect 19616 36320 19668 36372
rect 24768 36320 24820 36372
rect 25688 36320 25740 36372
rect 17224 36159 17276 36168
rect 17224 36125 17233 36159
rect 17233 36125 17267 36159
rect 17267 36125 17276 36159
rect 17224 36116 17276 36125
rect 19432 36252 19484 36304
rect 20352 36295 20404 36304
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 18788 36159 18840 36168
rect 18788 36125 18797 36159
rect 18797 36125 18831 36159
rect 18831 36125 18840 36159
rect 18788 36116 18840 36125
rect 19340 36116 19392 36168
rect 20352 36261 20361 36295
rect 20361 36261 20395 36295
rect 20395 36261 20404 36295
rect 20352 36252 20404 36261
rect 20720 36252 20772 36304
rect 20628 36227 20680 36236
rect 20628 36193 20637 36227
rect 20637 36193 20671 36227
rect 20671 36193 20680 36227
rect 20628 36184 20680 36193
rect 21548 36227 21600 36236
rect 21548 36193 21557 36227
rect 21557 36193 21591 36227
rect 21591 36193 21600 36227
rect 21548 36184 21600 36193
rect 20168 36116 20220 36168
rect 20536 36159 20588 36168
rect 20536 36125 20545 36159
rect 20545 36125 20579 36159
rect 20579 36125 20588 36159
rect 20536 36116 20588 36125
rect 21364 36159 21416 36168
rect 21364 36125 21373 36159
rect 21373 36125 21407 36159
rect 21407 36125 21416 36159
rect 21364 36116 21416 36125
rect 23204 36252 23256 36304
rect 22376 36184 22428 36236
rect 22928 36184 22980 36236
rect 24584 36184 24636 36236
rect 24492 36116 24544 36168
rect 26516 36252 26568 36304
rect 27068 36295 27120 36304
rect 27068 36261 27077 36295
rect 27077 36261 27111 36295
rect 27111 36261 27120 36295
rect 27068 36252 27120 36261
rect 28908 36320 28960 36372
rect 29000 36320 29052 36372
rect 30104 36320 30156 36372
rect 30840 36320 30892 36372
rect 31300 36320 31352 36372
rect 33140 36320 33192 36372
rect 28632 36252 28684 36304
rect 33416 36252 33468 36304
rect 33876 36252 33928 36304
rect 21916 36048 21968 36100
rect 23848 36091 23900 36100
rect 23848 36057 23857 36091
rect 23857 36057 23891 36091
rect 23891 36057 23900 36091
rect 23848 36048 23900 36057
rect 24216 36048 24268 36100
rect 25044 36159 25096 36168
rect 25044 36125 25053 36159
rect 25053 36125 25087 36159
rect 25087 36125 25096 36159
rect 25044 36116 25096 36125
rect 26424 36116 26476 36168
rect 26792 36159 26844 36168
rect 26792 36125 26801 36159
rect 26801 36125 26835 36159
rect 26835 36125 26844 36159
rect 26792 36116 26844 36125
rect 26884 36159 26936 36168
rect 26884 36125 26893 36159
rect 26893 36125 26927 36159
rect 26927 36125 26936 36159
rect 27620 36184 27672 36236
rect 26884 36116 26936 36125
rect 30656 36184 30708 36236
rect 25596 36048 25648 36100
rect 26976 36048 27028 36100
rect 19432 35980 19484 36032
rect 20720 36023 20772 36032
rect 20720 35989 20729 36023
rect 20729 35989 20763 36023
rect 20763 35989 20772 36023
rect 20720 35980 20772 35989
rect 22100 35980 22152 36032
rect 24768 35980 24820 36032
rect 24860 35980 24912 36032
rect 28264 36116 28316 36168
rect 28724 36091 28776 36100
rect 28724 36057 28733 36091
rect 28733 36057 28767 36091
rect 28767 36057 28776 36091
rect 28724 36048 28776 36057
rect 29184 36116 29236 36168
rect 30380 36116 30432 36168
rect 30564 36116 30616 36168
rect 32680 36227 32732 36236
rect 32680 36193 32689 36227
rect 32689 36193 32723 36227
rect 32723 36193 32732 36227
rect 32680 36184 32732 36193
rect 34704 36184 34756 36236
rect 31024 36159 31076 36168
rect 31024 36125 31033 36159
rect 31033 36125 31067 36159
rect 31067 36125 31076 36159
rect 31024 36116 31076 36125
rect 31484 36116 31536 36168
rect 32772 36159 32824 36168
rect 32772 36125 32781 36159
rect 32781 36125 32815 36159
rect 32815 36125 32824 36159
rect 32772 36116 32824 36125
rect 33140 36116 33192 36168
rect 33508 36116 33560 36168
rect 34336 36159 34388 36168
rect 34336 36125 34345 36159
rect 34345 36125 34379 36159
rect 34379 36125 34388 36159
rect 34336 36116 34388 36125
rect 34888 36159 34940 36168
rect 34888 36125 34897 36159
rect 34897 36125 34931 36159
rect 34931 36125 34940 36159
rect 34888 36116 34940 36125
rect 32128 36048 32180 36100
rect 35256 36159 35308 36168
rect 35256 36125 35265 36159
rect 35265 36125 35299 36159
rect 35299 36125 35308 36159
rect 35256 36116 35308 36125
rect 27896 35980 27948 36032
rect 30288 36023 30340 36032
rect 30288 35989 30297 36023
rect 30297 35989 30331 36023
rect 30331 35989 30340 36023
rect 30288 35980 30340 35989
rect 31944 35980 31996 36032
rect 33968 35980 34020 36032
rect 35164 35980 35216 36032
rect 36176 35980 36228 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 14280 35776 14332 35828
rect 15568 35776 15620 35828
rect 16120 35776 16172 35828
rect 23756 35776 23808 35828
rect 24492 35776 24544 35828
rect 28080 35819 28132 35828
rect 15200 35708 15252 35760
rect 15384 35708 15436 35760
rect 21456 35751 21508 35760
rect 14096 35683 14148 35692
rect 14096 35649 14105 35683
rect 14105 35649 14139 35683
rect 14139 35649 14148 35683
rect 14096 35640 14148 35649
rect 14924 35683 14976 35692
rect 14924 35649 14933 35683
rect 14933 35649 14967 35683
rect 14967 35649 14976 35683
rect 14924 35640 14976 35649
rect 15016 35683 15068 35692
rect 15016 35649 15025 35683
rect 15025 35649 15059 35683
rect 15059 35649 15068 35683
rect 15016 35640 15068 35649
rect 15752 35683 15804 35692
rect 15752 35649 15761 35683
rect 15761 35649 15795 35683
rect 15795 35649 15804 35683
rect 15752 35640 15804 35649
rect 21456 35717 21465 35751
rect 21465 35717 21499 35751
rect 21499 35717 21508 35751
rect 21456 35708 21508 35717
rect 22836 35751 22888 35760
rect 22836 35717 22845 35751
rect 22845 35717 22879 35751
rect 22879 35717 22888 35751
rect 22836 35708 22888 35717
rect 23112 35708 23164 35760
rect 24216 35751 24268 35760
rect 24216 35717 24225 35751
rect 24225 35717 24259 35751
rect 24259 35717 24268 35751
rect 24216 35708 24268 35717
rect 28080 35785 28089 35819
rect 28089 35785 28123 35819
rect 28123 35785 28132 35819
rect 28080 35776 28132 35785
rect 29000 35776 29052 35828
rect 15936 35683 15988 35692
rect 15936 35649 15945 35683
rect 15945 35649 15979 35683
rect 15979 35649 15988 35683
rect 15936 35640 15988 35649
rect 17040 35640 17092 35692
rect 17132 35615 17184 35624
rect 17132 35581 17141 35615
rect 17141 35581 17175 35615
rect 17175 35581 17184 35615
rect 17132 35572 17184 35581
rect 19524 35640 19576 35692
rect 19708 35640 19760 35692
rect 20076 35640 20128 35692
rect 20352 35640 20404 35692
rect 20536 35640 20588 35692
rect 22284 35640 22336 35692
rect 22744 35683 22796 35692
rect 22744 35649 22751 35683
rect 22751 35649 22796 35683
rect 20168 35615 20220 35624
rect 20168 35581 20177 35615
rect 20177 35581 20211 35615
rect 20211 35581 20220 35615
rect 20168 35572 20220 35581
rect 20904 35572 20956 35624
rect 22744 35640 22796 35649
rect 23020 35683 23072 35692
rect 23020 35649 23034 35683
rect 23034 35649 23068 35683
rect 23068 35649 23072 35683
rect 23020 35640 23072 35649
rect 23848 35640 23900 35692
rect 26148 35708 26200 35760
rect 27068 35708 27120 35760
rect 27344 35751 27396 35760
rect 27344 35717 27353 35751
rect 27353 35717 27387 35751
rect 27387 35717 27396 35751
rect 27344 35708 27396 35717
rect 23940 35572 23992 35624
rect 25688 35640 25740 35692
rect 25872 35640 25924 35692
rect 26884 35640 26936 35692
rect 25412 35572 25464 35624
rect 26332 35572 26384 35624
rect 28448 35640 28500 35692
rect 28908 35640 28960 35692
rect 29184 35683 29236 35692
rect 29184 35649 29193 35683
rect 29193 35649 29227 35683
rect 29227 35649 29236 35683
rect 29184 35640 29236 35649
rect 29092 35572 29144 35624
rect 18512 35436 18564 35488
rect 20076 35504 20128 35556
rect 25596 35504 25648 35556
rect 26608 35504 26660 35556
rect 29828 35708 29880 35760
rect 31392 35776 31444 35828
rect 32680 35819 32732 35828
rect 32680 35785 32689 35819
rect 32689 35785 32723 35819
rect 32723 35785 32732 35819
rect 32680 35776 32732 35785
rect 33508 35776 33560 35828
rect 34888 35776 34940 35828
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 29920 35640 29972 35649
rect 30288 35640 30340 35692
rect 29552 35615 29604 35624
rect 29552 35581 29561 35615
rect 29561 35581 29595 35615
rect 29595 35581 29604 35615
rect 31116 35683 31168 35692
rect 31116 35649 31125 35683
rect 31125 35649 31159 35683
rect 31159 35649 31168 35683
rect 31116 35640 31168 35649
rect 32404 35708 32456 35760
rect 29552 35572 29604 35581
rect 19432 35479 19484 35488
rect 19432 35445 19441 35479
rect 19441 35445 19475 35479
rect 19475 35445 19484 35479
rect 19432 35436 19484 35445
rect 23204 35479 23256 35488
rect 23204 35445 23213 35479
rect 23213 35445 23247 35479
rect 23247 35445 23256 35479
rect 23204 35436 23256 35445
rect 26148 35436 26200 35488
rect 27160 35436 27212 35488
rect 29092 35436 29144 35488
rect 30840 35436 30892 35488
rect 32956 35572 33008 35624
rect 34244 35708 34296 35760
rect 36176 35708 36228 35760
rect 34796 35683 34848 35692
rect 34796 35649 34805 35683
rect 34805 35649 34839 35683
rect 34839 35649 34848 35683
rect 34796 35640 34848 35649
rect 35164 35683 35216 35692
rect 35164 35649 35173 35683
rect 35173 35649 35207 35683
rect 35207 35649 35216 35683
rect 35164 35640 35216 35649
rect 35256 35640 35308 35692
rect 34520 35572 34572 35624
rect 35992 35572 36044 35624
rect 32496 35479 32548 35488
rect 32496 35445 32505 35479
rect 32505 35445 32539 35479
rect 32539 35445 32548 35479
rect 32496 35436 32548 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 14096 35232 14148 35284
rect 15016 35232 15068 35284
rect 19524 35275 19576 35284
rect 19524 35241 19533 35275
rect 19533 35241 19567 35275
rect 19567 35241 19576 35275
rect 19524 35232 19576 35241
rect 22744 35232 22796 35284
rect 15752 35096 15804 35148
rect 15568 35071 15620 35080
rect 15568 35037 15577 35071
rect 15577 35037 15611 35071
rect 15611 35037 15620 35071
rect 15568 35028 15620 35037
rect 17040 35071 17092 35080
rect 17040 35037 17049 35071
rect 17049 35037 17083 35071
rect 17083 35037 17092 35071
rect 17040 35028 17092 35037
rect 17132 35028 17184 35080
rect 19432 35164 19484 35216
rect 18236 35096 18288 35148
rect 19708 35096 19760 35148
rect 20352 35096 20404 35148
rect 19340 35028 19392 35080
rect 20536 35071 20588 35080
rect 20536 35037 20545 35071
rect 20545 35037 20579 35071
rect 20579 35037 20588 35071
rect 20536 35028 20588 35037
rect 14924 35003 14976 35012
rect 14924 34969 14933 35003
rect 14933 34969 14967 35003
rect 14967 34969 14976 35003
rect 14924 34960 14976 34969
rect 20904 35071 20956 35080
rect 20904 35037 20913 35071
rect 20913 35037 20947 35071
rect 20947 35037 20956 35071
rect 22928 35096 22980 35148
rect 25872 35232 25924 35284
rect 30840 35275 30892 35284
rect 30840 35241 30849 35275
rect 30849 35241 30883 35275
rect 30883 35241 30892 35275
rect 30840 35232 30892 35241
rect 29368 35164 29420 35216
rect 20904 35028 20956 35037
rect 22836 35071 22888 35080
rect 22836 35037 22845 35071
rect 22845 35037 22879 35071
rect 22879 35037 22888 35071
rect 22836 35028 22888 35037
rect 24952 35096 25004 35148
rect 24768 35071 24820 35080
rect 24768 35037 24777 35071
rect 24777 35037 24811 35071
rect 24811 35037 24820 35071
rect 24768 35028 24820 35037
rect 25044 35071 25096 35080
rect 25044 35037 25053 35071
rect 25053 35037 25087 35071
rect 25087 35037 25096 35071
rect 25044 35028 25096 35037
rect 28816 35096 28868 35148
rect 29460 35096 29512 35148
rect 29828 35139 29880 35148
rect 29828 35105 29837 35139
rect 29837 35105 29871 35139
rect 29871 35105 29880 35139
rect 29828 35096 29880 35105
rect 30104 35139 30156 35148
rect 30104 35105 30113 35139
rect 30113 35105 30147 35139
rect 30147 35105 30156 35139
rect 30104 35096 30156 35105
rect 31024 35096 31076 35148
rect 31484 35096 31536 35148
rect 26608 35071 26660 35080
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26608 35028 26660 35037
rect 27068 35071 27120 35080
rect 27068 35037 27077 35071
rect 27077 35037 27111 35071
rect 27111 35037 27120 35071
rect 27068 35028 27120 35037
rect 1676 34935 1728 34944
rect 1676 34901 1685 34935
rect 1685 34901 1719 34935
rect 1719 34901 1728 34935
rect 1676 34892 1728 34901
rect 2044 34892 2096 34944
rect 15200 34892 15252 34944
rect 15660 34892 15712 34944
rect 15936 34892 15988 34944
rect 21088 34892 21140 34944
rect 21640 34935 21692 34944
rect 21640 34901 21649 34935
rect 21649 34901 21683 34935
rect 21683 34901 21692 34935
rect 21640 34892 21692 34901
rect 21732 34892 21784 34944
rect 23388 34960 23440 35012
rect 25688 34960 25740 35012
rect 26332 35003 26384 35012
rect 26332 34969 26341 35003
rect 26341 34969 26375 35003
rect 26375 34969 26384 35003
rect 26332 34960 26384 34969
rect 26516 34960 26568 35012
rect 27804 34960 27856 35012
rect 23664 34892 23716 34944
rect 24584 34935 24636 34944
rect 24584 34901 24593 34935
rect 24593 34901 24627 34935
rect 24627 34901 24636 34935
rect 24584 34892 24636 34901
rect 26056 34935 26108 34944
rect 26056 34901 26065 34935
rect 26065 34901 26099 34935
rect 26099 34901 26108 34935
rect 26056 34892 26108 34901
rect 27252 34935 27304 34944
rect 27252 34901 27261 34935
rect 27261 34901 27295 34935
rect 27295 34901 27304 34935
rect 27252 34892 27304 34901
rect 28540 35071 28592 35080
rect 28540 35037 28549 35071
rect 28549 35037 28583 35071
rect 28583 35037 28592 35071
rect 28540 35028 28592 35037
rect 28908 35028 28960 35080
rect 29736 35028 29788 35080
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30840 35028 30892 35080
rect 31852 35139 31904 35148
rect 31852 35105 31861 35139
rect 31861 35105 31895 35139
rect 31895 35105 31904 35139
rect 33048 35164 33100 35216
rect 31852 35096 31904 35105
rect 33508 35096 33560 35148
rect 28724 34960 28776 35012
rect 29184 34960 29236 35012
rect 29000 34892 29052 34944
rect 30564 34960 30616 35012
rect 30932 34960 30984 35012
rect 31944 35071 31996 35080
rect 31944 35037 31953 35071
rect 31953 35037 31987 35071
rect 31987 35037 31996 35071
rect 31944 35028 31996 35037
rect 32128 35071 32180 35080
rect 32128 35037 32137 35071
rect 32137 35037 32171 35071
rect 32171 35037 32180 35071
rect 32128 35028 32180 35037
rect 32496 35028 32548 35080
rect 33048 35028 33100 35080
rect 33324 35071 33376 35080
rect 33324 35037 33333 35071
rect 33333 35037 33367 35071
rect 33367 35037 33376 35071
rect 33324 35028 33376 35037
rect 31852 34960 31904 35012
rect 33600 35028 33652 35080
rect 34796 35096 34848 35148
rect 34060 35028 34112 35080
rect 31116 34892 31168 34944
rect 31576 34892 31628 34944
rect 32680 34892 32732 34944
rect 33140 34892 33192 34944
rect 33324 34892 33376 34944
rect 33416 34892 33468 34944
rect 36912 34892 36964 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 14924 34688 14976 34740
rect 18236 34731 18288 34740
rect 18236 34697 18245 34731
rect 18245 34697 18279 34731
rect 18279 34697 18288 34731
rect 18236 34688 18288 34697
rect 20904 34688 20956 34740
rect 15200 34620 15252 34672
rect 18512 34620 18564 34672
rect 18788 34620 18840 34672
rect 20076 34620 20128 34672
rect 22376 34620 22428 34672
rect 22560 34688 22612 34740
rect 23020 34688 23072 34740
rect 23204 34620 23256 34672
rect 15108 34527 15160 34536
rect 15108 34493 15117 34527
rect 15117 34493 15151 34527
rect 15151 34493 15160 34527
rect 21732 34552 21784 34604
rect 23480 34552 23532 34604
rect 23664 34595 23716 34604
rect 23664 34561 23673 34595
rect 23673 34561 23707 34595
rect 23707 34561 23716 34595
rect 24952 34688 25004 34740
rect 25044 34688 25096 34740
rect 25228 34620 25280 34672
rect 26056 34620 26108 34672
rect 26792 34620 26844 34672
rect 27620 34620 27672 34672
rect 27896 34663 27948 34672
rect 27896 34629 27905 34663
rect 27905 34629 27939 34663
rect 27939 34629 27948 34663
rect 27896 34620 27948 34629
rect 29000 34688 29052 34740
rect 29828 34620 29880 34672
rect 23664 34552 23716 34561
rect 25596 34595 25648 34604
rect 15108 34484 15160 34493
rect 19248 34484 19300 34536
rect 21088 34527 21140 34536
rect 21088 34493 21097 34527
rect 21097 34493 21131 34527
rect 21131 34493 21140 34527
rect 21088 34484 21140 34493
rect 22008 34484 22060 34536
rect 22652 34484 22704 34536
rect 25596 34561 25605 34595
rect 25605 34561 25639 34595
rect 25639 34561 25648 34595
rect 25596 34552 25648 34561
rect 27252 34552 27304 34604
rect 25504 34484 25556 34536
rect 26424 34484 26476 34536
rect 27804 34552 27856 34604
rect 28080 34595 28132 34604
rect 28080 34561 28089 34595
rect 28089 34561 28123 34595
rect 28123 34561 28132 34595
rect 28816 34595 28868 34604
rect 28080 34552 28132 34561
rect 28816 34561 28825 34595
rect 28825 34561 28859 34595
rect 28859 34561 28868 34595
rect 28816 34552 28868 34561
rect 29276 34552 29328 34604
rect 29736 34595 29788 34604
rect 29736 34561 29745 34595
rect 29745 34561 29779 34595
rect 29779 34561 29788 34595
rect 29736 34552 29788 34561
rect 30196 34552 30248 34604
rect 31116 34595 31168 34604
rect 31116 34561 31125 34595
rect 31125 34561 31159 34595
rect 31159 34561 31168 34595
rect 31116 34552 31168 34561
rect 29920 34484 29972 34536
rect 30656 34527 30708 34536
rect 30656 34493 30665 34527
rect 30665 34493 30699 34527
rect 30699 34493 30708 34527
rect 30656 34484 30708 34493
rect 30932 34527 30984 34536
rect 30932 34493 30941 34527
rect 30941 34493 30975 34527
rect 30975 34493 30984 34527
rect 30932 34484 30984 34493
rect 31024 34527 31076 34536
rect 31024 34493 31033 34527
rect 31033 34493 31067 34527
rect 31067 34493 31076 34527
rect 57888 34688 57940 34740
rect 33140 34620 33192 34672
rect 34060 34620 34112 34672
rect 33324 34552 33376 34604
rect 33692 34552 33744 34604
rect 33876 34595 33928 34604
rect 33876 34561 33885 34595
rect 33885 34561 33919 34595
rect 33919 34561 33928 34595
rect 33876 34552 33928 34561
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 35532 34552 35584 34561
rect 35716 34595 35768 34604
rect 35716 34561 35725 34595
rect 35725 34561 35759 34595
rect 35759 34561 35768 34595
rect 35716 34552 35768 34561
rect 31024 34484 31076 34493
rect 31392 34484 31444 34536
rect 31944 34484 31996 34536
rect 33968 34527 34020 34536
rect 33968 34493 33977 34527
rect 33977 34493 34011 34527
rect 34011 34493 34020 34527
rect 33968 34484 34020 34493
rect 37464 34552 37516 34604
rect 36728 34484 36780 34536
rect 57428 34527 57480 34536
rect 57428 34493 57437 34527
rect 57437 34493 57471 34527
rect 57471 34493 57480 34527
rect 57428 34484 57480 34493
rect 21732 34416 21784 34468
rect 22744 34416 22796 34468
rect 26792 34416 26844 34468
rect 33048 34416 33100 34468
rect 38936 34416 38988 34468
rect 15384 34348 15436 34400
rect 20352 34391 20404 34400
rect 20352 34357 20361 34391
rect 20361 34357 20395 34391
rect 20395 34357 20404 34391
rect 20352 34348 20404 34357
rect 21088 34348 21140 34400
rect 27988 34348 28040 34400
rect 28264 34391 28316 34400
rect 28264 34357 28273 34391
rect 28273 34357 28307 34391
rect 28307 34357 28316 34391
rect 28264 34348 28316 34357
rect 29000 34348 29052 34400
rect 35624 34391 35676 34400
rect 35624 34357 35633 34391
rect 35633 34357 35667 34391
rect 35667 34357 35676 34391
rect 35624 34348 35676 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 15660 34187 15712 34196
rect 15660 34153 15669 34187
rect 15669 34153 15703 34187
rect 15703 34153 15712 34187
rect 15660 34144 15712 34153
rect 20352 34144 20404 34196
rect 21456 34144 21508 34196
rect 23572 34187 23624 34196
rect 23572 34153 23581 34187
rect 23581 34153 23615 34187
rect 23615 34153 23624 34187
rect 23572 34144 23624 34153
rect 17408 34119 17460 34128
rect 17408 34085 17417 34119
rect 17417 34085 17451 34119
rect 17451 34085 17460 34119
rect 17408 34076 17460 34085
rect 16212 34008 16264 34060
rect 15292 33983 15344 33992
rect 15292 33949 15301 33983
rect 15301 33949 15335 33983
rect 15335 33949 15344 33983
rect 15292 33940 15344 33949
rect 18512 34076 18564 34128
rect 19432 34008 19484 34060
rect 23480 34076 23532 34128
rect 20536 34008 20588 34060
rect 24952 34008 25004 34060
rect 25228 34051 25280 34060
rect 25228 34017 25237 34051
rect 25237 34017 25271 34051
rect 25271 34017 25280 34051
rect 25228 34008 25280 34017
rect 27160 34008 27212 34060
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 27712 34051 27764 34060
rect 27712 34017 27721 34051
rect 27721 34017 27755 34051
rect 27755 34017 27764 34051
rect 27712 34008 27764 34017
rect 29000 34008 29052 34060
rect 31024 34076 31076 34128
rect 31116 34076 31168 34128
rect 32128 34076 32180 34128
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 18512 33983 18564 33992
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 18604 33983 18656 33992
rect 18604 33949 18613 33983
rect 18613 33949 18647 33983
rect 18647 33949 18656 33983
rect 19984 33983 20036 33992
rect 18604 33940 18656 33949
rect 19984 33949 19993 33983
rect 19993 33949 20027 33983
rect 20027 33949 20036 33983
rect 19984 33940 20036 33949
rect 21640 33940 21692 33992
rect 22744 33983 22796 33992
rect 22744 33949 22753 33983
rect 22753 33949 22787 33983
rect 22787 33949 22796 33983
rect 22744 33940 22796 33949
rect 23020 33940 23072 33992
rect 25964 33940 26016 33992
rect 26608 33940 26660 33992
rect 26976 33940 27028 33992
rect 29092 33940 29144 33992
rect 29828 34008 29880 34060
rect 30932 34008 30984 34060
rect 31116 33940 31168 33992
rect 17960 33804 18012 33856
rect 18328 33804 18380 33856
rect 20260 33804 20312 33856
rect 21272 33847 21324 33856
rect 21272 33813 21281 33847
rect 21281 33813 21315 33847
rect 21315 33813 21324 33847
rect 21272 33804 21324 33813
rect 21456 33872 21508 33924
rect 22100 33915 22152 33924
rect 22100 33881 22109 33915
rect 22109 33881 22143 33915
rect 22143 33881 22152 33915
rect 23756 33915 23808 33924
rect 22100 33872 22152 33881
rect 23756 33881 23765 33915
rect 23765 33881 23799 33915
rect 23799 33881 23808 33915
rect 23756 33872 23808 33881
rect 24768 33872 24820 33924
rect 25688 33872 25740 33924
rect 22192 33804 22244 33856
rect 24032 33804 24084 33856
rect 24676 33804 24728 33856
rect 24952 33847 25004 33856
rect 24952 33813 24961 33847
rect 24961 33813 24995 33847
rect 24995 33813 25004 33847
rect 24952 33804 25004 33813
rect 25044 33804 25096 33856
rect 25780 33804 25832 33856
rect 27436 33804 27488 33856
rect 28448 33804 28500 33856
rect 28724 33847 28776 33856
rect 28724 33813 28733 33847
rect 28733 33813 28767 33847
rect 28767 33813 28776 33847
rect 28724 33804 28776 33813
rect 30564 33804 30616 33856
rect 31760 34008 31812 34060
rect 33416 34119 33468 34128
rect 33416 34085 33425 34119
rect 33425 34085 33459 34119
rect 33459 34085 33468 34119
rect 33416 34076 33468 34085
rect 35532 34144 35584 34196
rect 34980 34051 35032 34060
rect 34980 34017 34989 34051
rect 34989 34017 35023 34051
rect 35023 34017 35032 34051
rect 34980 34008 35032 34017
rect 31484 33983 31536 33992
rect 31484 33949 31493 33983
rect 31493 33949 31527 33983
rect 31527 33949 31536 33983
rect 32680 33983 32732 33992
rect 31484 33940 31536 33949
rect 32680 33949 32689 33983
rect 32689 33949 32723 33983
rect 32723 33949 32732 33983
rect 32680 33940 32732 33949
rect 33140 33983 33192 33992
rect 33140 33949 33149 33983
rect 33149 33949 33183 33983
rect 33183 33949 33192 33983
rect 33140 33940 33192 33949
rect 31392 33872 31444 33924
rect 31300 33804 31352 33856
rect 31852 33804 31904 33856
rect 32772 33804 32824 33856
rect 34428 33940 34480 33992
rect 35716 33940 35768 33992
rect 40224 34076 40276 34128
rect 36636 33940 36688 33992
rect 38936 33983 38988 33992
rect 38936 33949 38945 33983
rect 38945 33949 38979 33983
rect 38979 33949 38988 33983
rect 38936 33940 38988 33949
rect 38844 33872 38896 33924
rect 35808 33804 35860 33856
rect 38752 33847 38804 33856
rect 38752 33813 38761 33847
rect 38761 33813 38795 33847
rect 38795 33813 38804 33847
rect 38752 33804 38804 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 19432 33600 19484 33652
rect 21088 33600 21140 33652
rect 22192 33643 22244 33652
rect 22192 33609 22201 33643
rect 22201 33609 22235 33643
rect 22235 33609 22244 33643
rect 22192 33600 22244 33609
rect 23020 33643 23072 33652
rect 23020 33609 23029 33643
rect 23029 33609 23063 33643
rect 23063 33609 23072 33643
rect 23020 33600 23072 33609
rect 15200 33396 15252 33448
rect 15292 33396 15344 33448
rect 16212 33464 16264 33516
rect 23204 33532 23256 33584
rect 24032 33575 24084 33584
rect 17960 33507 18012 33516
rect 17960 33473 17969 33507
rect 17969 33473 18003 33507
rect 18003 33473 18012 33507
rect 17960 33464 18012 33473
rect 18512 33464 18564 33516
rect 20260 33464 20312 33516
rect 20720 33464 20772 33516
rect 20996 33507 21048 33516
rect 20996 33473 21005 33507
rect 21005 33473 21039 33507
rect 21039 33473 21048 33507
rect 20996 33464 21048 33473
rect 22376 33464 22428 33516
rect 23112 33464 23164 33516
rect 24032 33541 24041 33575
rect 24041 33541 24075 33575
rect 24075 33541 24084 33575
rect 24032 33532 24084 33541
rect 24584 33532 24636 33584
rect 24768 33575 24820 33584
rect 24768 33541 24777 33575
rect 24777 33541 24811 33575
rect 24811 33541 24820 33575
rect 24768 33532 24820 33541
rect 25596 33600 25648 33652
rect 26608 33600 26660 33652
rect 27252 33643 27304 33652
rect 27252 33609 27261 33643
rect 27261 33609 27295 33643
rect 27295 33609 27304 33643
rect 27252 33600 27304 33609
rect 28172 33643 28224 33652
rect 28172 33609 28181 33643
rect 28181 33609 28215 33643
rect 28215 33609 28224 33643
rect 28172 33600 28224 33609
rect 28724 33600 28776 33652
rect 31760 33600 31812 33652
rect 33876 33600 33928 33652
rect 34980 33600 35032 33652
rect 37464 33600 37516 33652
rect 38752 33600 38804 33652
rect 23572 33464 23624 33516
rect 23848 33507 23900 33516
rect 23848 33473 23857 33507
rect 23857 33473 23891 33507
rect 23891 33473 23900 33507
rect 25044 33532 25096 33584
rect 26424 33575 26476 33584
rect 26424 33541 26433 33575
rect 26433 33541 26467 33575
rect 26467 33541 26476 33575
rect 26424 33532 26476 33541
rect 25596 33507 25648 33516
rect 23848 33464 23900 33473
rect 25596 33473 25605 33507
rect 25605 33473 25639 33507
rect 25639 33473 25648 33507
rect 25596 33464 25648 33473
rect 27160 33507 27212 33516
rect 15660 33328 15712 33380
rect 22928 33439 22980 33448
rect 22928 33405 22937 33439
rect 22937 33405 22971 33439
rect 22971 33405 22980 33439
rect 22928 33396 22980 33405
rect 23664 33396 23716 33448
rect 24952 33396 25004 33448
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 30472 33532 30524 33584
rect 30288 33507 30340 33516
rect 30288 33473 30297 33507
rect 30297 33473 30331 33507
rect 30331 33473 30340 33507
rect 30288 33464 30340 33473
rect 31300 33532 31352 33584
rect 31208 33507 31260 33516
rect 31208 33473 31217 33507
rect 31217 33473 31251 33507
rect 31251 33473 31260 33507
rect 31208 33464 31260 33473
rect 31392 33464 31444 33516
rect 33140 33532 33192 33584
rect 33600 33575 33652 33584
rect 33600 33541 33609 33575
rect 33609 33541 33643 33575
rect 33643 33541 33652 33575
rect 33600 33532 33652 33541
rect 34152 33532 34204 33584
rect 32496 33507 32548 33516
rect 32496 33473 32505 33507
rect 32505 33473 32539 33507
rect 32539 33473 32548 33507
rect 32496 33464 32548 33473
rect 21640 33328 21692 33380
rect 15936 33260 15988 33312
rect 18420 33260 18472 33312
rect 20444 33260 20496 33312
rect 23572 33260 23624 33312
rect 26700 33328 26752 33380
rect 32220 33396 32272 33448
rect 32772 33464 32824 33516
rect 35624 33507 35676 33516
rect 35624 33473 35633 33507
rect 35633 33473 35667 33507
rect 35667 33473 35676 33507
rect 35624 33464 35676 33473
rect 35808 33507 35860 33516
rect 35808 33473 35817 33507
rect 35817 33473 35851 33507
rect 35851 33473 35860 33507
rect 35808 33464 35860 33473
rect 36636 33507 36688 33516
rect 36636 33473 36645 33507
rect 36645 33473 36679 33507
rect 36679 33473 36688 33507
rect 36636 33464 36688 33473
rect 37464 33507 37516 33516
rect 37464 33473 37473 33507
rect 37473 33473 37507 33507
rect 37507 33473 37516 33507
rect 37464 33464 37516 33473
rect 38844 33532 38896 33584
rect 29184 33371 29236 33380
rect 29184 33337 29193 33371
rect 29193 33337 29227 33371
rect 29227 33337 29236 33371
rect 35532 33396 35584 33448
rect 36728 33439 36780 33448
rect 36728 33405 36737 33439
rect 36737 33405 36771 33439
rect 36771 33405 36780 33439
rect 36728 33396 36780 33405
rect 29184 33328 29236 33337
rect 34428 33328 34480 33380
rect 38936 33464 38988 33516
rect 39672 33507 39724 33516
rect 39672 33473 39681 33507
rect 39681 33473 39715 33507
rect 39715 33473 39724 33507
rect 39672 33464 39724 33473
rect 40040 33507 40092 33516
rect 40040 33473 40049 33507
rect 40049 33473 40083 33507
rect 40083 33473 40092 33507
rect 40040 33464 40092 33473
rect 52276 33396 52328 33448
rect 26332 33260 26384 33312
rect 30840 33260 30892 33312
rect 32956 33303 33008 33312
rect 32956 33269 32965 33303
rect 32965 33269 32999 33303
rect 32999 33269 33008 33303
rect 32956 33260 33008 33269
rect 35716 33303 35768 33312
rect 35716 33269 35725 33303
rect 35725 33269 35759 33303
rect 35759 33269 35768 33303
rect 35716 33260 35768 33269
rect 36820 33260 36872 33312
rect 38752 33303 38804 33312
rect 38752 33269 38761 33303
rect 38761 33269 38795 33303
rect 38795 33269 38804 33303
rect 38752 33260 38804 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 21272 33056 21324 33108
rect 22836 33056 22888 33108
rect 26608 33056 26660 33108
rect 26792 33056 26844 33108
rect 31300 33099 31352 33108
rect 31300 33065 31309 33099
rect 31309 33065 31343 33099
rect 31343 33065 31352 33099
rect 31300 33056 31352 33065
rect 31944 33099 31996 33108
rect 31944 33065 31953 33099
rect 31953 33065 31987 33099
rect 31987 33065 31996 33099
rect 31944 33056 31996 33065
rect 32496 33056 32548 33108
rect 33232 33099 33284 33108
rect 33232 33065 33241 33099
rect 33241 33065 33275 33099
rect 33275 33065 33284 33099
rect 33232 33056 33284 33065
rect 34060 33099 34112 33108
rect 34060 33065 34069 33099
rect 34069 33065 34103 33099
rect 34103 33065 34112 33099
rect 34060 33056 34112 33065
rect 38844 33099 38896 33108
rect 38844 33065 38853 33099
rect 38853 33065 38887 33099
rect 38887 33065 38896 33099
rect 38844 33056 38896 33065
rect 40040 33056 40092 33108
rect 15200 32988 15252 33040
rect 20444 32988 20496 33040
rect 15660 32963 15712 32972
rect 15660 32929 15669 32963
rect 15669 32929 15703 32963
rect 15703 32929 15712 32963
rect 15660 32920 15712 32929
rect 18328 32920 18380 32972
rect 17408 32852 17460 32904
rect 17776 32852 17828 32904
rect 21272 32895 21324 32904
rect 19248 32784 19300 32836
rect 16120 32759 16172 32768
rect 16120 32725 16129 32759
rect 16129 32725 16163 32759
rect 16163 32725 16172 32759
rect 16120 32716 16172 32725
rect 18604 32716 18656 32768
rect 20628 32716 20680 32768
rect 21272 32861 21281 32895
rect 21281 32861 21315 32895
rect 21315 32861 21324 32895
rect 21272 32852 21324 32861
rect 22100 32920 22152 32972
rect 22836 32852 22888 32904
rect 23388 32988 23440 33040
rect 26056 32988 26108 33040
rect 26516 32988 26568 33040
rect 25688 32920 25740 32972
rect 25872 32920 25924 32972
rect 26700 32920 26752 32972
rect 23296 32895 23348 32904
rect 23296 32861 23305 32895
rect 23305 32861 23339 32895
rect 23339 32861 23348 32895
rect 23296 32852 23348 32861
rect 24676 32852 24728 32904
rect 24860 32895 24912 32904
rect 24860 32861 24869 32895
rect 24869 32861 24903 32895
rect 24903 32861 24912 32895
rect 24860 32852 24912 32861
rect 26332 32895 26384 32904
rect 26332 32861 26340 32895
rect 26340 32861 26374 32895
rect 26374 32861 26384 32895
rect 26332 32852 26384 32861
rect 27160 32852 27212 32904
rect 34428 32988 34480 33040
rect 28264 32920 28316 32972
rect 28816 32852 28868 32904
rect 29092 32920 29144 32972
rect 32220 32963 32272 32972
rect 32220 32929 32229 32963
rect 32229 32929 32263 32963
rect 32263 32929 32272 32963
rect 32220 32920 32272 32929
rect 32772 32920 32824 32972
rect 36636 32988 36688 33040
rect 31760 32852 31812 32904
rect 32128 32895 32180 32904
rect 32128 32861 32137 32895
rect 32137 32861 32171 32895
rect 32171 32861 32180 32895
rect 32128 32852 32180 32861
rect 32680 32852 32732 32904
rect 37280 32920 37332 32972
rect 35808 32895 35860 32904
rect 35808 32861 35817 32895
rect 35817 32861 35851 32895
rect 35851 32861 35860 32895
rect 35808 32852 35860 32861
rect 35992 32895 36044 32904
rect 35992 32861 36001 32895
rect 36001 32861 36035 32895
rect 36035 32861 36044 32895
rect 35992 32852 36044 32861
rect 36820 32895 36872 32904
rect 21364 32716 21416 32768
rect 21824 32716 21876 32768
rect 23020 32716 23072 32768
rect 23112 32716 23164 32768
rect 23388 32716 23440 32768
rect 24492 32716 24544 32768
rect 36820 32861 36829 32895
rect 36829 32861 36863 32895
rect 36863 32861 36872 32895
rect 36820 32852 36872 32861
rect 37556 32895 37608 32904
rect 37556 32861 37565 32895
rect 37565 32861 37599 32895
rect 37599 32861 37608 32895
rect 37556 32852 37608 32861
rect 40224 32895 40276 32904
rect 40224 32861 40233 32895
rect 40233 32861 40267 32895
rect 40267 32861 40276 32895
rect 40224 32852 40276 32861
rect 36728 32784 36780 32836
rect 38660 32827 38712 32836
rect 38660 32793 38669 32827
rect 38669 32793 38703 32827
rect 38703 32793 38712 32827
rect 38660 32784 38712 32793
rect 38936 32784 38988 32836
rect 25964 32716 26016 32768
rect 31116 32716 31168 32768
rect 31300 32716 31352 32768
rect 31760 32716 31812 32768
rect 32772 32716 32824 32768
rect 33600 32759 33652 32768
rect 33600 32725 33609 32759
rect 33609 32725 33643 32759
rect 33643 32725 33652 32759
rect 33600 32716 33652 32725
rect 35624 32716 35676 32768
rect 37924 32716 37976 32768
rect 39028 32759 39080 32768
rect 39028 32725 39037 32759
rect 39037 32725 39071 32759
rect 39071 32725 39080 32759
rect 39028 32716 39080 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 19248 32512 19300 32564
rect 25504 32512 25556 32564
rect 25964 32555 26016 32564
rect 25964 32521 25973 32555
rect 25973 32521 26007 32555
rect 26007 32521 26016 32555
rect 25964 32512 26016 32521
rect 26332 32512 26384 32564
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 24860 32487 24912 32496
rect 24860 32453 24869 32487
rect 24869 32453 24903 32487
rect 24903 32453 24912 32487
rect 24860 32444 24912 32453
rect 25688 32444 25740 32496
rect 27252 32487 27304 32496
rect 27252 32453 27261 32487
rect 27261 32453 27295 32487
rect 27295 32453 27304 32487
rect 27252 32444 27304 32453
rect 28356 32444 28408 32496
rect 20444 32419 20496 32428
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 20628 32419 20680 32428
rect 20628 32385 20637 32419
rect 20637 32385 20671 32419
rect 20671 32385 20680 32419
rect 20628 32376 20680 32385
rect 22836 32376 22888 32428
rect 22928 32376 22980 32428
rect 15844 32351 15896 32360
rect 15844 32317 15853 32351
rect 15853 32317 15887 32351
rect 15887 32317 15896 32351
rect 15844 32308 15896 32317
rect 18236 32351 18288 32360
rect 18236 32317 18245 32351
rect 18245 32317 18279 32351
rect 18279 32317 18288 32351
rect 18236 32308 18288 32317
rect 23296 32308 23348 32360
rect 15200 32240 15252 32292
rect 15384 32215 15436 32224
rect 15384 32181 15393 32215
rect 15393 32181 15427 32215
rect 15427 32181 15436 32215
rect 15384 32172 15436 32181
rect 18604 32215 18656 32224
rect 18604 32181 18613 32215
rect 18613 32181 18647 32215
rect 18647 32181 18656 32215
rect 18604 32172 18656 32181
rect 19984 32172 20036 32224
rect 21364 32215 21416 32224
rect 21364 32181 21373 32215
rect 21373 32181 21407 32215
rect 21407 32181 21416 32215
rect 21364 32172 21416 32181
rect 21456 32172 21508 32224
rect 23480 32419 23532 32428
rect 23480 32385 23489 32419
rect 23489 32385 23523 32419
rect 23523 32385 23532 32419
rect 23480 32376 23532 32385
rect 23664 32419 23716 32428
rect 23664 32385 23673 32419
rect 23673 32385 23707 32419
rect 23707 32385 23716 32419
rect 23664 32376 23716 32385
rect 24676 32376 24728 32428
rect 25780 32419 25832 32428
rect 23572 32351 23624 32360
rect 23572 32317 23581 32351
rect 23581 32317 23615 32351
rect 23615 32317 23624 32351
rect 23572 32308 23624 32317
rect 24492 32351 24544 32360
rect 24492 32317 24501 32351
rect 24501 32317 24535 32351
rect 24535 32317 24544 32351
rect 24492 32308 24544 32317
rect 24768 32308 24820 32360
rect 25780 32385 25789 32419
rect 25789 32385 25823 32419
rect 25823 32385 25832 32419
rect 25780 32376 25832 32385
rect 26608 32376 26660 32428
rect 27436 32419 27488 32428
rect 27436 32385 27445 32419
rect 27445 32385 27479 32419
rect 27479 32385 27488 32419
rect 27436 32376 27488 32385
rect 27528 32419 27580 32428
rect 27528 32385 27537 32419
rect 27537 32385 27571 32419
rect 27571 32385 27580 32419
rect 28816 32419 28868 32428
rect 27528 32376 27580 32385
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 30288 32512 30340 32564
rect 29368 32376 29420 32428
rect 30656 32444 30708 32496
rect 29092 32308 29144 32360
rect 30380 32351 30432 32360
rect 30380 32317 30389 32351
rect 30389 32317 30423 32351
rect 30423 32317 30432 32351
rect 30380 32308 30432 32317
rect 25688 32240 25740 32292
rect 30472 32240 30524 32292
rect 31208 32376 31260 32428
rect 32680 32376 32732 32428
rect 33232 32376 33284 32428
rect 33600 32419 33652 32428
rect 33600 32385 33609 32419
rect 33609 32385 33643 32419
rect 33643 32385 33652 32419
rect 33600 32376 33652 32385
rect 33784 32376 33836 32428
rect 32128 32308 32180 32360
rect 33508 32308 33560 32360
rect 34060 32376 34112 32428
rect 33692 32240 33744 32292
rect 34428 32308 34480 32360
rect 35992 32512 36044 32564
rect 35716 32376 35768 32428
rect 37648 32419 37700 32428
rect 37648 32385 37657 32419
rect 37657 32385 37691 32419
rect 37691 32385 37700 32419
rect 37648 32376 37700 32385
rect 37924 32419 37976 32428
rect 37924 32385 37933 32419
rect 37933 32385 37967 32419
rect 37967 32385 37976 32419
rect 37924 32376 37976 32385
rect 38752 32444 38804 32496
rect 39672 32512 39724 32564
rect 39028 32376 39080 32428
rect 26976 32172 27028 32224
rect 27252 32215 27304 32224
rect 27252 32181 27261 32215
rect 27261 32181 27295 32215
rect 27295 32181 27304 32215
rect 27252 32172 27304 32181
rect 31116 32172 31168 32224
rect 33600 32172 33652 32224
rect 33876 32172 33928 32224
rect 35808 32172 35860 32224
rect 36452 32240 36504 32292
rect 37464 32215 37516 32224
rect 37464 32181 37473 32215
rect 37473 32181 37507 32215
rect 37507 32181 37516 32215
rect 37464 32172 37516 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 18236 31968 18288 32020
rect 23664 31968 23716 32020
rect 24676 31968 24728 32020
rect 26976 32011 27028 32020
rect 26976 31977 26985 32011
rect 26985 31977 27019 32011
rect 27019 31977 27028 32011
rect 26976 31968 27028 31977
rect 28356 32011 28408 32020
rect 28356 31977 28365 32011
rect 28365 31977 28399 32011
rect 28399 31977 28408 32011
rect 28356 31968 28408 31977
rect 30380 32011 30432 32020
rect 30380 31977 30389 32011
rect 30389 31977 30423 32011
rect 30423 31977 30432 32011
rect 30380 31968 30432 31977
rect 30472 31968 30524 32020
rect 16672 31875 16724 31884
rect 16672 31841 16681 31875
rect 16681 31841 16715 31875
rect 16715 31841 16724 31875
rect 16672 31832 16724 31841
rect 18052 31900 18104 31952
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 15384 31764 15436 31816
rect 17684 31832 17736 31884
rect 18604 31875 18656 31884
rect 18052 31807 18104 31816
rect 18052 31773 18061 31807
rect 18061 31773 18095 31807
rect 18095 31773 18104 31807
rect 18052 31764 18104 31773
rect 18604 31841 18613 31875
rect 18613 31841 18647 31875
rect 18647 31841 18656 31875
rect 18604 31832 18656 31841
rect 19984 31875 20036 31884
rect 19984 31841 19993 31875
rect 19993 31841 20027 31875
rect 20027 31841 20036 31875
rect 19984 31832 20036 31841
rect 20444 31875 20496 31884
rect 20444 31841 20453 31875
rect 20453 31841 20487 31875
rect 20487 31841 20496 31875
rect 20444 31832 20496 31841
rect 20904 31807 20956 31816
rect 14648 31696 14700 31748
rect 20904 31773 20913 31807
rect 20913 31773 20947 31807
rect 20947 31773 20956 31807
rect 20904 31764 20956 31773
rect 25780 31900 25832 31952
rect 26884 31943 26936 31952
rect 26884 31909 26893 31943
rect 26893 31909 26927 31943
rect 26927 31909 26936 31943
rect 26884 31900 26936 31909
rect 27252 31900 27304 31952
rect 35440 31968 35492 32020
rect 37648 32011 37700 32020
rect 37648 31977 37657 32011
rect 37657 31977 37691 32011
rect 37691 31977 37700 32011
rect 37648 31968 37700 31977
rect 25872 31832 25924 31884
rect 27160 31832 27212 31884
rect 21456 31764 21508 31816
rect 21732 31807 21784 31816
rect 21732 31773 21741 31807
rect 21741 31773 21775 31807
rect 21775 31773 21784 31807
rect 21732 31764 21784 31773
rect 22284 31764 22336 31816
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 24768 31807 24820 31816
rect 24768 31773 24777 31807
rect 24777 31773 24811 31807
rect 24811 31773 24820 31807
rect 24768 31764 24820 31773
rect 21640 31696 21692 31748
rect 24492 31696 24544 31748
rect 25320 31764 25372 31816
rect 25596 31764 25648 31816
rect 26332 31764 26384 31816
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 30564 31832 30616 31884
rect 31208 31875 31260 31884
rect 31208 31841 31217 31875
rect 31217 31841 31251 31875
rect 31251 31841 31260 31875
rect 31208 31832 31260 31841
rect 26976 31764 27028 31773
rect 25872 31696 25924 31748
rect 27068 31696 27120 31748
rect 27804 31739 27856 31748
rect 27804 31705 27813 31739
rect 27813 31705 27847 31739
rect 27847 31705 27856 31739
rect 27804 31696 27856 31705
rect 29184 31696 29236 31748
rect 31116 31764 31168 31816
rect 32956 31832 33008 31884
rect 32680 31807 32732 31816
rect 32680 31773 32689 31807
rect 32689 31773 32723 31807
rect 32723 31773 32732 31807
rect 32680 31764 32732 31773
rect 33784 31875 33836 31884
rect 33784 31841 33793 31875
rect 33793 31841 33827 31875
rect 33827 31841 33836 31875
rect 33784 31832 33836 31841
rect 33876 31875 33928 31884
rect 33876 31841 33885 31875
rect 33885 31841 33919 31875
rect 33919 31841 33928 31875
rect 33876 31832 33928 31841
rect 34060 31832 34112 31884
rect 36452 31875 36504 31884
rect 33508 31764 33560 31816
rect 35440 31807 35492 31816
rect 35440 31773 35449 31807
rect 35449 31773 35483 31807
rect 35483 31773 35492 31807
rect 35440 31764 35492 31773
rect 35624 31807 35676 31816
rect 35624 31773 35633 31807
rect 35633 31773 35667 31807
rect 35667 31773 35676 31807
rect 35624 31764 35676 31773
rect 36452 31841 36461 31875
rect 36461 31841 36495 31875
rect 36495 31841 36504 31875
rect 36452 31832 36504 31841
rect 37280 31807 37332 31816
rect 37280 31773 37289 31807
rect 37289 31773 37323 31807
rect 37323 31773 37332 31807
rect 37280 31764 37332 31773
rect 37556 31900 37608 31952
rect 18512 31671 18564 31680
rect 18512 31637 18521 31671
rect 18521 31637 18555 31671
rect 18555 31637 18564 31671
rect 18512 31628 18564 31637
rect 22744 31628 22796 31680
rect 26056 31628 26108 31680
rect 26516 31628 26568 31680
rect 28632 31628 28684 31680
rect 32588 31671 32640 31680
rect 32588 31637 32597 31671
rect 32597 31637 32631 31671
rect 32631 31637 32640 31671
rect 32588 31628 32640 31637
rect 34060 31671 34112 31680
rect 34060 31637 34069 31671
rect 34069 31637 34103 31671
rect 34103 31637 34112 31671
rect 34060 31628 34112 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 15844 31424 15896 31476
rect 21640 31424 21692 31476
rect 24492 31424 24544 31476
rect 26976 31424 27028 31476
rect 15200 31288 15252 31340
rect 16672 31356 16724 31408
rect 32680 31467 32732 31476
rect 32680 31433 32689 31467
rect 32689 31433 32723 31467
rect 32723 31433 32732 31467
rect 32680 31424 32732 31433
rect 27436 31399 27488 31408
rect 15936 31331 15988 31340
rect 15936 31297 15945 31331
rect 15945 31297 15979 31331
rect 15979 31297 15988 31331
rect 15936 31288 15988 31297
rect 16120 31288 16172 31340
rect 18236 31288 18288 31340
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 24768 31288 24820 31340
rect 27436 31365 27463 31399
rect 27463 31365 27488 31399
rect 27436 31356 27488 31365
rect 27620 31399 27672 31408
rect 27620 31365 27629 31399
rect 27629 31365 27663 31399
rect 27663 31365 27672 31399
rect 27620 31356 27672 31365
rect 25872 31331 25924 31340
rect 25872 31297 25881 31331
rect 25881 31297 25915 31331
rect 25915 31297 25924 31331
rect 25872 31288 25924 31297
rect 26056 31331 26108 31340
rect 26056 31297 26065 31331
rect 26065 31297 26099 31331
rect 26099 31297 26108 31331
rect 26056 31288 26108 31297
rect 31392 31356 31444 31408
rect 32956 31356 33008 31408
rect 34060 31424 34112 31476
rect 34244 31356 34296 31408
rect 15292 31220 15344 31272
rect 17684 31263 17736 31272
rect 17684 31229 17693 31263
rect 17693 31229 17727 31263
rect 17727 31229 17736 31263
rect 17684 31220 17736 31229
rect 18420 31220 18472 31272
rect 25964 31263 26016 31272
rect 25964 31229 25973 31263
rect 25973 31229 26007 31263
rect 26007 31229 26016 31263
rect 25964 31220 26016 31229
rect 28632 31288 28684 31340
rect 29184 31331 29236 31340
rect 29184 31297 29193 31331
rect 29193 31297 29227 31331
rect 29227 31297 29236 31331
rect 29184 31288 29236 31297
rect 29644 31288 29696 31340
rect 31024 31331 31076 31340
rect 31024 31297 31033 31331
rect 31033 31297 31067 31331
rect 31067 31297 31076 31331
rect 31024 31288 31076 31297
rect 31484 31288 31536 31340
rect 35348 31331 35400 31340
rect 35348 31297 35357 31331
rect 35357 31297 35391 31331
rect 35391 31297 35400 31331
rect 35348 31288 35400 31297
rect 35900 31288 35952 31340
rect 28540 31263 28592 31272
rect 28540 31229 28549 31263
rect 28549 31229 28583 31263
rect 28583 31229 28592 31263
rect 28540 31220 28592 31229
rect 30104 31263 30156 31272
rect 30104 31229 30113 31263
rect 30113 31229 30147 31263
rect 30147 31229 30156 31263
rect 30104 31220 30156 31229
rect 33968 31220 34020 31272
rect 34796 31220 34848 31272
rect 18880 31152 18932 31204
rect 57428 31152 57480 31204
rect 16948 31084 17000 31136
rect 22560 31084 22612 31136
rect 24584 31127 24636 31136
rect 24584 31093 24593 31127
rect 24593 31093 24627 31127
rect 24627 31093 24636 31127
rect 24584 31084 24636 31093
rect 27160 31084 27212 31136
rect 28356 31084 28408 31136
rect 32956 31084 33008 31136
rect 34336 31127 34388 31136
rect 34336 31093 34345 31127
rect 34345 31093 34379 31127
rect 34379 31093 34388 31127
rect 34336 31084 34388 31093
rect 35992 31084 36044 31136
rect 37188 31084 37240 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15200 30880 15252 30932
rect 15936 30880 15988 30932
rect 20444 30880 20496 30932
rect 25964 30923 26016 30932
rect 25964 30889 25973 30923
rect 25973 30889 26007 30923
rect 26007 30889 26016 30923
rect 25964 30880 26016 30889
rect 26884 30880 26936 30932
rect 22284 30812 22336 30864
rect 24768 30812 24820 30864
rect 16120 30787 16172 30796
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 17960 30787 18012 30796
rect 17960 30753 17969 30787
rect 17969 30753 18003 30787
rect 18003 30753 18012 30787
rect 17960 30744 18012 30753
rect 16672 30676 16724 30728
rect 20260 30744 20312 30796
rect 18880 30719 18932 30728
rect 18880 30685 18889 30719
rect 18889 30685 18923 30719
rect 18923 30685 18932 30719
rect 18880 30676 18932 30685
rect 20168 30676 20220 30728
rect 20536 30651 20588 30660
rect 19432 30540 19484 30592
rect 20536 30617 20563 30651
rect 20563 30617 20588 30651
rect 20536 30608 20588 30617
rect 20720 30651 20772 30660
rect 20720 30617 20729 30651
rect 20729 30617 20763 30651
rect 20763 30617 20772 30651
rect 24308 30744 24360 30796
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 22560 30719 22612 30728
rect 22560 30685 22569 30719
rect 22569 30685 22603 30719
rect 22603 30685 22612 30719
rect 22560 30676 22612 30685
rect 22744 30719 22796 30728
rect 22744 30685 22753 30719
rect 22753 30685 22787 30719
rect 22787 30685 22796 30719
rect 22744 30676 22796 30685
rect 20720 30608 20772 30617
rect 22100 30651 22152 30660
rect 22100 30617 22109 30651
rect 22109 30617 22143 30651
rect 22143 30617 22152 30651
rect 22100 30608 22152 30617
rect 20996 30540 21048 30592
rect 24676 30676 24728 30728
rect 25688 30744 25740 30796
rect 29184 30880 29236 30932
rect 31484 30923 31536 30932
rect 31484 30889 31493 30923
rect 31493 30889 31527 30923
rect 31527 30889 31536 30923
rect 31484 30880 31536 30889
rect 34152 30923 34204 30932
rect 34152 30889 34161 30923
rect 34161 30889 34195 30923
rect 34195 30889 34204 30923
rect 34152 30880 34204 30889
rect 35348 30880 35400 30932
rect 36452 30880 36504 30932
rect 25320 30676 25372 30728
rect 26424 30719 26476 30728
rect 26424 30685 26433 30719
rect 26433 30685 26467 30719
rect 26467 30685 26476 30719
rect 26424 30676 26476 30685
rect 26976 30676 27028 30728
rect 28264 30719 28316 30728
rect 26516 30608 26568 30660
rect 28264 30685 28273 30719
rect 28273 30685 28307 30719
rect 28307 30685 28316 30719
rect 28264 30676 28316 30685
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 28724 30676 28776 30728
rect 32128 30812 32180 30864
rect 32496 30812 32548 30864
rect 30840 30744 30892 30796
rect 31024 30744 31076 30796
rect 31392 30719 31444 30728
rect 31392 30685 31401 30719
rect 31401 30685 31435 30719
rect 31435 30685 31444 30719
rect 31392 30676 31444 30685
rect 32588 30676 32640 30728
rect 32956 30719 33008 30728
rect 32956 30685 32965 30719
rect 32965 30685 32999 30719
rect 32999 30685 33008 30719
rect 32956 30676 33008 30685
rect 34244 30744 34296 30796
rect 33968 30676 34020 30728
rect 26332 30540 26384 30592
rect 26884 30540 26936 30592
rect 27068 30540 27120 30592
rect 27436 30540 27488 30592
rect 27804 30583 27856 30592
rect 27804 30549 27813 30583
rect 27813 30549 27847 30583
rect 27847 30549 27856 30583
rect 27804 30540 27856 30549
rect 28448 30540 28500 30592
rect 33600 30608 33652 30660
rect 35716 30719 35768 30728
rect 35716 30685 35725 30719
rect 35725 30685 35759 30719
rect 35759 30685 35768 30719
rect 36084 30744 36136 30796
rect 37280 30787 37332 30796
rect 37280 30753 37289 30787
rect 37289 30753 37323 30787
rect 37323 30753 37332 30787
rect 37280 30744 37332 30753
rect 41328 30744 41380 30796
rect 35716 30676 35768 30685
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 37188 30719 37240 30728
rect 35992 30676 36044 30685
rect 37188 30685 37197 30719
rect 37197 30685 37231 30719
rect 37231 30685 37240 30719
rect 37188 30676 37240 30685
rect 29276 30540 29328 30592
rect 29552 30540 29604 30592
rect 30932 30583 30984 30592
rect 30932 30549 30941 30583
rect 30941 30549 30975 30583
rect 30975 30549 30984 30583
rect 30932 30540 30984 30549
rect 35900 30540 35952 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 17960 30379 18012 30388
rect 17960 30345 17969 30379
rect 17969 30345 18003 30379
rect 18003 30345 18012 30379
rect 17960 30336 18012 30345
rect 20444 30336 20496 30388
rect 26240 30379 26292 30388
rect 26240 30345 26249 30379
rect 26249 30345 26283 30379
rect 26283 30345 26292 30379
rect 26240 30336 26292 30345
rect 26424 30336 26476 30388
rect 27528 30336 27580 30388
rect 28632 30336 28684 30388
rect 18052 30200 18104 30252
rect 18512 30200 18564 30252
rect 19432 30200 19484 30252
rect 20720 30268 20772 30320
rect 20536 30200 20588 30252
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 20996 30243 21048 30252
rect 20996 30209 21005 30243
rect 21005 30209 21039 30243
rect 21039 30209 21048 30243
rect 20996 30200 21048 30209
rect 22560 30200 22612 30252
rect 23940 30200 23992 30252
rect 24216 30200 24268 30252
rect 24584 30200 24636 30252
rect 24768 30200 24820 30252
rect 20812 30132 20864 30184
rect 22652 30175 22704 30184
rect 22652 30141 22661 30175
rect 22661 30141 22695 30175
rect 22695 30141 22704 30175
rect 22652 30132 22704 30141
rect 27068 30268 27120 30320
rect 26332 30200 26384 30252
rect 26608 30200 26660 30252
rect 20168 30107 20220 30116
rect 20168 30073 20177 30107
rect 20177 30073 20211 30107
rect 20211 30073 20220 30107
rect 20168 30064 20220 30073
rect 23756 30064 23808 30116
rect 27620 30132 27672 30184
rect 28448 30243 28500 30252
rect 28448 30209 28457 30243
rect 28457 30209 28491 30243
rect 28491 30209 28500 30243
rect 29368 30311 29420 30320
rect 29368 30277 29377 30311
rect 29377 30277 29411 30311
rect 29411 30277 29420 30311
rect 29368 30268 29420 30277
rect 34796 30336 34848 30388
rect 33968 30311 34020 30320
rect 28448 30200 28500 30209
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 29000 30132 29052 30184
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 32772 30243 32824 30252
rect 32772 30209 32781 30243
rect 32781 30209 32815 30243
rect 32815 30209 32824 30243
rect 32772 30200 32824 30209
rect 32128 30132 32180 30184
rect 33968 30277 33977 30311
rect 33977 30277 34011 30311
rect 34011 30277 34020 30311
rect 33968 30268 34020 30277
rect 34152 30311 34204 30320
rect 34152 30277 34193 30311
rect 34193 30277 34204 30311
rect 34152 30268 34204 30277
rect 35440 30268 35492 30320
rect 35992 30268 36044 30320
rect 34060 30200 34112 30252
rect 35900 30243 35952 30252
rect 34336 30132 34388 30184
rect 35900 30209 35909 30243
rect 35909 30209 35943 30243
rect 35943 30209 35952 30243
rect 35900 30200 35952 30209
rect 36084 30243 36136 30252
rect 36084 30209 36093 30243
rect 36093 30209 36127 30243
rect 36127 30209 36136 30243
rect 36084 30200 36136 30209
rect 21088 30039 21140 30048
rect 21088 30005 21097 30039
rect 21097 30005 21131 30039
rect 21131 30005 21140 30039
rect 21088 29996 21140 30005
rect 21732 29996 21784 30048
rect 25320 29996 25372 30048
rect 37280 30268 37332 30320
rect 36636 30243 36688 30252
rect 36636 30209 36645 30243
rect 36645 30209 36679 30243
rect 36679 30209 36688 30243
rect 36636 30200 36688 30209
rect 28908 30039 28960 30048
rect 28908 30005 28917 30039
rect 28917 30005 28951 30039
rect 28951 30005 28960 30039
rect 28908 29996 28960 30005
rect 32496 29996 32548 30048
rect 33600 29996 33652 30048
rect 36084 30064 36136 30116
rect 36636 30064 36688 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 20996 29792 21048 29844
rect 22100 29792 22152 29844
rect 27528 29792 27580 29844
rect 29092 29792 29144 29844
rect 31300 29792 31352 29844
rect 33692 29792 33744 29844
rect 18512 29724 18564 29776
rect 21088 29724 21140 29776
rect 24768 29724 24820 29776
rect 20904 29656 20956 29708
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 25044 29656 25096 29708
rect 34060 29724 34112 29776
rect 19432 29588 19484 29640
rect 20076 29588 20128 29640
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 21732 29631 21784 29640
rect 21732 29597 21741 29631
rect 21741 29597 21775 29631
rect 21775 29597 21784 29631
rect 21732 29588 21784 29597
rect 22468 29588 22520 29640
rect 22652 29588 22704 29640
rect 24584 29588 24636 29640
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 26884 29631 26936 29640
rect 26884 29597 26893 29631
rect 26893 29597 26927 29631
rect 26927 29597 26936 29631
rect 26884 29588 26936 29597
rect 29000 29656 29052 29708
rect 29276 29656 29328 29708
rect 28908 29588 28960 29640
rect 29644 29588 29696 29640
rect 30104 29588 30156 29640
rect 20628 29520 20680 29572
rect 30840 29563 30892 29572
rect 30840 29529 30849 29563
rect 30849 29529 30883 29563
rect 30883 29529 30892 29563
rect 30840 29520 30892 29529
rect 19340 29452 19392 29504
rect 19984 29452 20036 29504
rect 20812 29452 20864 29504
rect 23848 29495 23900 29504
rect 23848 29461 23857 29495
rect 23857 29461 23891 29495
rect 23891 29461 23900 29495
rect 23848 29452 23900 29461
rect 24124 29452 24176 29504
rect 31576 29520 31628 29572
rect 33416 29656 33468 29708
rect 33048 29588 33100 29640
rect 31300 29495 31352 29504
rect 31300 29461 31309 29495
rect 31309 29461 31343 29495
rect 31343 29461 31352 29495
rect 31300 29452 31352 29461
rect 32404 29452 32456 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 24124 29248 24176 29300
rect 25964 29248 26016 29300
rect 29000 29291 29052 29300
rect 29000 29257 29009 29291
rect 29009 29257 29043 29291
rect 29043 29257 29052 29291
rect 29000 29248 29052 29257
rect 16948 29223 17000 29232
rect 16948 29189 16957 29223
rect 16957 29189 16991 29223
rect 16991 29189 17000 29223
rect 16948 29180 17000 29189
rect 18052 29044 18104 29096
rect 18512 29180 18564 29232
rect 20904 29223 20956 29232
rect 20904 29189 20913 29223
rect 20913 29189 20947 29223
rect 20947 29189 20956 29223
rect 20904 29180 20956 29189
rect 25136 29180 25188 29232
rect 33140 29248 33192 29300
rect 30840 29180 30892 29232
rect 30932 29223 30984 29232
rect 30932 29189 30941 29223
rect 30941 29189 30975 29223
rect 30975 29189 30984 29223
rect 30932 29180 30984 29189
rect 19984 29155 20036 29164
rect 19432 29044 19484 29096
rect 19984 29121 19993 29155
rect 19993 29121 20027 29155
rect 20027 29121 20036 29155
rect 19984 29112 20036 29121
rect 20076 29155 20128 29164
rect 20076 29121 20085 29155
rect 20085 29121 20119 29155
rect 20119 29121 20128 29155
rect 20076 29112 20128 29121
rect 20812 29112 20864 29164
rect 21364 29112 21416 29164
rect 23756 29155 23808 29164
rect 20996 29044 21048 29096
rect 1676 29019 1728 29028
rect 1676 28985 1685 29019
rect 1685 28985 1719 29019
rect 1719 28985 1728 29019
rect 1676 28976 1728 28985
rect 18880 28976 18932 29028
rect 19616 28976 19668 29028
rect 17868 28951 17920 28960
rect 17868 28917 17877 28951
rect 17877 28917 17911 28951
rect 17911 28917 17920 28951
rect 17868 28908 17920 28917
rect 19432 28908 19484 28960
rect 20260 28976 20312 29028
rect 20628 29019 20680 29028
rect 20628 28985 20637 29019
rect 20637 28985 20671 29019
rect 20671 28985 20680 29019
rect 20628 28976 20680 28985
rect 23756 29121 23765 29155
rect 23765 29121 23799 29155
rect 23799 29121 23808 29155
rect 23756 29112 23808 29121
rect 25320 29112 25372 29164
rect 27436 29112 27488 29164
rect 24308 29087 24360 29096
rect 24308 29053 24317 29087
rect 24317 29053 24351 29087
rect 24351 29053 24360 29087
rect 24308 29044 24360 29053
rect 26976 29044 27028 29096
rect 27528 29087 27580 29096
rect 27528 29053 27537 29087
rect 27537 29053 27571 29087
rect 27571 29053 27580 29087
rect 27528 29044 27580 29053
rect 27620 29044 27672 29096
rect 28540 29155 28592 29164
rect 28540 29121 28549 29155
rect 28549 29121 28583 29155
rect 28583 29121 28592 29155
rect 28540 29112 28592 29121
rect 29644 29155 29696 29164
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 30104 29112 30156 29164
rect 28172 29044 28224 29096
rect 31300 29112 31352 29164
rect 31484 29180 31536 29232
rect 34060 29223 34112 29232
rect 34060 29189 34069 29223
rect 34069 29189 34103 29223
rect 34103 29189 34112 29223
rect 34060 29180 34112 29189
rect 37188 29180 37240 29232
rect 23848 28976 23900 29028
rect 26240 28976 26292 29028
rect 29828 28976 29880 29028
rect 32312 29044 32364 29096
rect 33784 29087 33836 29096
rect 33784 29053 33793 29087
rect 33793 29053 33827 29087
rect 33827 29053 33836 29087
rect 33784 29044 33836 29053
rect 36084 29112 36136 29164
rect 32680 28976 32732 29028
rect 35532 29044 35584 29096
rect 57888 28976 57940 29028
rect 23572 28908 23624 28960
rect 25136 28908 25188 28960
rect 30104 28951 30156 28960
rect 30104 28917 30113 28951
rect 30113 28917 30147 28951
rect 30147 28917 30156 28951
rect 30104 28908 30156 28917
rect 30380 28908 30432 28960
rect 32588 28908 32640 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19616 28747 19668 28756
rect 19616 28713 19625 28747
rect 19625 28713 19659 28747
rect 19659 28713 19668 28747
rect 19616 28704 19668 28713
rect 16948 28636 17000 28688
rect 18880 28543 18932 28552
rect 18880 28509 18889 28543
rect 18889 28509 18923 28543
rect 18923 28509 18932 28543
rect 18880 28500 18932 28509
rect 19248 28500 19300 28552
rect 25596 28636 25648 28688
rect 20628 28611 20680 28620
rect 20628 28577 20637 28611
rect 20637 28577 20671 28611
rect 20671 28577 20680 28611
rect 20628 28568 20680 28577
rect 23572 28611 23624 28620
rect 22284 28543 22336 28552
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 22468 28543 22520 28552
rect 22468 28509 22477 28543
rect 22477 28509 22511 28543
rect 22511 28509 22520 28543
rect 23572 28577 23581 28611
rect 23581 28577 23615 28611
rect 23615 28577 23624 28611
rect 23572 28568 23624 28577
rect 26240 28611 26292 28620
rect 26240 28577 26249 28611
rect 26249 28577 26283 28611
rect 26283 28577 26292 28611
rect 26240 28568 26292 28577
rect 31484 28636 31536 28688
rect 22468 28500 22520 28509
rect 25044 28500 25096 28552
rect 27620 28543 27672 28552
rect 27620 28509 27629 28543
rect 27629 28509 27663 28543
rect 27663 28509 27672 28543
rect 27620 28500 27672 28509
rect 28172 28543 28224 28552
rect 17868 28432 17920 28484
rect 20904 28432 20956 28484
rect 20996 28475 21048 28484
rect 20996 28441 21005 28475
rect 21005 28441 21039 28475
rect 21039 28441 21048 28475
rect 25136 28475 25188 28484
rect 20996 28432 21048 28441
rect 25136 28441 25145 28475
rect 25145 28441 25179 28475
rect 25179 28441 25188 28475
rect 25136 28432 25188 28441
rect 28172 28509 28181 28543
rect 28181 28509 28215 28543
rect 28215 28509 28224 28543
rect 28172 28500 28224 28509
rect 28540 28500 28592 28552
rect 29092 28500 29144 28552
rect 30748 28500 30800 28552
rect 30932 28543 30984 28552
rect 30932 28509 30941 28543
rect 30941 28509 30975 28543
rect 30975 28509 30984 28543
rect 32496 28543 32548 28552
rect 30932 28500 30984 28509
rect 32496 28509 32505 28543
rect 32505 28509 32539 28543
rect 32539 28509 32548 28543
rect 32496 28500 32548 28509
rect 32772 28543 32824 28552
rect 32772 28509 32781 28543
rect 32781 28509 32815 28543
rect 32815 28509 32824 28543
rect 32772 28500 32824 28509
rect 33784 28500 33836 28552
rect 33968 28500 34020 28552
rect 18604 28407 18656 28416
rect 18604 28373 18613 28407
rect 18613 28373 18647 28407
rect 18647 28373 18656 28407
rect 18604 28364 18656 28373
rect 22284 28364 22336 28416
rect 25412 28364 25464 28416
rect 26976 28407 27028 28416
rect 26976 28373 26985 28407
rect 26985 28373 27019 28407
rect 27019 28373 27028 28407
rect 26976 28364 27028 28373
rect 27528 28364 27580 28416
rect 29184 28432 29236 28484
rect 30104 28432 30156 28484
rect 33600 28432 33652 28484
rect 35532 28475 35584 28484
rect 35532 28441 35541 28475
rect 35541 28441 35575 28475
rect 35575 28441 35584 28475
rect 35532 28432 35584 28441
rect 37188 28432 37240 28484
rect 31116 28364 31168 28416
rect 36544 28364 36596 28416
rect 39488 28432 39540 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 19340 28092 19392 28144
rect 22192 28092 22244 28144
rect 9864 28024 9916 28076
rect 20904 28067 20956 28076
rect 20904 28033 20913 28067
rect 20913 28033 20947 28067
rect 20947 28033 20956 28067
rect 20904 28024 20956 28033
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 22468 28092 22520 28144
rect 28540 28160 28592 28212
rect 25136 28024 25188 28076
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 27620 28092 27672 28144
rect 29000 28092 29052 28144
rect 29184 28092 29236 28144
rect 31116 28135 31168 28144
rect 31116 28101 31125 28135
rect 31125 28101 31159 28135
rect 31159 28101 31168 28135
rect 31116 28092 31168 28101
rect 34152 28092 34204 28144
rect 34704 28092 34756 28144
rect 27528 28024 27580 28076
rect 33140 28067 33192 28076
rect 33140 28033 33149 28067
rect 33149 28033 33183 28067
rect 33183 28033 33192 28067
rect 33140 28024 33192 28033
rect 33600 28067 33652 28076
rect 33600 28033 33609 28067
rect 33609 28033 33643 28067
rect 33643 28033 33652 28067
rect 33600 28024 33652 28033
rect 34796 28067 34848 28076
rect 34796 28033 34805 28067
rect 34805 28033 34839 28067
rect 34839 28033 34848 28067
rect 34796 28024 34848 28033
rect 19248 27999 19300 28008
rect 19248 27965 19257 27999
rect 19257 27965 19291 27999
rect 19291 27965 19300 27999
rect 19248 27956 19300 27965
rect 19432 27956 19484 28008
rect 27252 27956 27304 28008
rect 31760 27956 31812 28008
rect 32404 27956 32456 28008
rect 35624 28024 35676 28076
rect 35348 27956 35400 28008
rect 21364 27820 21416 27872
rect 25596 27820 25648 27872
rect 29828 27820 29880 27872
rect 35440 27863 35492 27872
rect 35440 27829 35449 27863
rect 35449 27829 35483 27863
rect 35483 27829 35492 27863
rect 35440 27820 35492 27829
rect 36452 27863 36504 27872
rect 36452 27829 36461 27863
rect 36461 27829 36495 27863
rect 36495 27829 36504 27863
rect 36452 27820 36504 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 28172 27616 28224 27668
rect 35440 27616 35492 27668
rect 2872 27548 2924 27600
rect 22192 27480 22244 27532
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 22468 27412 22520 27464
rect 24032 27412 24084 27464
rect 25136 27412 25188 27464
rect 25596 27455 25648 27464
rect 25596 27421 25605 27455
rect 25605 27421 25639 27455
rect 25639 27421 25648 27455
rect 26976 27548 27028 27600
rect 30380 27548 30432 27600
rect 30748 27591 30800 27600
rect 30748 27557 30757 27591
rect 30757 27557 30791 27591
rect 30791 27557 30800 27591
rect 30748 27548 30800 27557
rect 33232 27548 33284 27600
rect 25596 27412 25648 27421
rect 19340 27344 19392 27396
rect 24584 27387 24636 27396
rect 20904 27276 20956 27328
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 26976 27276 27028 27328
rect 27436 27276 27488 27328
rect 28172 27276 28224 27328
rect 31024 27412 31076 27464
rect 31300 27455 31352 27464
rect 31300 27421 31309 27455
rect 31309 27421 31343 27455
rect 31343 27421 31352 27455
rect 31300 27412 31352 27421
rect 31484 27319 31536 27328
rect 31484 27285 31493 27319
rect 31493 27285 31527 27319
rect 31527 27285 31536 27319
rect 31484 27276 31536 27285
rect 31944 27276 31996 27328
rect 35900 27455 35952 27464
rect 35900 27421 35909 27455
rect 35909 27421 35943 27455
rect 35943 27421 35952 27455
rect 35900 27412 35952 27421
rect 33232 27319 33284 27328
rect 33232 27285 33241 27319
rect 33241 27285 33275 27319
rect 33275 27285 33284 27319
rect 33232 27276 33284 27285
rect 33784 27276 33836 27328
rect 34244 27319 34296 27328
rect 34244 27285 34253 27319
rect 34253 27285 34287 27319
rect 34287 27285 34296 27319
rect 34244 27276 34296 27285
rect 34704 27276 34756 27328
rect 35348 27344 35400 27396
rect 37188 27344 37240 27396
rect 37924 27387 37976 27396
rect 37924 27353 37933 27387
rect 37933 27353 37967 27387
rect 37967 27353 37976 27387
rect 37924 27344 37976 27353
rect 38384 27387 38436 27396
rect 38384 27353 38393 27387
rect 38393 27353 38427 27387
rect 38427 27353 38436 27387
rect 38384 27344 38436 27353
rect 36452 27276 36504 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 20996 27004 21048 27056
rect 24584 27072 24636 27124
rect 23388 27004 23440 27056
rect 27160 27072 27212 27124
rect 27436 27047 27488 27056
rect 27436 27013 27445 27047
rect 27445 27013 27479 27047
rect 27479 27013 27488 27047
rect 27436 27004 27488 27013
rect 27528 27004 27580 27056
rect 31208 27004 31260 27056
rect 31484 27047 31536 27056
rect 31484 27013 31493 27047
rect 31493 27013 31527 27047
rect 31527 27013 31536 27047
rect 31484 27004 31536 27013
rect 34612 27072 34664 27124
rect 34244 27004 34296 27056
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 31760 26979 31812 26988
rect 31760 26945 31769 26979
rect 31769 26945 31803 26979
rect 31803 26945 31812 26979
rect 31760 26936 31812 26945
rect 33784 26979 33836 26988
rect 33784 26945 33793 26979
rect 33793 26945 33827 26979
rect 33827 26945 33836 26979
rect 33784 26936 33836 26945
rect 33968 26979 34020 26988
rect 33968 26945 33977 26979
rect 33977 26945 34011 26979
rect 34011 26945 34020 26979
rect 33968 26936 34020 26945
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 35532 27072 35584 27124
rect 36912 27072 36964 27124
rect 37188 27072 37240 27124
rect 39488 27115 39540 27124
rect 39488 27081 39497 27115
rect 39497 27081 39531 27115
rect 39531 27081 39540 27115
rect 39488 27072 39540 27081
rect 20444 26911 20496 26920
rect 20444 26877 20453 26911
rect 20453 26877 20487 26911
rect 20487 26877 20496 26911
rect 20444 26868 20496 26877
rect 24584 26868 24636 26920
rect 27160 26911 27212 26920
rect 27160 26877 27169 26911
rect 27169 26877 27203 26911
rect 27203 26877 27212 26911
rect 27160 26868 27212 26877
rect 35440 26936 35492 26988
rect 38384 26936 38436 26988
rect 35532 26868 35584 26920
rect 38844 26868 38896 26920
rect 43996 26868 44048 26920
rect 57612 26868 57664 26920
rect 33784 26800 33836 26852
rect 34060 26800 34112 26852
rect 39488 26800 39540 26852
rect 57152 26800 57204 26852
rect 24216 26732 24268 26784
rect 29460 26732 29512 26784
rect 33232 26732 33284 26784
rect 35900 26732 35952 26784
rect 36820 26775 36872 26784
rect 36820 26741 36829 26775
rect 36829 26741 36863 26775
rect 36863 26741 36872 26775
rect 36820 26732 36872 26741
rect 38752 26732 38804 26784
rect 41880 26775 41932 26784
rect 41880 26741 41889 26775
rect 41889 26741 41923 26775
rect 41923 26741 41932 26775
rect 41880 26732 41932 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 23388 26528 23440 26580
rect 23848 26528 23900 26580
rect 27436 26460 27488 26512
rect 24584 26435 24636 26444
rect 24584 26401 24593 26435
rect 24593 26401 24627 26435
rect 24627 26401 24636 26435
rect 24584 26392 24636 26401
rect 26332 26392 26384 26444
rect 26792 26392 26844 26444
rect 24124 26324 24176 26376
rect 27068 26324 27120 26376
rect 31300 26528 31352 26580
rect 33416 26571 33468 26580
rect 33416 26537 33425 26571
rect 33425 26537 33459 26571
rect 33459 26537 33468 26571
rect 33416 26528 33468 26537
rect 34796 26528 34848 26580
rect 35348 26528 35400 26580
rect 30472 26435 30524 26444
rect 30472 26401 30481 26435
rect 30481 26401 30515 26435
rect 30515 26401 30524 26435
rect 30472 26392 30524 26401
rect 36176 26528 36228 26580
rect 37188 26528 37240 26580
rect 58164 26528 58216 26580
rect 40224 26460 40276 26512
rect 33968 26392 34020 26444
rect 33232 26367 33284 26376
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33232 26324 33284 26333
rect 24216 26256 24268 26308
rect 27344 26256 27396 26308
rect 31208 26256 31260 26308
rect 32588 26256 32640 26308
rect 34336 26324 34388 26376
rect 30656 26188 30708 26240
rect 34796 26256 34848 26308
rect 37280 26392 37332 26444
rect 38384 26392 38436 26444
rect 39212 26367 39264 26376
rect 39212 26333 39221 26367
rect 39221 26333 39255 26367
rect 39255 26333 39264 26367
rect 39212 26324 39264 26333
rect 40040 26324 40092 26376
rect 41880 26324 41932 26376
rect 36084 26299 36136 26308
rect 36084 26265 36093 26299
rect 36093 26265 36127 26299
rect 36127 26265 36136 26299
rect 36084 26256 36136 26265
rect 38016 26256 38068 26308
rect 38752 26256 38804 26308
rect 41052 26256 41104 26308
rect 33876 26188 33928 26240
rect 35900 26188 35952 26240
rect 40132 26188 40184 26240
rect 43444 26256 43496 26308
rect 44824 26188 44876 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 24124 26027 24176 26036
rect 24124 25993 24133 26027
rect 24133 25993 24167 26027
rect 24167 25993 24176 26027
rect 24124 25984 24176 25993
rect 27160 25984 27212 26036
rect 30472 25984 30524 26036
rect 33416 25984 33468 26036
rect 33876 25984 33928 26036
rect 29460 25959 29512 25968
rect 29460 25925 29469 25959
rect 29469 25925 29503 25959
rect 29503 25925 29512 25959
rect 29460 25916 29512 25925
rect 31208 25916 31260 25968
rect 27528 25848 27580 25900
rect 33600 25891 33652 25900
rect 33600 25857 33609 25891
rect 33609 25857 33643 25891
rect 33643 25857 33652 25891
rect 33600 25848 33652 25857
rect 26332 25823 26384 25832
rect 26332 25789 26341 25823
rect 26341 25789 26375 25823
rect 26375 25789 26384 25823
rect 26332 25780 26384 25789
rect 27252 25780 27304 25832
rect 27068 25644 27120 25696
rect 33416 25780 33468 25832
rect 34244 25712 34296 25764
rect 35440 25984 35492 26036
rect 36084 25984 36136 26036
rect 39212 25984 39264 26036
rect 41052 26027 41104 26036
rect 41052 25993 41061 26027
rect 41061 25993 41095 26027
rect 41095 25993 41104 26027
rect 41052 25984 41104 25993
rect 35440 25891 35492 25900
rect 35440 25857 35449 25891
rect 35449 25857 35483 25891
rect 35483 25857 35492 25891
rect 35440 25848 35492 25857
rect 35532 25891 35584 25900
rect 35532 25857 35541 25891
rect 35541 25857 35575 25891
rect 35575 25857 35584 25891
rect 42800 25916 42852 25968
rect 43628 25916 43680 25968
rect 35532 25848 35584 25857
rect 39488 25891 39540 25900
rect 39488 25857 39497 25891
rect 39497 25857 39531 25891
rect 39531 25857 39540 25891
rect 39488 25848 39540 25857
rect 40132 25891 40184 25900
rect 40132 25857 40141 25891
rect 40141 25857 40175 25891
rect 40175 25857 40184 25891
rect 40132 25848 40184 25857
rect 42064 25848 42116 25900
rect 43444 25891 43496 25900
rect 43444 25857 43453 25891
rect 43453 25857 43487 25891
rect 43487 25857 43496 25891
rect 43444 25848 43496 25857
rect 43536 25891 43588 25900
rect 43536 25857 43545 25891
rect 43545 25857 43579 25891
rect 43579 25857 43588 25891
rect 43536 25848 43588 25857
rect 44824 25848 44876 25900
rect 46112 25848 46164 25900
rect 38016 25780 38068 25832
rect 38384 25712 38436 25764
rect 41144 25712 41196 25764
rect 27528 25644 27580 25696
rect 30656 25644 30708 25696
rect 30932 25687 30984 25696
rect 30932 25653 30941 25687
rect 30941 25653 30975 25687
rect 30975 25653 30984 25687
rect 30932 25644 30984 25653
rect 33140 25644 33192 25696
rect 39948 25644 40000 25696
rect 41052 25644 41104 25696
rect 41972 25687 42024 25696
rect 41972 25653 41981 25687
rect 41981 25653 42015 25687
rect 42015 25653 42024 25687
rect 41972 25644 42024 25653
rect 43352 25644 43404 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 27528 25483 27580 25492
rect 27528 25449 27537 25483
rect 27537 25449 27571 25483
rect 27571 25449 27580 25483
rect 27528 25440 27580 25449
rect 33600 25440 33652 25492
rect 33876 25483 33928 25492
rect 33876 25449 33885 25483
rect 33885 25449 33919 25483
rect 33919 25449 33928 25483
rect 33876 25440 33928 25449
rect 30932 25415 30984 25424
rect 30932 25381 30941 25415
rect 30941 25381 30975 25415
rect 30975 25381 30984 25415
rect 30932 25372 30984 25381
rect 33140 25347 33192 25356
rect 33140 25313 33149 25347
rect 33149 25313 33183 25347
rect 33183 25313 33192 25347
rect 33140 25304 33192 25313
rect 33968 25372 34020 25424
rect 35808 25440 35860 25492
rect 39212 25440 39264 25492
rect 41052 25483 41104 25492
rect 41052 25449 41061 25483
rect 41061 25449 41095 25483
rect 41095 25449 41104 25483
rect 41052 25440 41104 25449
rect 30472 25279 30524 25288
rect 30472 25245 30481 25279
rect 30481 25245 30515 25279
rect 30515 25245 30524 25279
rect 30472 25236 30524 25245
rect 33416 25279 33468 25288
rect 33416 25245 33425 25279
rect 33425 25245 33459 25279
rect 33459 25245 33468 25279
rect 35532 25372 35584 25424
rect 38016 25372 38068 25424
rect 41144 25372 41196 25424
rect 35440 25304 35492 25356
rect 39304 25304 39356 25356
rect 43996 25372 44048 25424
rect 33416 25236 33468 25245
rect 27068 25168 27120 25220
rect 31392 25211 31444 25220
rect 31392 25177 31401 25211
rect 31401 25177 31435 25211
rect 31435 25177 31444 25211
rect 31392 25168 31444 25177
rect 32680 25168 32732 25220
rect 34060 25211 34112 25220
rect 34060 25177 34087 25211
rect 34087 25177 34112 25211
rect 34060 25168 34112 25177
rect 34244 25211 34296 25220
rect 34244 25177 34253 25211
rect 34253 25177 34287 25211
rect 34287 25177 34296 25211
rect 34244 25168 34296 25177
rect 35256 25279 35308 25288
rect 35256 25245 35265 25279
rect 35265 25245 35299 25279
rect 35299 25245 35308 25279
rect 35256 25236 35308 25245
rect 35900 25279 35952 25288
rect 35900 25245 35909 25279
rect 35909 25245 35943 25279
rect 35943 25245 35952 25279
rect 35900 25236 35952 25245
rect 37280 25236 37332 25288
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 40224 25279 40276 25288
rect 40224 25245 40233 25279
rect 40233 25245 40267 25279
rect 40267 25245 40276 25279
rect 40224 25236 40276 25245
rect 40776 25236 40828 25288
rect 28356 25100 28408 25152
rect 35532 25100 35584 25152
rect 35716 25168 35768 25220
rect 38844 25211 38896 25220
rect 38844 25177 38853 25211
rect 38853 25177 38887 25211
rect 38887 25177 38896 25211
rect 38844 25168 38896 25177
rect 40132 25168 40184 25220
rect 43444 25304 43496 25356
rect 41236 25236 41288 25288
rect 41972 25236 42024 25288
rect 42432 25279 42484 25288
rect 42432 25245 42441 25279
rect 42441 25245 42475 25279
rect 42475 25245 42484 25279
rect 42432 25236 42484 25245
rect 43352 25279 43404 25288
rect 43352 25245 43361 25279
rect 43361 25245 43395 25279
rect 43395 25245 43404 25279
rect 43352 25236 43404 25245
rect 43904 25236 43956 25288
rect 46112 25236 46164 25288
rect 42984 25168 43036 25220
rect 43812 25168 43864 25220
rect 45468 25211 45520 25220
rect 45468 25177 45477 25211
rect 45477 25177 45511 25211
rect 45511 25177 45520 25211
rect 45468 25168 45520 25177
rect 37648 25143 37700 25152
rect 37648 25109 37657 25143
rect 37657 25109 37691 25143
rect 37691 25109 37700 25143
rect 37648 25100 37700 25109
rect 38108 25100 38160 25152
rect 39212 25100 39264 25152
rect 40316 25100 40368 25152
rect 40868 25143 40920 25152
rect 40868 25109 40877 25143
rect 40877 25109 40911 25143
rect 40911 25109 40920 25143
rect 40868 25100 40920 25109
rect 42156 25143 42208 25152
rect 42156 25109 42165 25143
rect 42165 25109 42199 25143
rect 42199 25109 42208 25143
rect 42156 25100 42208 25109
rect 43352 25100 43404 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 30472 24896 30524 24948
rect 34060 24896 34112 24948
rect 35256 24896 35308 24948
rect 35992 24896 36044 24948
rect 40500 24896 40552 24948
rect 41052 24939 41104 24948
rect 33968 24828 34020 24880
rect 24952 24760 25004 24812
rect 33324 24760 33376 24812
rect 37648 24828 37700 24880
rect 38752 24828 38804 24880
rect 40592 24828 40644 24880
rect 41052 24905 41061 24939
rect 41061 24905 41095 24939
rect 41095 24905 41104 24939
rect 41052 24896 41104 24905
rect 41696 24896 41748 24948
rect 42156 24896 42208 24948
rect 42984 24939 43036 24948
rect 42984 24905 43011 24939
rect 43011 24905 43036 24939
rect 42984 24896 43036 24905
rect 42432 24828 42484 24880
rect 43536 24828 43588 24880
rect 2044 24692 2096 24744
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 33876 24735 33928 24744
rect 33876 24701 33885 24735
rect 33885 24701 33919 24735
rect 33919 24701 33928 24735
rect 33876 24692 33928 24701
rect 34336 24803 34388 24812
rect 34336 24769 34345 24803
rect 34345 24769 34379 24803
rect 34379 24769 34388 24803
rect 34336 24760 34388 24769
rect 34520 24803 34572 24812
rect 34520 24769 34529 24803
rect 34529 24769 34563 24803
rect 34563 24769 34572 24803
rect 34520 24760 34572 24769
rect 34796 24760 34848 24812
rect 35348 24692 35400 24744
rect 35532 24735 35584 24744
rect 35532 24701 35541 24735
rect 35541 24701 35575 24735
rect 35575 24701 35584 24735
rect 35532 24692 35584 24701
rect 35900 24760 35952 24812
rect 36544 24760 36596 24812
rect 36820 24760 36872 24812
rect 37924 24803 37976 24812
rect 37924 24769 37933 24803
rect 37933 24769 37967 24803
rect 37967 24769 37976 24803
rect 37924 24760 37976 24769
rect 38016 24760 38068 24812
rect 38568 24803 38620 24812
rect 38568 24769 38577 24803
rect 38577 24769 38611 24803
rect 38611 24769 38620 24803
rect 38568 24760 38620 24769
rect 38844 24760 38896 24812
rect 39672 24760 39724 24812
rect 40960 24803 41012 24812
rect 35624 24667 35676 24676
rect 28448 24556 28500 24608
rect 33600 24556 33652 24608
rect 34244 24556 34296 24608
rect 35624 24633 35633 24667
rect 35633 24633 35667 24667
rect 35667 24633 35676 24667
rect 35624 24624 35676 24633
rect 36820 24667 36872 24676
rect 36820 24633 36829 24667
rect 36829 24633 36863 24667
rect 36863 24633 36872 24667
rect 36820 24624 36872 24633
rect 37280 24556 37332 24608
rect 38752 24692 38804 24744
rect 40960 24769 40969 24803
rect 40969 24769 41003 24803
rect 41003 24769 41012 24803
rect 40960 24760 41012 24769
rect 41604 24760 41656 24812
rect 43628 24760 43680 24812
rect 44272 24760 44324 24812
rect 44824 24803 44876 24812
rect 44824 24769 44833 24803
rect 44833 24769 44867 24803
rect 44867 24769 44876 24803
rect 44824 24760 44876 24769
rect 45468 24828 45520 24880
rect 45560 24760 45612 24812
rect 41236 24692 41288 24744
rect 41512 24692 41564 24744
rect 38568 24624 38620 24676
rect 42616 24624 42668 24676
rect 39212 24556 39264 24608
rect 40224 24556 40276 24608
rect 40684 24599 40736 24608
rect 40684 24565 40693 24599
rect 40693 24565 40727 24599
rect 40727 24565 40736 24599
rect 40684 24556 40736 24565
rect 43444 24624 43496 24676
rect 44088 24624 44140 24676
rect 45468 24667 45520 24676
rect 45468 24633 45477 24667
rect 45477 24633 45511 24667
rect 45511 24633 45520 24667
rect 45468 24624 45520 24633
rect 43812 24556 43864 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 34336 24352 34388 24404
rect 37832 24352 37884 24404
rect 37924 24352 37976 24404
rect 40132 24352 40184 24404
rect 40684 24395 40736 24404
rect 40684 24361 40693 24395
rect 40693 24361 40727 24395
rect 40727 24361 40736 24395
rect 40684 24352 40736 24361
rect 34520 24284 34572 24336
rect 29000 24216 29052 24268
rect 25964 24191 26016 24200
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 26424 24148 26476 24200
rect 27436 24123 27488 24132
rect 27436 24089 27445 24123
rect 27445 24089 27479 24123
rect 27479 24089 27488 24123
rect 27436 24080 27488 24089
rect 28264 24148 28316 24200
rect 29092 24148 29144 24200
rect 30748 24216 30800 24268
rect 33876 24216 33928 24268
rect 33968 24216 34020 24268
rect 38752 24284 38804 24336
rect 40040 24284 40092 24336
rect 42248 24352 42300 24404
rect 41144 24284 41196 24336
rect 43996 24352 44048 24404
rect 30104 24148 30156 24200
rect 31668 24148 31720 24200
rect 33416 24148 33468 24200
rect 33692 24148 33744 24200
rect 35440 24148 35492 24200
rect 35900 24148 35952 24200
rect 36544 24148 36596 24200
rect 36820 24148 36872 24200
rect 37280 24191 37332 24200
rect 28448 24080 28500 24132
rect 32588 24080 32640 24132
rect 27804 24012 27856 24064
rect 27988 24012 28040 24064
rect 32220 24012 32272 24064
rect 37280 24157 37289 24191
rect 37289 24157 37323 24191
rect 37323 24157 37332 24191
rect 37280 24148 37332 24157
rect 39304 24148 39356 24200
rect 40408 24148 40460 24200
rect 40868 24216 40920 24268
rect 40960 24216 41012 24268
rect 42616 24259 42668 24268
rect 41512 24191 41564 24200
rect 41512 24157 41521 24191
rect 41521 24157 41555 24191
rect 41555 24157 41564 24191
rect 41512 24148 41564 24157
rect 42616 24225 42625 24259
rect 42625 24225 42659 24259
rect 42659 24225 42668 24259
rect 42616 24216 42668 24225
rect 45468 24284 45520 24336
rect 44272 24216 44324 24268
rect 37188 24080 37240 24132
rect 38844 24123 38896 24132
rect 38844 24089 38853 24123
rect 38853 24089 38887 24123
rect 38887 24089 38896 24123
rect 38844 24080 38896 24089
rect 41696 24157 41705 24178
rect 41705 24157 41739 24178
rect 41739 24157 41748 24178
rect 41696 24126 41748 24157
rect 41972 24148 42024 24200
rect 42064 24148 42116 24200
rect 43536 24123 43588 24132
rect 43536 24089 43545 24123
rect 43545 24089 43579 24123
rect 43579 24089 43588 24123
rect 43536 24080 43588 24089
rect 43996 24148 44048 24200
rect 46112 24148 46164 24200
rect 44180 24080 44232 24132
rect 35348 24055 35400 24064
rect 35348 24021 35357 24055
rect 35357 24021 35391 24055
rect 35391 24021 35400 24055
rect 35348 24012 35400 24021
rect 35808 24012 35860 24064
rect 40132 24055 40184 24064
rect 40132 24021 40141 24055
rect 40141 24021 40175 24055
rect 40175 24021 40184 24055
rect 40132 24012 40184 24021
rect 40316 24055 40368 24064
rect 40316 24021 40325 24055
rect 40325 24021 40359 24055
rect 40359 24021 40368 24055
rect 40316 24012 40368 24021
rect 41236 24055 41288 24064
rect 41236 24021 41245 24055
rect 41245 24021 41279 24055
rect 41279 24021 41288 24055
rect 41236 24012 41288 24021
rect 41604 24012 41656 24064
rect 42616 24012 42668 24064
rect 45008 24012 45060 24064
rect 46020 24080 46072 24132
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 29092 23851 29144 23860
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 25044 23740 25096 23792
rect 25412 23740 25464 23792
rect 27896 23740 27948 23792
rect 28448 23783 28500 23792
rect 28448 23749 28457 23783
rect 28457 23749 28491 23783
rect 28491 23749 28500 23783
rect 28448 23740 28500 23749
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 2504 23468 2556 23520
rect 24952 23672 25004 23724
rect 25964 23672 26016 23724
rect 27988 23672 28040 23724
rect 28908 23672 28960 23724
rect 30288 23672 30340 23724
rect 34336 23808 34388 23860
rect 39304 23808 39356 23860
rect 41512 23808 41564 23860
rect 42432 23808 42484 23860
rect 43352 23851 43404 23860
rect 43352 23817 43361 23851
rect 43361 23817 43395 23851
rect 43395 23817 43404 23851
rect 43352 23808 43404 23817
rect 44548 23851 44600 23860
rect 44548 23817 44566 23851
rect 44566 23817 44600 23851
rect 44548 23808 44600 23817
rect 43536 23740 43588 23792
rect 43812 23740 43864 23792
rect 32956 23715 33008 23724
rect 32956 23681 32965 23715
rect 32965 23681 32999 23715
rect 32999 23681 33008 23715
rect 32956 23672 33008 23681
rect 33508 23672 33560 23724
rect 33692 23672 33744 23724
rect 25136 23647 25188 23656
rect 25136 23613 25145 23647
rect 25145 23613 25179 23647
rect 25179 23613 25188 23647
rect 25136 23604 25188 23613
rect 25596 23604 25648 23656
rect 26148 23536 26200 23588
rect 27252 23536 27304 23588
rect 28264 23604 28316 23656
rect 24860 23468 24912 23520
rect 25228 23468 25280 23520
rect 30748 23536 30800 23588
rect 31760 23604 31812 23656
rect 33600 23647 33652 23656
rect 33600 23613 33609 23647
rect 33609 23613 33643 23647
rect 33643 23613 33652 23647
rect 33600 23604 33652 23613
rect 35532 23672 35584 23724
rect 35808 23715 35860 23724
rect 35808 23681 35817 23715
rect 35817 23681 35851 23715
rect 35851 23681 35860 23715
rect 35808 23672 35860 23681
rect 36728 23672 36780 23724
rect 30564 23511 30616 23520
rect 30564 23477 30573 23511
rect 30573 23477 30607 23511
rect 30607 23477 30616 23511
rect 30564 23468 30616 23477
rect 35256 23604 35308 23656
rect 37372 23672 37424 23724
rect 38016 23672 38068 23724
rect 39488 23672 39540 23724
rect 39672 23715 39724 23724
rect 39672 23681 39681 23715
rect 39681 23681 39715 23715
rect 39715 23681 39724 23715
rect 39672 23672 39724 23681
rect 39764 23672 39816 23724
rect 41144 23715 41196 23724
rect 37004 23604 37056 23656
rect 37924 23647 37976 23656
rect 37924 23613 37933 23647
rect 37933 23613 37967 23647
rect 37967 23613 37976 23647
rect 37924 23604 37976 23613
rect 38568 23604 38620 23656
rect 39856 23604 39908 23656
rect 40684 23647 40736 23656
rect 40684 23613 40693 23647
rect 40693 23613 40727 23647
rect 40727 23613 40736 23647
rect 40684 23604 40736 23613
rect 41144 23681 41153 23715
rect 41153 23681 41187 23715
rect 41187 23681 41196 23715
rect 41144 23672 41196 23681
rect 43168 23715 43220 23724
rect 43168 23681 43177 23715
rect 43177 23681 43211 23715
rect 43211 23681 43220 23715
rect 43168 23672 43220 23681
rect 43444 23715 43496 23724
rect 43444 23681 43453 23715
rect 43453 23681 43487 23715
rect 43487 23681 43496 23715
rect 43444 23672 43496 23681
rect 43628 23672 43680 23724
rect 44180 23672 44232 23724
rect 46112 23672 46164 23724
rect 42064 23604 42116 23656
rect 42708 23604 42760 23656
rect 44916 23647 44968 23656
rect 39764 23536 39816 23588
rect 44916 23613 44925 23647
rect 44925 23613 44959 23647
rect 44959 23613 44968 23647
rect 44916 23604 44968 23613
rect 45560 23536 45612 23588
rect 33784 23511 33836 23520
rect 33784 23477 33793 23511
rect 33793 23477 33827 23511
rect 33827 23477 33836 23511
rect 33784 23468 33836 23477
rect 34428 23468 34480 23520
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 34704 23468 34756 23520
rect 35256 23468 35308 23520
rect 35992 23511 36044 23520
rect 35992 23477 36001 23511
rect 36001 23477 36035 23511
rect 36035 23477 36044 23511
rect 35992 23468 36044 23477
rect 36452 23468 36504 23520
rect 36544 23468 36596 23520
rect 36820 23468 36872 23520
rect 39212 23468 39264 23520
rect 40132 23468 40184 23520
rect 40868 23468 40920 23520
rect 41512 23468 41564 23520
rect 42984 23511 43036 23520
rect 42984 23477 42993 23511
rect 42993 23477 43027 23511
rect 43027 23477 43036 23511
rect 42984 23468 43036 23477
rect 43536 23468 43588 23520
rect 44916 23468 44968 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 24860 23264 24912 23316
rect 25412 23264 25464 23316
rect 33784 23264 33836 23316
rect 34244 23307 34296 23316
rect 34244 23273 34253 23307
rect 34253 23273 34287 23307
rect 34287 23273 34296 23307
rect 34244 23264 34296 23273
rect 35440 23264 35492 23316
rect 38660 23264 38712 23316
rect 38844 23264 38896 23316
rect 39488 23264 39540 23316
rect 45008 23264 45060 23316
rect 23848 23196 23900 23248
rect 26424 23171 26476 23180
rect 26424 23137 26433 23171
rect 26433 23137 26467 23171
rect 26467 23137 26476 23171
rect 26424 23128 26476 23137
rect 27160 23128 27212 23180
rect 27896 23171 27948 23180
rect 27896 23137 27905 23171
rect 27905 23137 27939 23171
rect 27939 23137 27948 23171
rect 27896 23128 27948 23137
rect 28908 23128 28960 23180
rect 22836 23060 22888 23112
rect 23572 23060 23624 23112
rect 25228 23060 25280 23112
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 22284 22992 22336 23044
rect 24584 22992 24636 23044
rect 26148 23060 26200 23112
rect 27804 23103 27856 23112
rect 27804 23069 27813 23103
rect 27813 23069 27847 23103
rect 27847 23069 27856 23103
rect 27804 23060 27856 23069
rect 29000 23060 29052 23112
rect 30288 23103 30340 23112
rect 30288 23069 30297 23103
rect 30297 23069 30331 23103
rect 30331 23069 30340 23103
rect 30288 23060 30340 23069
rect 30564 23128 30616 23180
rect 32404 23171 32456 23180
rect 32404 23137 32413 23171
rect 32413 23137 32447 23171
rect 32447 23137 32456 23171
rect 32404 23128 32456 23137
rect 31392 23060 31444 23112
rect 31760 23060 31812 23112
rect 33232 23103 33284 23112
rect 33232 23069 33241 23103
rect 33241 23069 33275 23103
rect 33275 23069 33284 23103
rect 33232 23060 33284 23069
rect 35256 23196 35308 23248
rect 35716 23196 35768 23248
rect 37188 23196 37240 23248
rect 39120 23196 39172 23248
rect 40592 23196 40644 23248
rect 43352 23196 43404 23248
rect 43536 23239 43588 23248
rect 43536 23205 43545 23239
rect 43545 23205 43579 23239
rect 43579 23205 43588 23239
rect 43536 23196 43588 23205
rect 34244 23128 34296 23180
rect 21732 22967 21784 22976
rect 21732 22933 21741 22967
rect 21741 22933 21775 22967
rect 21775 22933 21784 22967
rect 21732 22924 21784 22933
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 24768 22924 24820 22976
rect 25136 22924 25188 22976
rect 34612 23060 34664 23112
rect 35440 23128 35492 23180
rect 35348 23060 35400 23112
rect 35624 22992 35676 23044
rect 35716 23035 35768 23044
rect 35716 23001 35725 23035
rect 35725 23001 35759 23035
rect 35759 23001 35768 23035
rect 35716 22992 35768 23001
rect 36360 22992 36412 23044
rect 36728 23103 36780 23112
rect 36728 23069 36737 23103
rect 36737 23069 36771 23103
rect 36771 23069 36780 23103
rect 38476 23128 38528 23180
rect 36728 23060 36780 23069
rect 37280 23060 37332 23112
rect 36912 22992 36964 23044
rect 39304 23103 39356 23112
rect 39304 23069 39313 23103
rect 39313 23069 39347 23103
rect 39347 23069 39356 23103
rect 39304 23060 39356 23069
rect 39488 23060 39540 23112
rect 32772 22924 32824 22976
rect 33416 22924 33468 22976
rect 36084 22967 36136 22976
rect 36084 22933 36093 22967
rect 36093 22933 36127 22967
rect 36127 22933 36136 22967
rect 36084 22924 36136 22933
rect 37188 22924 37240 22976
rect 39948 23060 40000 23112
rect 40592 23060 40644 23112
rect 40868 23060 40920 23112
rect 41236 23103 41288 23112
rect 41236 23069 41245 23103
rect 41245 23069 41279 23103
rect 41279 23069 41288 23103
rect 41236 23060 41288 23069
rect 41420 23103 41472 23112
rect 41420 23069 41429 23103
rect 41429 23069 41463 23103
rect 41463 23069 41472 23103
rect 42984 23128 43036 23180
rect 41420 23060 41472 23069
rect 42708 23103 42760 23112
rect 38660 22924 38712 22976
rect 40040 22967 40092 22976
rect 40040 22933 40049 22967
rect 40049 22933 40083 22967
rect 40083 22933 40092 22967
rect 40040 22924 40092 22933
rect 41144 22992 41196 23044
rect 40960 22924 41012 22976
rect 41788 22992 41840 23044
rect 42708 23069 42717 23103
rect 42717 23069 42751 23103
rect 42751 23069 42760 23103
rect 42708 23060 42760 23069
rect 45560 23103 45612 23112
rect 45560 23069 45569 23103
rect 45569 23069 45603 23103
rect 45603 23069 45612 23103
rect 46112 23103 46164 23112
rect 45560 23060 45612 23069
rect 46112 23069 46121 23103
rect 46121 23069 46155 23103
rect 46155 23069 46164 23103
rect 46112 23060 46164 23069
rect 43812 23035 43864 23044
rect 43812 23001 43821 23035
rect 43821 23001 43855 23035
rect 43855 23001 43864 23035
rect 43812 22992 43864 23001
rect 44640 22992 44692 23044
rect 43168 22924 43220 22976
rect 43628 22924 43680 22976
rect 43996 22924 44048 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 22836 22763 22888 22772
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 24584 22763 24636 22772
rect 24584 22729 24593 22763
rect 24593 22729 24627 22763
rect 24627 22729 24636 22763
rect 24584 22720 24636 22729
rect 24952 22763 25004 22772
rect 24952 22729 24961 22763
rect 24961 22729 24995 22763
rect 24995 22729 25004 22763
rect 24952 22720 25004 22729
rect 27252 22763 27304 22772
rect 27252 22729 27261 22763
rect 27261 22729 27295 22763
rect 27295 22729 27304 22763
rect 27252 22720 27304 22729
rect 27896 22720 27948 22772
rect 32404 22763 32456 22772
rect 32404 22729 32413 22763
rect 32413 22729 32447 22763
rect 32447 22729 32456 22763
rect 32404 22720 32456 22729
rect 32772 22763 32824 22772
rect 32772 22729 32781 22763
rect 32781 22729 32815 22763
rect 32815 22729 32824 22763
rect 32772 22720 32824 22729
rect 26148 22652 26200 22704
rect 29000 22695 29052 22704
rect 29000 22661 29009 22695
rect 29009 22661 29043 22695
rect 29043 22661 29052 22695
rect 29000 22652 29052 22661
rect 32312 22652 32364 22704
rect 23572 22627 23624 22636
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 24768 22627 24820 22636
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25044 22584 25096 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 28172 22627 28224 22636
rect 25136 22559 25188 22568
rect 25136 22525 25145 22559
rect 25145 22525 25179 22559
rect 25179 22525 25188 22559
rect 25136 22516 25188 22525
rect 26976 22516 27028 22568
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 28172 22584 28224 22593
rect 29828 22559 29880 22568
rect 29828 22525 29837 22559
rect 29837 22525 29871 22559
rect 29871 22525 29880 22559
rect 29828 22516 29880 22525
rect 31852 22584 31904 22636
rect 32220 22584 32272 22636
rect 32588 22627 32640 22636
rect 32588 22593 32597 22627
rect 32597 22593 32631 22627
rect 32631 22593 32640 22627
rect 32588 22584 32640 22593
rect 34060 22720 34112 22772
rect 34244 22720 34296 22772
rect 34612 22720 34664 22772
rect 36268 22720 36320 22772
rect 39488 22763 39540 22772
rect 34428 22627 34480 22636
rect 29276 22448 29328 22500
rect 30840 22448 30892 22500
rect 31208 22380 31260 22432
rect 31392 22423 31444 22432
rect 31392 22389 31401 22423
rect 31401 22389 31435 22423
rect 31435 22389 31444 22423
rect 31392 22380 31444 22389
rect 33600 22380 33652 22432
rect 33876 22380 33928 22432
rect 34428 22593 34437 22627
rect 34437 22593 34471 22627
rect 34471 22593 34480 22627
rect 34428 22584 34480 22593
rect 34612 22584 34664 22636
rect 35256 22627 35308 22636
rect 35256 22593 35265 22627
rect 35265 22593 35299 22627
rect 35299 22593 35308 22627
rect 35256 22584 35308 22593
rect 34520 22448 34572 22500
rect 35716 22380 35768 22432
rect 35900 22627 35952 22636
rect 35900 22593 35909 22627
rect 35909 22593 35943 22627
rect 35943 22593 35952 22627
rect 37188 22652 37240 22704
rect 39488 22729 39497 22763
rect 39497 22729 39531 22763
rect 39531 22729 39540 22763
rect 39488 22720 39540 22729
rect 41144 22720 41196 22772
rect 39304 22652 39356 22704
rect 39764 22652 39816 22704
rect 39948 22652 40000 22704
rect 35900 22584 35952 22593
rect 36452 22584 36504 22636
rect 36636 22584 36688 22636
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 38660 22584 38712 22636
rect 39580 22584 39632 22636
rect 40868 22652 40920 22704
rect 41144 22627 41196 22636
rect 41144 22593 41153 22627
rect 41153 22593 41187 22627
rect 41187 22593 41196 22627
rect 41144 22584 41196 22593
rect 41788 22627 41840 22636
rect 35992 22559 36044 22568
rect 35992 22525 36001 22559
rect 36001 22525 36035 22559
rect 36035 22525 36044 22559
rect 35992 22516 36044 22525
rect 36176 22448 36228 22500
rect 37556 22516 37608 22568
rect 39028 22559 39080 22568
rect 39028 22525 39037 22559
rect 39037 22525 39071 22559
rect 39071 22525 39080 22559
rect 39028 22516 39080 22525
rect 39120 22559 39172 22568
rect 39120 22525 39129 22559
rect 39129 22525 39163 22559
rect 39163 22525 39172 22559
rect 39120 22516 39172 22525
rect 39948 22516 40000 22568
rect 40132 22559 40184 22568
rect 40132 22525 40141 22559
rect 40141 22525 40175 22559
rect 40175 22525 40184 22559
rect 40132 22516 40184 22525
rect 40224 22559 40276 22568
rect 40224 22525 40233 22559
rect 40233 22525 40267 22559
rect 40267 22525 40276 22559
rect 40224 22516 40276 22525
rect 39488 22448 39540 22500
rect 40592 22448 40644 22500
rect 41052 22448 41104 22500
rect 41788 22593 41797 22627
rect 41797 22593 41831 22627
rect 41831 22593 41840 22627
rect 41788 22584 41840 22593
rect 42984 22652 43036 22704
rect 43352 22652 43404 22704
rect 42340 22584 42392 22636
rect 41696 22448 41748 22500
rect 42616 22559 42668 22568
rect 42616 22525 42625 22559
rect 42625 22525 42659 22559
rect 42659 22525 42668 22559
rect 42616 22516 42668 22525
rect 42800 22516 42852 22568
rect 44640 22584 44692 22636
rect 45008 22627 45060 22636
rect 45008 22593 45017 22627
rect 45017 22593 45051 22627
rect 45051 22593 45060 22627
rect 45008 22584 45060 22593
rect 44088 22516 44140 22568
rect 45468 22516 45520 22568
rect 45744 22584 45796 22636
rect 45100 22448 45152 22500
rect 58256 22491 58308 22500
rect 58256 22457 58265 22491
rect 58265 22457 58299 22491
rect 58299 22457 58308 22491
rect 58256 22448 58308 22457
rect 38292 22380 38344 22432
rect 39120 22380 39172 22432
rect 43076 22423 43128 22432
rect 43076 22389 43085 22423
rect 43085 22389 43119 22423
rect 43119 22389 43128 22423
rect 43076 22380 43128 22389
rect 43996 22380 44048 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 24860 22176 24912 22228
rect 32588 22176 32640 22228
rect 33048 22176 33100 22228
rect 35992 22176 36044 22228
rect 25964 22108 26016 22160
rect 33416 22108 33468 22160
rect 34612 22108 34664 22160
rect 37740 22176 37792 22228
rect 38016 22176 38068 22228
rect 38614 22176 38666 22228
rect 39488 22176 39540 22228
rect 43168 22176 43220 22228
rect 36176 22108 36228 22160
rect 38384 22108 38436 22160
rect 22836 22040 22888 22092
rect 21732 21972 21784 22024
rect 1952 21904 2004 21956
rect 22284 21972 22336 22024
rect 23388 21947 23440 21956
rect 23388 21913 23397 21947
rect 23397 21913 23431 21947
rect 23431 21913 23440 21947
rect 23388 21904 23440 21913
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 25688 22040 25740 22092
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 29276 22040 29328 22092
rect 33232 22040 33284 22092
rect 25596 22015 25648 22024
rect 23756 21947 23808 21956
rect 23756 21913 23765 21947
rect 23765 21913 23799 21947
rect 23799 21913 23808 21947
rect 23756 21904 23808 21913
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 27160 21972 27212 22024
rect 30656 21972 30708 22024
rect 31024 21972 31076 22024
rect 31484 22015 31536 22024
rect 31484 21981 31493 22015
rect 31493 21981 31527 22015
rect 31527 21981 31536 22015
rect 31484 21972 31536 21981
rect 26516 21904 26568 21956
rect 30472 21836 30524 21888
rect 31852 21972 31904 22024
rect 33140 22015 33192 22024
rect 33140 21981 33149 22015
rect 33149 21981 33183 22015
rect 33183 21981 33192 22015
rect 33140 21972 33192 21981
rect 33324 21972 33376 22024
rect 35440 22040 35492 22092
rect 35716 22083 35768 22092
rect 35716 22049 35725 22083
rect 35725 22049 35759 22083
rect 35759 22049 35768 22083
rect 35716 22040 35768 22049
rect 34704 21972 34756 22024
rect 32588 21904 32640 21956
rect 34520 21904 34572 21956
rect 35072 21972 35124 22024
rect 36452 22040 36504 22092
rect 37004 22040 37056 22092
rect 41696 22108 41748 22160
rect 41788 22108 41840 22160
rect 45928 22108 45980 22160
rect 38660 22083 38712 22092
rect 38660 22049 38669 22083
rect 38669 22049 38703 22083
rect 38703 22049 38712 22083
rect 39304 22083 39356 22092
rect 38660 22040 38712 22049
rect 36820 21972 36872 22024
rect 38016 21972 38068 22024
rect 38200 21972 38252 22024
rect 39304 22049 39313 22083
rect 39313 22049 39347 22083
rect 39347 22049 39356 22083
rect 39304 22040 39356 22049
rect 39948 22040 40000 22092
rect 40960 22040 41012 22092
rect 36268 21904 36320 21956
rect 36728 21904 36780 21956
rect 37740 21947 37792 21956
rect 37740 21913 37749 21947
rect 37749 21913 37783 21947
rect 37783 21913 37792 21947
rect 37740 21904 37792 21913
rect 39764 21972 39816 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40040 21972 40092 21981
rect 40224 22015 40276 22024
rect 40224 21981 40233 22015
rect 40233 21981 40267 22015
rect 40267 21981 40276 22015
rect 40224 21972 40276 21981
rect 41144 21972 41196 22024
rect 41972 22040 42024 22092
rect 43628 22040 43680 22092
rect 33232 21836 33284 21888
rect 33876 21836 33928 21888
rect 35532 21836 35584 21888
rect 35808 21836 35860 21888
rect 36452 21836 36504 21888
rect 37372 21836 37424 21888
rect 40316 21904 40368 21956
rect 40960 21904 41012 21956
rect 39028 21836 39080 21888
rect 39856 21836 39908 21888
rect 40132 21836 40184 21888
rect 41236 21879 41288 21888
rect 41236 21845 41245 21879
rect 41245 21845 41279 21879
rect 41279 21845 41288 21879
rect 41236 21836 41288 21845
rect 42800 21972 42852 22024
rect 43352 22015 43404 22024
rect 43076 21904 43128 21956
rect 43352 21981 43361 22015
rect 43361 21981 43395 22015
rect 43395 21981 43404 22015
rect 43352 21972 43404 21981
rect 43996 21972 44048 22024
rect 43720 21904 43772 21956
rect 44272 21972 44324 22024
rect 45744 22040 45796 22092
rect 45376 22015 45428 22024
rect 45376 21981 45385 22015
rect 45385 21981 45419 22015
rect 45419 21981 45428 22015
rect 45376 21972 45428 21981
rect 45468 21972 45520 22024
rect 45836 22015 45888 22024
rect 45836 21981 45845 22015
rect 45845 21981 45879 22015
rect 45879 21981 45888 22015
rect 45836 21972 45888 21981
rect 44456 21904 44508 21956
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 23664 21675 23716 21684
rect 23664 21641 23673 21675
rect 23673 21641 23707 21675
rect 23707 21641 23716 21675
rect 23664 21632 23716 21641
rect 23756 21675 23808 21684
rect 23756 21641 23765 21675
rect 23765 21641 23799 21675
rect 23799 21641 23808 21675
rect 23756 21632 23808 21641
rect 25596 21632 25648 21684
rect 27896 21632 27948 21684
rect 28172 21632 28224 21684
rect 31024 21675 31076 21684
rect 31024 21641 31033 21675
rect 31033 21641 31067 21675
rect 31067 21641 31076 21675
rect 31024 21632 31076 21641
rect 33324 21632 33376 21684
rect 34060 21632 34112 21684
rect 34704 21632 34756 21684
rect 35440 21632 35492 21684
rect 36176 21632 36228 21684
rect 36820 21632 36872 21684
rect 37556 21632 37608 21684
rect 37832 21632 37884 21684
rect 38200 21632 38252 21684
rect 39304 21632 39356 21684
rect 44824 21675 44876 21684
rect 44824 21641 44833 21675
rect 44833 21641 44867 21675
rect 44867 21641 44876 21675
rect 44824 21632 44876 21641
rect 23296 21564 23348 21616
rect 23940 21564 23992 21616
rect 23480 21496 23532 21548
rect 23848 21496 23900 21548
rect 25688 21539 25740 21548
rect 25688 21505 25697 21539
rect 25697 21505 25731 21539
rect 25731 21505 25740 21539
rect 25688 21496 25740 21505
rect 28356 21496 28408 21548
rect 29828 21564 29880 21616
rect 32588 21607 32640 21616
rect 32588 21573 32597 21607
rect 32597 21573 32631 21607
rect 32631 21573 32640 21607
rect 32588 21564 32640 21573
rect 35072 21564 35124 21616
rect 36084 21564 36136 21616
rect 31208 21539 31260 21548
rect 31208 21505 31217 21539
rect 31217 21505 31251 21539
rect 31251 21505 31260 21539
rect 31208 21496 31260 21505
rect 22192 21428 22244 21480
rect 22836 21471 22888 21480
rect 22836 21437 22845 21471
rect 22845 21437 22879 21471
rect 22879 21437 22888 21471
rect 22836 21428 22888 21437
rect 23756 21428 23808 21480
rect 26056 21428 26108 21480
rect 29092 21471 29144 21480
rect 29092 21437 29101 21471
rect 29101 21437 29135 21471
rect 29135 21437 29144 21471
rect 29092 21428 29144 21437
rect 30472 21471 30524 21480
rect 25044 21360 25096 21412
rect 30472 21437 30481 21471
rect 30481 21437 30515 21471
rect 30515 21437 30524 21471
rect 30472 21428 30524 21437
rect 31484 21496 31536 21548
rect 32220 21496 32272 21548
rect 32404 21496 32456 21548
rect 33968 21539 34020 21548
rect 32772 21428 32824 21480
rect 33968 21505 33977 21539
rect 33977 21505 34011 21539
rect 34011 21505 34020 21539
rect 33968 21496 34020 21505
rect 34520 21496 34572 21548
rect 34704 21539 34756 21548
rect 34704 21505 34713 21539
rect 34713 21505 34747 21539
rect 34747 21505 34756 21539
rect 34704 21496 34756 21505
rect 35440 21496 35492 21548
rect 35624 21496 35676 21548
rect 35716 21539 35768 21548
rect 35716 21505 35725 21539
rect 35725 21505 35759 21539
rect 35759 21505 35768 21539
rect 36636 21564 36688 21616
rect 37004 21564 37056 21616
rect 35716 21496 35768 21505
rect 37188 21496 37240 21548
rect 37280 21428 37332 21480
rect 37648 21496 37700 21548
rect 38200 21539 38252 21548
rect 38200 21505 38209 21539
rect 38209 21505 38243 21539
rect 38243 21505 38252 21539
rect 38200 21496 38252 21505
rect 38568 21539 38620 21548
rect 38568 21505 38577 21539
rect 38577 21505 38611 21539
rect 38611 21505 38620 21539
rect 38568 21496 38620 21505
rect 38844 21496 38896 21548
rect 39764 21564 39816 21616
rect 39212 21496 39264 21548
rect 39856 21539 39908 21548
rect 37924 21428 37976 21480
rect 38476 21428 38528 21480
rect 39488 21428 39540 21480
rect 39856 21505 39865 21539
rect 39865 21505 39899 21539
rect 39899 21505 39908 21539
rect 39856 21496 39908 21505
rect 40408 21496 40460 21548
rect 41972 21564 42024 21616
rect 43536 21564 43588 21616
rect 44088 21564 44140 21616
rect 45836 21632 45888 21684
rect 45928 21675 45980 21684
rect 45928 21641 45937 21675
rect 45937 21641 45971 21675
rect 45971 21641 45980 21675
rect 45928 21632 45980 21641
rect 40868 21539 40920 21548
rect 40868 21505 40877 21539
rect 40877 21505 40911 21539
rect 40911 21505 40920 21539
rect 40868 21496 40920 21505
rect 41328 21496 41380 21548
rect 43260 21496 43312 21548
rect 43812 21496 43864 21548
rect 44180 21496 44232 21548
rect 44456 21496 44508 21548
rect 45468 21564 45520 21616
rect 45008 21539 45060 21548
rect 45008 21505 45017 21539
rect 45017 21505 45051 21539
rect 45051 21505 45060 21539
rect 45008 21496 45060 21505
rect 45284 21539 45336 21548
rect 45284 21505 45293 21539
rect 45293 21505 45327 21539
rect 45327 21505 45336 21539
rect 45284 21496 45336 21505
rect 40500 21428 40552 21480
rect 43720 21428 43772 21480
rect 44088 21428 44140 21480
rect 25964 21292 26016 21344
rect 27896 21292 27948 21344
rect 28908 21292 28960 21344
rect 31852 21360 31904 21412
rect 32312 21360 32364 21412
rect 35992 21360 36044 21412
rect 35716 21292 35768 21344
rect 35900 21292 35952 21344
rect 37188 21360 37240 21412
rect 39948 21360 40000 21412
rect 39396 21335 39448 21344
rect 39396 21301 39405 21335
rect 39405 21301 39439 21335
rect 39439 21301 39448 21335
rect 39396 21292 39448 21301
rect 39856 21292 39908 21344
rect 40132 21292 40184 21344
rect 40776 21292 40828 21344
rect 41052 21360 41104 21412
rect 41696 21403 41748 21412
rect 41696 21369 41705 21403
rect 41705 21369 41739 21403
rect 41739 21369 41748 21403
rect 41696 21360 41748 21369
rect 43260 21360 43312 21412
rect 43628 21360 43680 21412
rect 42708 21292 42760 21344
rect 42892 21292 42944 21344
rect 44640 21292 44692 21344
rect 46664 21335 46716 21344
rect 46664 21301 46673 21335
rect 46673 21301 46707 21335
rect 46707 21301 46716 21335
rect 46664 21292 46716 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 23388 21088 23440 21140
rect 25780 21131 25832 21140
rect 25780 21097 25789 21131
rect 25789 21097 25823 21131
rect 25823 21097 25832 21131
rect 25780 21088 25832 21097
rect 25688 20952 25740 21004
rect 31208 21088 31260 21140
rect 32404 21131 32456 21140
rect 32404 21097 32413 21131
rect 32413 21097 32447 21131
rect 32447 21097 32456 21131
rect 32404 21088 32456 21097
rect 32772 21088 32824 21140
rect 35624 21088 35676 21140
rect 36176 21088 36228 21140
rect 36728 21088 36780 21140
rect 36820 21088 36872 21140
rect 37648 21088 37700 21140
rect 37740 21088 37792 21140
rect 38384 21088 38436 21140
rect 27712 21020 27764 21072
rect 28356 21063 28408 21072
rect 28356 21029 28365 21063
rect 28365 21029 28399 21063
rect 28399 21029 28408 21063
rect 28356 21020 28408 21029
rect 23756 20884 23808 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 33232 20952 33284 21004
rect 23848 20884 23900 20893
rect 25596 20816 25648 20868
rect 25964 20884 26016 20936
rect 32220 20884 32272 20936
rect 26056 20859 26108 20868
rect 26056 20825 26065 20859
rect 26065 20825 26099 20859
rect 26099 20825 26108 20859
rect 26056 20816 26108 20825
rect 27896 20816 27948 20868
rect 30196 20816 30248 20868
rect 32956 20816 33008 20868
rect 33968 20884 34020 20936
rect 34888 20884 34940 20936
rect 35532 20884 35584 20936
rect 35992 20884 36044 20936
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25688 20748 25740 20800
rect 27528 20748 27580 20800
rect 29736 20791 29788 20800
rect 29736 20757 29745 20791
rect 29745 20757 29779 20791
rect 29779 20757 29788 20791
rect 29736 20748 29788 20757
rect 31852 20791 31904 20800
rect 31852 20757 31861 20791
rect 31861 20757 31895 20791
rect 31895 20757 31904 20791
rect 31852 20748 31904 20757
rect 32404 20748 32456 20800
rect 34060 20816 34112 20868
rect 35808 20816 35860 20868
rect 36084 20816 36136 20868
rect 36360 20952 36412 21004
rect 37188 20952 37240 21004
rect 37648 20952 37700 21004
rect 40592 21088 40644 21140
rect 41236 21088 41288 21140
rect 42708 21088 42760 21140
rect 39212 21020 39264 21072
rect 39856 21020 39908 21072
rect 40500 21020 40552 21072
rect 45100 21088 45152 21140
rect 39396 20952 39448 21004
rect 36452 20884 36504 20936
rect 36636 20927 36688 20936
rect 36636 20893 36645 20927
rect 36645 20893 36679 20927
rect 36679 20893 36688 20927
rect 36636 20884 36688 20893
rect 37280 20884 37332 20936
rect 37740 20884 37792 20936
rect 38844 20884 38896 20936
rect 39120 20927 39172 20936
rect 39120 20893 39129 20927
rect 39129 20893 39163 20927
rect 39163 20893 39172 20927
rect 41972 20952 42024 21004
rect 39120 20884 39172 20893
rect 37464 20859 37516 20868
rect 37464 20825 37473 20859
rect 37473 20825 37507 20859
rect 37507 20825 37516 20859
rect 37464 20816 37516 20825
rect 38568 20816 38620 20868
rect 39212 20816 39264 20868
rect 33600 20791 33652 20800
rect 33600 20757 33609 20791
rect 33609 20757 33643 20791
rect 33643 20757 33652 20791
rect 33600 20748 33652 20757
rect 35532 20791 35584 20800
rect 35532 20757 35541 20791
rect 35541 20757 35575 20791
rect 35575 20757 35584 20791
rect 35532 20748 35584 20757
rect 35992 20748 36044 20800
rect 36820 20791 36872 20800
rect 36820 20757 36829 20791
rect 36829 20757 36863 20791
rect 36863 20757 36872 20791
rect 36820 20748 36872 20757
rect 37280 20748 37332 20800
rect 37556 20748 37608 20800
rect 39120 20748 39172 20800
rect 40040 20816 40092 20868
rect 39948 20748 40000 20800
rect 42524 20884 42576 20936
rect 43536 20952 43588 21004
rect 43812 20884 43864 20936
rect 44180 20884 44232 20936
rect 45192 20884 45244 20936
rect 45652 20884 45704 20936
rect 40500 20791 40552 20800
rect 40500 20757 40509 20791
rect 40509 20757 40543 20791
rect 40543 20757 40552 20791
rect 40500 20748 40552 20757
rect 42156 20748 42208 20800
rect 42524 20748 42576 20800
rect 42800 20748 42852 20800
rect 44456 20816 44508 20868
rect 43720 20748 43772 20800
rect 43996 20748 44048 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 26976 20544 27028 20596
rect 35532 20544 35584 20596
rect 37556 20587 37608 20596
rect 37556 20553 37565 20587
rect 37565 20553 37599 20587
rect 37599 20553 37608 20587
rect 37556 20544 37608 20553
rect 38476 20544 38528 20596
rect 39028 20544 39080 20596
rect 39304 20544 39356 20596
rect 39488 20544 39540 20596
rect 23572 20476 23624 20528
rect 23020 20408 23072 20460
rect 25596 20408 25648 20460
rect 25688 20451 25740 20460
rect 25688 20417 25697 20451
rect 25697 20417 25731 20451
rect 25731 20417 25740 20451
rect 25688 20408 25740 20417
rect 27252 20408 27304 20460
rect 27896 20408 27948 20460
rect 29920 20408 29972 20460
rect 30196 20451 30248 20460
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30196 20408 30248 20417
rect 30380 20451 30432 20460
rect 30380 20417 30389 20451
rect 30389 20417 30423 20451
rect 30423 20417 30432 20451
rect 30380 20408 30432 20417
rect 22836 20383 22888 20392
rect 22836 20349 22845 20383
rect 22845 20349 22879 20383
rect 22879 20349 22888 20383
rect 22836 20340 22888 20349
rect 28724 20383 28776 20392
rect 28724 20349 28733 20383
rect 28733 20349 28767 20383
rect 28767 20349 28776 20383
rect 28724 20340 28776 20349
rect 29736 20340 29788 20392
rect 27528 20315 27580 20324
rect 27528 20281 27537 20315
rect 27537 20281 27571 20315
rect 27571 20281 27580 20315
rect 27528 20272 27580 20281
rect 29736 20247 29788 20256
rect 29736 20213 29745 20247
rect 29745 20213 29779 20247
rect 29779 20213 29788 20247
rect 29736 20204 29788 20213
rect 30288 20247 30340 20256
rect 30288 20213 30297 20247
rect 30297 20213 30331 20247
rect 30331 20213 30340 20247
rect 30288 20204 30340 20213
rect 32496 20476 32548 20528
rect 35992 20476 36044 20528
rect 36084 20476 36136 20528
rect 40684 20544 40736 20596
rect 41144 20544 41196 20596
rect 41788 20544 41840 20596
rect 41972 20544 42024 20596
rect 31852 20272 31904 20324
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33048 20408 33100 20460
rect 33876 20451 33928 20460
rect 33876 20417 33885 20451
rect 33885 20417 33919 20451
rect 33919 20417 33928 20451
rect 33876 20408 33928 20417
rect 34888 20408 34940 20460
rect 35900 20451 35952 20460
rect 35900 20417 35909 20451
rect 35909 20417 35943 20451
rect 35943 20417 35952 20451
rect 35900 20408 35952 20417
rect 36360 20451 36412 20460
rect 36360 20417 36369 20451
rect 36369 20417 36403 20451
rect 36403 20417 36412 20451
rect 36360 20408 36412 20417
rect 34796 20340 34848 20392
rect 35716 20340 35768 20392
rect 36636 20408 36688 20460
rect 37464 20451 37516 20460
rect 37464 20417 37473 20451
rect 37473 20417 37507 20451
rect 37507 20417 37516 20451
rect 37464 20408 37516 20417
rect 39304 20408 39356 20460
rect 39948 20408 40000 20460
rect 40224 20476 40276 20528
rect 40500 20476 40552 20528
rect 40868 20408 40920 20460
rect 41052 20408 41104 20460
rect 41880 20408 41932 20460
rect 42248 20408 42300 20460
rect 42432 20408 42484 20460
rect 43444 20544 43496 20596
rect 43812 20544 43864 20596
rect 42892 20451 42944 20460
rect 42892 20417 42901 20451
rect 42901 20417 42935 20451
rect 42935 20417 42944 20451
rect 42892 20408 42944 20417
rect 43352 20408 43404 20460
rect 43720 20408 43772 20460
rect 44180 20408 44232 20460
rect 45100 20476 45152 20528
rect 45192 20451 45244 20460
rect 45192 20417 45201 20451
rect 45201 20417 45235 20451
rect 45235 20417 45244 20451
rect 45192 20408 45244 20417
rect 45652 20451 45704 20460
rect 45652 20417 45661 20451
rect 45661 20417 45695 20451
rect 45695 20417 45704 20451
rect 45652 20408 45704 20417
rect 33416 20204 33468 20256
rect 33692 20247 33744 20256
rect 33692 20213 33701 20247
rect 33701 20213 33735 20247
rect 33735 20213 33744 20247
rect 33692 20204 33744 20213
rect 34060 20247 34112 20256
rect 34060 20213 34069 20247
rect 34069 20213 34103 20247
rect 34103 20213 34112 20247
rect 34060 20204 34112 20213
rect 34336 20272 34388 20324
rect 37740 20315 37792 20324
rect 37740 20281 37749 20315
rect 37749 20281 37783 20315
rect 37783 20281 37792 20315
rect 37740 20272 37792 20281
rect 41236 20340 41288 20392
rect 42064 20340 42116 20392
rect 40224 20272 40276 20324
rect 35440 20204 35492 20256
rect 36360 20204 36412 20256
rect 36636 20204 36688 20256
rect 39304 20204 39356 20256
rect 40132 20204 40184 20256
rect 41052 20272 41104 20324
rect 43628 20315 43680 20324
rect 43628 20281 43637 20315
rect 43637 20281 43671 20315
rect 43671 20281 43680 20315
rect 43628 20272 43680 20281
rect 44272 20272 44324 20324
rect 45928 20272 45980 20324
rect 40592 20204 40644 20256
rect 41144 20247 41196 20256
rect 41144 20213 41153 20247
rect 41153 20213 41187 20247
rect 41187 20213 41196 20247
rect 41144 20204 41196 20213
rect 41696 20204 41748 20256
rect 44364 20247 44416 20256
rect 44364 20213 44373 20247
rect 44373 20213 44407 20247
rect 44407 20213 44416 20247
rect 44364 20204 44416 20213
rect 44548 20247 44600 20256
rect 44548 20213 44557 20247
rect 44557 20213 44591 20247
rect 44591 20213 44600 20247
rect 44548 20204 44600 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 23664 20043 23716 20052
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 23756 20000 23808 20052
rect 26056 20000 26108 20052
rect 27252 20043 27304 20052
rect 27252 20009 27261 20043
rect 27261 20009 27295 20043
rect 27295 20009 27304 20043
rect 27252 20000 27304 20009
rect 25412 19932 25464 19984
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 28264 20000 28316 20052
rect 30748 20043 30800 20052
rect 30748 20009 30757 20043
rect 30757 20009 30791 20043
rect 30791 20009 30800 20043
rect 30748 20000 30800 20009
rect 32496 20000 32548 20052
rect 33140 20000 33192 20052
rect 34060 20000 34112 20052
rect 35624 20000 35676 20052
rect 35808 20000 35860 20052
rect 40776 20000 40828 20052
rect 32864 19932 32916 19984
rect 35900 19975 35952 19984
rect 35900 19941 35909 19975
rect 35909 19941 35943 19975
rect 35943 19941 35952 19975
rect 35900 19932 35952 19941
rect 35992 19932 36044 19984
rect 36452 19932 36504 19984
rect 37004 19932 37056 19984
rect 40684 19932 40736 19984
rect 27896 19864 27948 19916
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 23480 19796 23532 19848
rect 23756 19796 23808 19848
rect 24952 19796 25004 19848
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 29092 19864 29144 19916
rect 25320 19771 25372 19780
rect 25320 19737 25329 19771
rect 25329 19737 25363 19771
rect 25363 19737 25372 19771
rect 25320 19728 25372 19737
rect 27620 19728 27672 19780
rect 29736 19796 29788 19848
rect 30288 19839 30340 19848
rect 30288 19805 30292 19839
rect 30292 19805 30326 19839
rect 30326 19805 30340 19839
rect 30288 19796 30340 19805
rect 30564 19796 30616 19848
rect 35532 19864 35584 19916
rect 33048 19796 33100 19848
rect 33508 19839 33560 19848
rect 33508 19805 33517 19839
rect 33517 19805 33551 19839
rect 33551 19805 33560 19839
rect 33508 19796 33560 19805
rect 33784 19839 33836 19848
rect 33784 19805 33793 19839
rect 33793 19805 33827 19839
rect 33827 19805 33836 19839
rect 33784 19796 33836 19805
rect 34244 19796 34296 19848
rect 35348 19796 35400 19848
rect 35440 19796 35492 19848
rect 36084 19839 36136 19848
rect 36084 19805 36093 19839
rect 36093 19805 36127 19839
rect 36127 19805 36136 19839
rect 36084 19796 36136 19805
rect 33968 19728 34020 19780
rect 34060 19728 34112 19780
rect 35808 19728 35860 19780
rect 36360 19796 36412 19848
rect 37464 19839 37516 19848
rect 37464 19805 37473 19839
rect 37473 19805 37507 19839
rect 37507 19805 37516 19839
rect 37464 19796 37516 19805
rect 37832 19796 37884 19848
rect 38200 19796 38252 19848
rect 38476 19796 38528 19848
rect 39028 19771 39080 19780
rect 29736 19660 29788 19712
rect 30380 19660 30432 19712
rect 31852 19660 31904 19712
rect 33324 19660 33376 19712
rect 35440 19703 35492 19712
rect 35440 19669 35449 19703
rect 35449 19669 35483 19703
rect 35483 19669 35492 19703
rect 35440 19660 35492 19669
rect 35532 19660 35584 19712
rect 36452 19660 36504 19712
rect 37372 19703 37424 19712
rect 37372 19669 37381 19703
rect 37381 19669 37415 19703
rect 37415 19669 37424 19703
rect 37372 19660 37424 19669
rect 37464 19660 37516 19712
rect 39028 19737 39037 19771
rect 39037 19737 39071 19771
rect 39071 19737 39080 19771
rect 39028 19728 39080 19737
rect 39488 19796 39540 19848
rect 40040 19839 40092 19848
rect 40040 19805 40049 19839
rect 40049 19805 40083 19839
rect 40083 19805 40092 19839
rect 40040 19796 40092 19805
rect 40224 19839 40276 19848
rect 40224 19805 40233 19839
rect 40233 19805 40267 19839
rect 40267 19805 40276 19839
rect 40224 19796 40276 19805
rect 41144 19864 41196 19916
rect 40500 19839 40552 19848
rect 40500 19805 40509 19839
rect 40509 19805 40543 19839
rect 40543 19805 40552 19839
rect 40500 19796 40552 19805
rect 40592 19839 40644 19848
rect 40592 19805 40601 19839
rect 40601 19805 40635 19839
rect 40635 19805 40644 19839
rect 41972 20000 42024 20052
rect 44824 20000 44876 20052
rect 46020 20000 46072 20052
rect 41696 19975 41748 19984
rect 41696 19941 41705 19975
rect 41705 19941 41739 19975
rect 41739 19941 41748 19975
rect 41696 19932 41748 19941
rect 41880 19932 41932 19984
rect 42340 19932 42392 19984
rect 41512 19839 41564 19848
rect 40592 19796 40644 19805
rect 41512 19805 41521 19839
rect 41521 19805 41555 19839
rect 41555 19805 41564 19839
rect 41512 19796 41564 19805
rect 41788 19839 41840 19848
rect 41788 19805 41797 19839
rect 41797 19805 41831 19839
rect 41831 19805 41840 19839
rect 41788 19796 41840 19805
rect 41972 19839 42024 19848
rect 41972 19805 41981 19839
rect 41981 19805 42015 19839
rect 42015 19805 42024 19839
rect 41972 19796 42024 19805
rect 42616 19796 42668 19848
rect 44088 19864 44140 19916
rect 44272 19907 44324 19916
rect 44272 19873 44281 19907
rect 44281 19873 44315 19907
rect 44315 19873 44324 19907
rect 44272 19864 44324 19873
rect 44456 19907 44508 19916
rect 44456 19873 44465 19907
rect 44465 19873 44499 19907
rect 44499 19873 44508 19907
rect 44456 19864 44508 19873
rect 45192 19907 45244 19916
rect 45192 19873 45201 19907
rect 45201 19873 45235 19907
rect 45235 19873 45244 19907
rect 45192 19864 45244 19873
rect 42892 19728 42944 19780
rect 39488 19660 39540 19712
rect 41328 19703 41380 19712
rect 41328 19669 41337 19703
rect 41337 19669 41371 19703
rect 41371 19669 41380 19703
rect 41328 19660 41380 19669
rect 41696 19660 41748 19712
rect 43444 19796 43496 19848
rect 44180 19796 44232 19848
rect 46664 19864 46716 19916
rect 44088 19728 44140 19780
rect 45468 19839 45520 19848
rect 45468 19805 45477 19839
rect 45477 19805 45511 19839
rect 45511 19805 45520 19839
rect 45468 19796 45520 19805
rect 43352 19660 43404 19712
rect 45100 19728 45152 19780
rect 45468 19660 45520 19712
rect 45560 19660 45612 19712
rect 45928 19796 45980 19848
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 23848 19456 23900 19508
rect 26608 19456 26660 19508
rect 30196 19456 30248 19508
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 23664 19320 23716 19329
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 24216 19363 24268 19372
rect 23756 19320 23808 19329
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 24216 19320 24268 19329
rect 24400 19363 24452 19372
rect 24400 19329 24409 19363
rect 24409 19329 24443 19363
rect 24443 19329 24452 19363
rect 24400 19320 24452 19329
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 25688 19320 25740 19372
rect 27620 19388 27672 19440
rect 27896 19320 27948 19372
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 25412 19295 25464 19304
rect 25412 19261 25421 19295
rect 25421 19261 25455 19295
rect 25455 19261 25464 19295
rect 25412 19252 25464 19261
rect 28724 19252 28776 19304
rect 24308 19159 24360 19168
rect 24308 19125 24317 19159
rect 24317 19125 24351 19159
rect 24351 19125 24360 19159
rect 24308 19116 24360 19125
rect 25780 19116 25832 19168
rect 28448 19159 28500 19168
rect 28448 19125 28457 19159
rect 28457 19125 28491 19159
rect 28491 19125 28500 19159
rect 28448 19116 28500 19125
rect 29920 19320 29972 19372
rect 31852 19320 31904 19372
rect 37740 19456 37792 19508
rect 38108 19456 38160 19508
rect 38660 19456 38712 19508
rect 39764 19456 39816 19508
rect 40500 19499 40552 19508
rect 40500 19465 40509 19499
rect 40509 19465 40543 19499
rect 40543 19465 40552 19499
rect 40500 19456 40552 19465
rect 40684 19456 40736 19508
rect 43076 19456 43128 19508
rect 43260 19456 43312 19508
rect 46020 19499 46072 19508
rect 46020 19465 46029 19499
rect 46029 19465 46063 19499
rect 46063 19465 46072 19499
rect 46020 19456 46072 19465
rect 33232 19388 33284 19440
rect 33324 19320 33376 19372
rect 35992 19388 36044 19440
rect 36084 19388 36136 19440
rect 37372 19388 37424 19440
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 35348 19363 35400 19372
rect 34428 19320 34480 19329
rect 34520 19295 34572 19304
rect 34520 19261 34529 19295
rect 34529 19261 34563 19295
rect 34563 19261 34572 19295
rect 34520 19252 34572 19261
rect 34612 19329 34621 19338
rect 34621 19329 34655 19338
rect 34655 19329 34664 19338
rect 34612 19286 34664 19329
rect 35348 19329 35357 19363
rect 35357 19329 35391 19363
rect 35391 19329 35400 19363
rect 35348 19320 35400 19329
rect 35440 19363 35492 19372
rect 35440 19329 35449 19363
rect 35449 19329 35483 19363
rect 35483 19329 35492 19363
rect 35440 19320 35492 19329
rect 35808 19320 35860 19372
rect 36360 19363 36412 19372
rect 31392 19184 31444 19236
rect 32864 19227 32916 19236
rect 32864 19193 32873 19227
rect 32873 19193 32907 19227
rect 32907 19193 32916 19227
rect 32864 19184 32916 19193
rect 30564 19116 30616 19168
rect 33324 19116 33376 19168
rect 34336 19116 34388 19168
rect 35256 19116 35308 19168
rect 35992 19252 36044 19304
rect 36360 19329 36369 19363
rect 36369 19329 36403 19363
rect 36403 19329 36412 19363
rect 36360 19320 36412 19329
rect 36636 19320 36688 19372
rect 37740 19363 37792 19372
rect 37740 19329 37749 19363
rect 37749 19329 37783 19363
rect 37783 19329 37792 19363
rect 37740 19320 37792 19329
rect 37372 19252 37424 19304
rect 37924 19363 37976 19372
rect 37924 19329 37933 19363
rect 37933 19329 37967 19363
rect 37967 19329 37976 19363
rect 40224 19388 40276 19440
rect 37924 19320 37976 19329
rect 38936 19320 38988 19372
rect 38200 19252 38252 19304
rect 39304 19363 39356 19372
rect 39304 19329 39313 19363
rect 39313 19329 39347 19363
rect 39347 19329 39356 19363
rect 39304 19320 39356 19329
rect 39488 19363 39540 19372
rect 39488 19329 39497 19363
rect 39497 19329 39531 19363
rect 39531 19329 39540 19363
rect 39488 19320 39540 19329
rect 40316 19320 40368 19372
rect 42064 19431 42116 19440
rect 42064 19397 42073 19431
rect 42073 19397 42107 19431
rect 42107 19397 42116 19431
rect 42064 19388 42116 19397
rect 40868 19320 40920 19372
rect 41880 19320 41932 19372
rect 42432 19320 42484 19372
rect 42708 19320 42760 19372
rect 43168 19388 43220 19440
rect 43352 19388 43404 19440
rect 43444 19388 43496 19440
rect 43260 19363 43312 19372
rect 43260 19329 43269 19363
rect 43269 19329 43303 19363
rect 43303 19329 43312 19363
rect 43260 19320 43312 19329
rect 43904 19363 43956 19372
rect 43904 19329 43913 19363
rect 43913 19329 43947 19363
rect 43947 19329 43956 19363
rect 43904 19320 43956 19329
rect 41420 19252 41472 19304
rect 41512 19295 41564 19304
rect 41512 19261 41521 19295
rect 41521 19261 41555 19295
rect 41555 19261 41564 19295
rect 41512 19252 41564 19261
rect 41788 19252 41840 19304
rect 36636 19184 36688 19236
rect 36452 19116 36504 19168
rect 37556 19116 37608 19168
rect 37924 19116 37976 19168
rect 38384 19116 38436 19168
rect 38844 19159 38896 19168
rect 38844 19125 38853 19159
rect 38853 19125 38887 19159
rect 38887 19125 38896 19159
rect 38844 19116 38896 19125
rect 41052 19184 41104 19236
rect 45836 19320 45888 19372
rect 44272 19184 44324 19236
rect 45376 19252 45428 19304
rect 41788 19116 41840 19168
rect 43076 19159 43128 19168
rect 43076 19125 43085 19159
rect 43085 19125 43119 19159
rect 43119 19125 43128 19159
rect 43076 19116 43128 19125
rect 44088 19116 44140 19168
rect 44916 19116 44968 19168
rect 45284 19159 45336 19168
rect 45284 19125 45293 19159
rect 45293 19125 45327 19159
rect 45327 19125 45336 19159
rect 45284 19116 45336 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 23480 18912 23532 18964
rect 25964 18955 26016 18964
rect 25964 18921 25973 18955
rect 25973 18921 26007 18955
rect 26007 18921 26016 18955
rect 25964 18912 26016 18921
rect 27620 18955 27672 18964
rect 27620 18921 27629 18955
rect 27629 18921 27663 18955
rect 27663 18921 27672 18955
rect 27620 18912 27672 18921
rect 27804 18887 27856 18896
rect 27804 18853 27813 18887
rect 27813 18853 27847 18887
rect 27847 18853 27856 18887
rect 27804 18844 27856 18853
rect 33048 18912 33100 18964
rect 36084 18912 36136 18964
rect 35532 18844 35584 18896
rect 39028 18912 39080 18964
rect 39304 18912 39356 18964
rect 36360 18844 36412 18896
rect 36636 18844 36688 18896
rect 37464 18887 37516 18896
rect 37464 18853 37473 18887
rect 37473 18853 37507 18887
rect 37507 18853 37516 18887
rect 37464 18844 37516 18853
rect 38200 18844 38252 18896
rect 38936 18844 38988 18896
rect 41144 18844 41196 18896
rect 41512 18912 41564 18964
rect 42432 18912 42484 18964
rect 44180 18912 44232 18964
rect 46112 18912 46164 18964
rect 43444 18887 43496 18896
rect 23572 18776 23624 18828
rect 28448 18776 28500 18828
rect 31760 18776 31812 18828
rect 24308 18708 24360 18760
rect 24584 18708 24636 18760
rect 25044 18708 25096 18760
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 25964 18751 26016 18760
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 25964 18708 26016 18717
rect 31024 18751 31076 18760
rect 31024 18717 31033 18751
rect 31033 18717 31067 18751
rect 31067 18717 31076 18751
rect 31024 18708 31076 18717
rect 31392 18751 31444 18760
rect 28080 18683 28132 18692
rect 28080 18649 28089 18683
rect 28089 18649 28123 18683
rect 28123 18649 28132 18683
rect 28080 18640 28132 18649
rect 31392 18717 31401 18751
rect 31401 18717 31435 18751
rect 31435 18717 31444 18751
rect 31392 18708 31444 18717
rect 32220 18751 32272 18760
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 33048 18751 33100 18760
rect 33048 18717 33057 18751
rect 33057 18717 33091 18751
rect 33091 18717 33100 18751
rect 33048 18708 33100 18717
rect 33600 18708 33652 18760
rect 37924 18776 37976 18828
rect 38844 18776 38896 18828
rect 39488 18776 39540 18828
rect 41880 18819 41932 18828
rect 41880 18785 41889 18819
rect 41889 18785 41923 18819
rect 41923 18785 41932 18819
rect 41880 18776 41932 18785
rect 34336 18751 34388 18760
rect 34336 18717 34345 18751
rect 34345 18717 34379 18751
rect 34379 18717 34388 18751
rect 34336 18708 34388 18717
rect 34612 18708 34664 18760
rect 35532 18751 35584 18760
rect 35532 18717 35541 18751
rect 35541 18717 35575 18751
rect 35575 18717 35584 18751
rect 35532 18708 35584 18717
rect 37381 18745 37433 18757
rect 37381 18711 37390 18745
rect 37390 18711 37424 18745
rect 37424 18711 37433 18745
rect 37648 18751 37700 18760
rect 37381 18705 37433 18711
rect 37648 18717 37657 18751
rect 37657 18717 37691 18751
rect 37691 18717 37700 18751
rect 37648 18708 37700 18717
rect 37740 18708 37792 18760
rect 40776 18751 40828 18760
rect 32036 18683 32088 18692
rect 32036 18649 32045 18683
rect 32045 18649 32079 18683
rect 32079 18649 32088 18683
rect 32036 18640 32088 18649
rect 33324 18640 33376 18692
rect 23848 18572 23900 18624
rect 24216 18572 24268 18624
rect 25596 18572 25648 18624
rect 31116 18572 31168 18624
rect 32680 18572 32732 18624
rect 35348 18572 35400 18624
rect 36452 18640 36504 18692
rect 36636 18640 36688 18692
rect 38384 18640 38436 18692
rect 39212 18640 39264 18692
rect 38200 18572 38252 18624
rect 38568 18572 38620 18624
rect 39028 18572 39080 18624
rect 40500 18640 40552 18692
rect 40776 18717 40788 18751
rect 40788 18717 40828 18751
rect 40776 18708 40828 18717
rect 41052 18708 41104 18760
rect 43444 18853 43453 18887
rect 43453 18853 43487 18887
rect 43487 18853 43496 18887
rect 43444 18844 43496 18853
rect 44272 18844 44324 18896
rect 42800 18776 42852 18828
rect 43720 18776 43772 18828
rect 42524 18683 42576 18692
rect 42524 18649 42533 18683
rect 42533 18649 42567 18683
rect 42567 18649 42576 18683
rect 42524 18640 42576 18649
rect 43628 18751 43680 18760
rect 43628 18717 43637 18751
rect 43637 18717 43671 18751
rect 43671 18717 43680 18751
rect 43628 18708 43680 18717
rect 43812 18751 43864 18760
rect 43812 18717 43821 18751
rect 43821 18717 43855 18751
rect 43855 18717 43864 18751
rect 43812 18708 43864 18717
rect 44916 18708 44968 18760
rect 45836 18708 45888 18760
rect 41512 18572 41564 18624
rect 43536 18572 43588 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 32128 18368 32180 18420
rect 33232 18411 33284 18420
rect 33232 18377 33241 18411
rect 33241 18377 33275 18411
rect 33275 18377 33284 18411
rect 33232 18368 33284 18377
rect 34704 18368 34756 18420
rect 30564 18343 30616 18352
rect 30564 18309 30573 18343
rect 30573 18309 30607 18343
rect 30607 18309 30616 18343
rect 30564 18300 30616 18309
rect 31116 18343 31168 18352
rect 31116 18309 31125 18343
rect 31125 18309 31159 18343
rect 31159 18309 31168 18343
rect 31116 18300 31168 18309
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 24400 18232 24452 18284
rect 25780 18232 25832 18284
rect 27528 18275 27580 18284
rect 27528 18241 27537 18275
rect 27537 18241 27571 18275
rect 27571 18241 27580 18275
rect 27528 18232 27580 18241
rect 29920 18232 29972 18284
rect 32036 18232 32088 18284
rect 32496 18232 32548 18284
rect 34060 18300 34112 18352
rect 24308 18139 24360 18148
rect 24308 18105 24317 18139
rect 24317 18105 24351 18139
rect 24351 18105 24360 18139
rect 24308 18096 24360 18105
rect 27804 18164 27856 18216
rect 28724 18207 28776 18216
rect 28724 18173 28733 18207
rect 28733 18173 28767 18207
rect 28767 18173 28776 18207
rect 28724 18164 28776 18173
rect 32220 18164 32272 18216
rect 25964 18096 26016 18148
rect 25504 18028 25556 18080
rect 27252 18071 27304 18080
rect 27252 18037 27261 18071
rect 27261 18037 27295 18071
rect 27295 18037 27304 18071
rect 27252 18028 27304 18037
rect 30012 18028 30064 18080
rect 30196 18071 30248 18080
rect 30196 18037 30205 18071
rect 30205 18037 30239 18071
rect 30239 18037 30248 18071
rect 30196 18028 30248 18037
rect 31944 18096 31996 18148
rect 32956 18096 33008 18148
rect 33324 18232 33376 18284
rect 34428 18232 34480 18284
rect 31392 18028 31444 18080
rect 32588 18071 32640 18080
rect 32588 18037 32597 18071
rect 32597 18037 32631 18071
rect 32631 18037 32640 18071
rect 32588 18028 32640 18037
rect 33876 18071 33928 18080
rect 33876 18037 33885 18071
rect 33885 18037 33919 18071
rect 33919 18037 33928 18071
rect 33876 18028 33928 18037
rect 35440 18232 35492 18284
rect 35808 18232 35860 18284
rect 37832 18368 37884 18420
rect 36912 18300 36964 18352
rect 36176 18275 36228 18284
rect 36176 18241 36185 18275
rect 36185 18241 36219 18275
rect 36219 18241 36228 18275
rect 36176 18232 36228 18241
rect 36544 18232 36596 18284
rect 37372 18232 37424 18284
rect 37832 18232 37884 18284
rect 38384 18368 38436 18420
rect 39304 18368 39356 18420
rect 39764 18411 39816 18420
rect 39764 18377 39773 18411
rect 39773 18377 39807 18411
rect 39807 18377 39816 18411
rect 39764 18368 39816 18377
rect 40408 18368 40460 18420
rect 40592 18368 40644 18420
rect 42800 18411 42852 18420
rect 42800 18377 42809 18411
rect 42809 18377 42843 18411
rect 42843 18377 42852 18411
rect 42800 18368 42852 18377
rect 43536 18368 43588 18420
rect 42984 18300 43036 18352
rect 43444 18300 43496 18352
rect 38384 18232 38436 18284
rect 38660 18232 38712 18284
rect 39488 18275 39540 18284
rect 39488 18241 39497 18275
rect 39497 18241 39531 18275
rect 39531 18241 39540 18275
rect 39488 18232 39540 18241
rect 39580 18232 39632 18284
rect 41328 18232 41380 18284
rect 42892 18232 42944 18284
rect 43260 18232 43312 18284
rect 43812 18275 43864 18284
rect 43812 18241 43821 18275
rect 43821 18241 43855 18275
rect 43855 18241 43864 18275
rect 43812 18232 43864 18241
rect 44272 18232 44324 18284
rect 44916 18232 44968 18284
rect 37740 18164 37792 18216
rect 38844 18164 38896 18216
rect 40316 18164 40368 18216
rect 41512 18164 41564 18216
rect 42524 18164 42576 18216
rect 44548 18164 44600 18216
rect 45192 18164 45244 18216
rect 35624 18096 35676 18148
rect 38660 18139 38712 18148
rect 38660 18105 38669 18139
rect 38669 18105 38703 18139
rect 38703 18105 38712 18139
rect 38660 18096 38712 18105
rect 46480 18096 46532 18148
rect 35440 18028 35492 18080
rect 35900 18028 35952 18080
rect 36452 18028 36504 18080
rect 38200 18028 38252 18080
rect 38476 18028 38528 18080
rect 38936 18071 38988 18080
rect 38936 18037 38945 18071
rect 38945 18037 38979 18071
rect 38979 18037 38988 18071
rect 38936 18028 38988 18037
rect 39028 18028 39080 18080
rect 43168 18028 43220 18080
rect 45744 18028 45796 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 24400 17824 24452 17876
rect 27528 17824 27580 17876
rect 29736 17867 29788 17876
rect 29736 17833 29745 17867
rect 29745 17833 29779 17867
rect 29779 17833 29788 17867
rect 29736 17824 29788 17833
rect 32956 17867 33008 17876
rect 32956 17833 32965 17867
rect 32965 17833 32999 17867
rect 32999 17833 33008 17867
rect 32956 17824 33008 17833
rect 33416 17867 33468 17876
rect 33416 17833 33425 17867
rect 33425 17833 33459 17867
rect 33459 17833 33468 17867
rect 33416 17824 33468 17833
rect 36176 17824 36228 17876
rect 37372 17824 37424 17876
rect 38200 17867 38252 17876
rect 38200 17833 38209 17867
rect 38209 17833 38243 17867
rect 38243 17833 38252 17867
rect 38200 17824 38252 17833
rect 38384 17824 38436 17876
rect 40684 17824 40736 17876
rect 41512 17867 41564 17876
rect 41512 17833 41521 17867
rect 41521 17833 41555 17867
rect 41555 17833 41564 17867
rect 41512 17824 41564 17833
rect 42064 17824 42116 17876
rect 42524 17824 42576 17876
rect 43444 17824 43496 17876
rect 25412 17756 25464 17808
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 25044 17620 25096 17672
rect 25504 17620 25556 17672
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 25964 17663 26016 17672
rect 25964 17629 25973 17663
rect 25973 17629 26007 17663
rect 26007 17629 26016 17663
rect 28080 17756 28132 17808
rect 25964 17620 26016 17629
rect 26516 17620 26568 17672
rect 27804 17552 27856 17604
rect 26056 17484 26108 17536
rect 30196 17756 30248 17808
rect 36820 17756 36872 17808
rect 29920 17663 29972 17672
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 29920 17620 29972 17629
rect 31392 17663 31444 17672
rect 28724 17552 28776 17604
rect 29460 17552 29512 17604
rect 31392 17629 31401 17663
rect 31401 17629 31435 17663
rect 31435 17629 31444 17663
rect 31392 17620 31444 17629
rect 31944 17688 31996 17740
rect 34704 17688 34756 17740
rect 35440 17731 35492 17740
rect 35440 17697 35449 17731
rect 35449 17697 35483 17731
rect 35483 17697 35492 17731
rect 35440 17688 35492 17697
rect 31852 17595 31904 17604
rect 31852 17561 31861 17595
rect 31861 17561 31895 17595
rect 31895 17561 31904 17595
rect 31852 17552 31904 17561
rect 32128 17663 32180 17672
rect 32128 17629 32137 17663
rect 32137 17629 32171 17663
rect 32171 17629 32180 17663
rect 32128 17620 32180 17629
rect 33416 17620 33468 17672
rect 34428 17620 34480 17672
rect 36268 17688 36320 17740
rect 36728 17620 36780 17672
rect 37556 17688 37608 17740
rect 37740 17688 37792 17740
rect 38108 17688 38160 17740
rect 40500 17688 40552 17740
rect 41696 17756 41748 17808
rect 38844 17663 38896 17672
rect 37188 17595 37240 17604
rect 28448 17484 28500 17536
rect 31116 17484 31168 17536
rect 31392 17484 31444 17536
rect 33784 17527 33836 17536
rect 33784 17493 33793 17527
rect 33793 17493 33827 17527
rect 33827 17493 33836 17527
rect 33784 17484 33836 17493
rect 34060 17484 34112 17536
rect 35900 17527 35952 17536
rect 35900 17493 35909 17527
rect 35909 17493 35943 17527
rect 35943 17493 35952 17527
rect 35900 17484 35952 17493
rect 36084 17527 36136 17536
rect 36084 17493 36093 17527
rect 36093 17493 36127 17527
rect 36127 17493 36136 17527
rect 36084 17484 36136 17493
rect 37188 17561 37197 17595
rect 37197 17561 37231 17595
rect 37231 17561 37240 17595
rect 37188 17552 37240 17561
rect 37648 17552 37700 17604
rect 38844 17629 38853 17663
rect 38853 17629 38887 17663
rect 38887 17629 38896 17663
rect 38844 17620 38896 17629
rect 39120 17663 39172 17672
rect 39120 17629 39129 17663
rect 39129 17629 39163 17663
rect 39163 17629 39172 17663
rect 39120 17620 39172 17629
rect 39948 17620 40000 17672
rect 40132 17663 40184 17672
rect 40132 17629 40141 17663
rect 40141 17629 40175 17663
rect 40175 17629 40184 17663
rect 40132 17620 40184 17629
rect 41420 17688 41472 17740
rect 41512 17688 41564 17740
rect 42800 17756 42852 17808
rect 42892 17756 42944 17808
rect 41236 17663 41288 17672
rect 38476 17552 38528 17604
rect 40224 17552 40276 17604
rect 39212 17484 39264 17536
rect 40316 17527 40368 17536
rect 40316 17493 40325 17527
rect 40325 17493 40359 17527
rect 40359 17493 40368 17527
rect 40316 17484 40368 17493
rect 41236 17629 41245 17663
rect 41245 17629 41279 17663
rect 41279 17629 41288 17663
rect 41236 17620 41288 17629
rect 42432 17620 42484 17672
rect 42708 17663 42760 17672
rect 42708 17629 42717 17663
rect 42717 17629 42751 17663
rect 42751 17629 42760 17663
rect 42708 17620 42760 17629
rect 43168 17620 43220 17672
rect 44916 17688 44968 17740
rect 45100 17620 45152 17672
rect 45468 17620 45520 17672
rect 45836 17663 45888 17672
rect 45836 17629 45845 17663
rect 45845 17629 45879 17663
rect 45879 17629 45888 17663
rect 45836 17620 45888 17629
rect 41972 17484 42024 17536
rect 42524 17595 42576 17604
rect 42524 17561 42533 17595
rect 42533 17561 42567 17595
rect 42567 17561 42576 17595
rect 42524 17552 42576 17561
rect 42616 17595 42668 17604
rect 42616 17561 42625 17595
rect 42625 17561 42659 17595
rect 42659 17561 42668 17595
rect 43536 17595 43588 17604
rect 42616 17552 42668 17561
rect 43536 17561 43563 17595
rect 43563 17561 43588 17595
rect 43536 17552 43588 17561
rect 43996 17552 44048 17604
rect 44180 17595 44232 17604
rect 44180 17561 44189 17595
rect 44189 17561 44223 17595
rect 44223 17561 44232 17595
rect 44180 17552 44232 17561
rect 42800 17484 42852 17536
rect 43260 17484 43312 17536
rect 44548 17484 44600 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 31944 17280 31996 17332
rect 33416 17323 33468 17332
rect 33416 17289 33425 17323
rect 33425 17289 33459 17323
rect 33459 17289 33468 17323
rect 33416 17280 33468 17289
rect 34060 17323 34112 17332
rect 34060 17289 34069 17323
rect 34069 17289 34103 17323
rect 34103 17289 34112 17323
rect 34060 17280 34112 17289
rect 34244 17280 34296 17332
rect 2504 17212 2556 17264
rect 31392 17212 31444 17264
rect 33232 17255 33284 17264
rect 16856 17144 16908 17196
rect 23664 17187 23716 17196
rect 23664 17153 23673 17187
rect 23673 17153 23707 17187
rect 23707 17153 23716 17187
rect 23664 17144 23716 17153
rect 23940 17144 23992 17196
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 25044 17144 25096 17196
rect 26056 17187 26108 17196
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 30104 17187 30156 17196
rect 30104 17153 30113 17187
rect 30113 17153 30147 17187
rect 30147 17153 30156 17187
rect 30104 17144 30156 17153
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 33232 17221 33241 17255
rect 33241 17221 33275 17255
rect 33275 17221 33284 17255
rect 33232 17212 33284 17221
rect 32588 17187 32640 17196
rect 32588 17153 32597 17187
rect 32597 17153 32631 17187
rect 32631 17153 32640 17187
rect 32588 17144 32640 17153
rect 32956 17144 33008 17196
rect 35348 17212 35400 17264
rect 33968 17076 34020 17128
rect 34336 17187 34388 17196
rect 34336 17153 34345 17187
rect 34345 17153 34379 17187
rect 34379 17153 34388 17187
rect 34336 17144 34388 17153
rect 34520 17144 34572 17196
rect 36544 17280 36596 17332
rect 36820 17280 36872 17332
rect 37556 17280 37608 17332
rect 37924 17280 37976 17332
rect 38108 17280 38160 17332
rect 39396 17280 39448 17332
rect 39488 17280 39540 17332
rect 40776 17323 40828 17332
rect 40776 17289 40785 17323
rect 40785 17289 40819 17323
rect 40819 17289 40828 17323
rect 40776 17280 40828 17289
rect 41512 17280 41564 17332
rect 42064 17323 42116 17332
rect 42064 17289 42073 17323
rect 42073 17289 42107 17323
rect 42107 17289 42116 17323
rect 42064 17280 42116 17289
rect 1676 17051 1728 17060
rect 1676 17017 1685 17051
rect 1685 17017 1719 17051
rect 1719 17017 1728 17051
rect 1676 17008 1728 17017
rect 27252 17051 27304 17060
rect 27252 17017 27261 17051
rect 27261 17017 27295 17051
rect 27295 17017 27304 17051
rect 27252 17008 27304 17017
rect 39028 17212 39080 17264
rect 36636 17144 36688 17196
rect 37556 17144 37608 17196
rect 37740 17187 37792 17196
rect 37740 17153 37749 17187
rect 37749 17153 37783 17187
rect 37783 17153 37792 17187
rect 37740 17144 37792 17153
rect 38384 17076 38436 17128
rect 38660 17144 38712 17196
rect 39304 17144 39356 17196
rect 40500 17212 40552 17264
rect 39580 17144 39632 17196
rect 40684 17187 40736 17196
rect 40684 17153 40693 17187
rect 40693 17153 40727 17187
rect 40727 17153 40736 17187
rect 40684 17144 40736 17153
rect 40960 17187 41012 17196
rect 40960 17153 40969 17187
rect 40969 17153 41003 17187
rect 41003 17153 41012 17187
rect 40960 17144 41012 17153
rect 41328 17144 41380 17196
rect 42616 17187 42668 17196
rect 42616 17153 42625 17187
rect 42625 17153 42659 17187
rect 42659 17153 42668 17187
rect 42616 17144 42668 17153
rect 42800 17187 42852 17196
rect 42800 17153 42809 17187
rect 42809 17153 42843 17187
rect 42843 17153 42852 17187
rect 42800 17144 42852 17153
rect 42892 17187 42944 17196
rect 42892 17153 42901 17187
rect 42901 17153 42935 17187
rect 42935 17153 42944 17187
rect 42892 17144 42944 17153
rect 43076 17144 43128 17196
rect 43536 17144 43588 17196
rect 45008 17212 45060 17264
rect 44916 17187 44968 17196
rect 44916 17153 44925 17187
rect 44925 17153 44959 17187
rect 44959 17153 44968 17187
rect 44916 17144 44968 17153
rect 39120 17076 39172 17128
rect 36636 17008 36688 17060
rect 36912 17008 36964 17060
rect 37188 17008 37240 17060
rect 37648 17008 37700 17060
rect 37924 17008 37976 17060
rect 38568 17008 38620 17060
rect 57428 17119 57480 17128
rect 57428 17085 57437 17119
rect 57437 17085 57471 17119
rect 57471 17085 57480 17119
rect 57428 17076 57480 17085
rect 40132 17008 40184 17060
rect 41420 17008 41472 17060
rect 41972 17008 42024 17060
rect 43536 17008 43588 17060
rect 43996 17008 44048 17060
rect 58256 17051 58308 17060
rect 58256 17017 58265 17051
rect 58265 17017 58299 17051
rect 58299 17017 58308 17051
rect 58256 17008 58308 17017
rect 2320 16940 2372 16992
rect 25964 16940 26016 16992
rect 33324 16940 33376 16992
rect 33968 16940 34020 16992
rect 36268 16940 36320 16992
rect 36544 16983 36596 16992
rect 36544 16949 36553 16983
rect 36553 16949 36587 16983
rect 36587 16949 36596 16983
rect 36544 16940 36596 16949
rect 36728 16940 36780 16992
rect 37740 16940 37792 16992
rect 38016 16940 38068 16992
rect 38108 16940 38160 16992
rect 40040 16940 40092 16992
rect 40408 16940 40460 16992
rect 40960 16983 41012 16992
rect 40960 16949 40969 16983
rect 40969 16949 41003 16983
rect 41003 16949 41012 16983
rect 40960 16940 41012 16949
rect 41328 16940 41380 16992
rect 43168 16940 43220 16992
rect 43904 16940 43956 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 25136 16736 25188 16788
rect 24584 16668 24636 16720
rect 25872 16668 25924 16720
rect 28356 16736 28408 16788
rect 29184 16736 29236 16788
rect 33784 16736 33836 16788
rect 34336 16736 34388 16788
rect 37280 16736 37332 16788
rect 37372 16736 37424 16788
rect 38016 16736 38068 16788
rect 27252 16600 27304 16652
rect 27436 16600 27488 16652
rect 24952 16532 25004 16584
rect 25412 16532 25464 16584
rect 27620 16532 27672 16584
rect 27896 16532 27948 16584
rect 28540 16575 28592 16584
rect 28540 16541 28549 16575
rect 28549 16541 28583 16575
rect 28583 16541 28592 16575
rect 28540 16532 28592 16541
rect 31576 16575 31628 16584
rect 31576 16541 31585 16575
rect 31585 16541 31619 16575
rect 31619 16541 31628 16575
rect 31576 16532 31628 16541
rect 32220 16575 32272 16584
rect 25320 16396 25372 16448
rect 25412 16396 25464 16448
rect 28356 16464 28408 16516
rect 27436 16396 27488 16448
rect 32220 16541 32229 16575
rect 32229 16541 32263 16575
rect 32263 16541 32272 16575
rect 32220 16532 32272 16541
rect 32404 16575 32456 16584
rect 32404 16541 32413 16575
rect 32413 16541 32447 16575
rect 32447 16541 32456 16575
rect 32404 16532 32456 16541
rect 33324 16668 33376 16720
rect 35532 16668 35584 16720
rect 38200 16711 38252 16720
rect 38200 16677 38209 16711
rect 38209 16677 38243 16711
rect 38243 16677 38252 16711
rect 38200 16668 38252 16677
rect 38384 16668 38436 16720
rect 36636 16600 36688 16652
rect 37648 16600 37700 16652
rect 38936 16736 38988 16788
rect 39304 16736 39356 16788
rect 41328 16736 41380 16788
rect 43628 16736 43680 16788
rect 44088 16736 44140 16788
rect 38844 16668 38896 16720
rect 33048 16575 33100 16584
rect 33048 16541 33057 16575
rect 33057 16541 33091 16575
rect 33091 16541 33100 16575
rect 33324 16575 33376 16584
rect 33048 16532 33100 16541
rect 33324 16541 33333 16575
rect 33333 16541 33367 16575
rect 33367 16541 33376 16575
rect 33324 16532 33376 16541
rect 33968 16575 34020 16584
rect 33968 16541 33977 16575
rect 33977 16541 34011 16575
rect 34011 16541 34020 16575
rect 33968 16532 34020 16541
rect 35256 16464 35308 16516
rect 36084 16532 36136 16584
rect 36452 16532 36504 16584
rect 37280 16532 37332 16584
rect 39488 16600 39540 16652
rect 40316 16643 40368 16652
rect 40316 16609 40325 16643
rect 40325 16609 40359 16643
rect 40359 16609 40368 16643
rect 40316 16600 40368 16609
rect 40776 16600 40828 16652
rect 37832 16464 37884 16516
rect 38844 16532 38896 16584
rect 38936 16532 38988 16584
rect 40132 16532 40184 16584
rect 34520 16396 34572 16448
rect 37648 16396 37700 16448
rect 40500 16575 40552 16584
rect 40500 16541 40509 16575
rect 40509 16541 40543 16575
rect 40543 16541 40552 16575
rect 40500 16532 40552 16541
rect 41236 16575 41288 16584
rect 41236 16541 41245 16575
rect 41245 16541 41279 16575
rect 41279 16541 41288 16575
rect 41236 16532 41288 16541
rect 41696 16532 41748 16584
rect 41420 16464 41472 16516
rect 42248 16575 42300 16584
rect 42248 16541 42257 16575
rect 42257 16541 42291 16575
rect 42291 16541 42300 16575
rect 43168 16600 43220 16652
rect 43352 16575 43404 16584
rect 42248 16532 42300 16541
rect 43352 16541 43361 16575
rect 43361 16541 43395 16575
rect 43395 16541 43404 16575
rect 43352 16532 43404 16541
rect 43444 16575 43496 16584
rect 43444 16541 43453 16575
rect 43453 16541 43487 16575
rect 43487 16541 43496 16575
rect 43628 16575 43680 16584
rect 43444 16532 43496 16541
rect 43628 16541 43637 16575
rect 43637 16541 43671 16575
rect 43671 16541 43680 16575
rect 43628 16532 43680 16541
rect 43720 16575 43772 16584
rect 43720 16541 43729 16575
rect 43729 16541 43763 16575
rect 43763 16541 43772 16575
rect 43720 16532 43772 16541
rect 44548 16575 44600 16584
rect 44548 16541 44557 16575
rect 44557 16541 44591 16575
rect 44591 16541 44600 16575
rect 44548 16532 44600 16541
rect 42340 16464 42392 16516
rect 42800 16396 42852 16448
rect 43628 16396 43680 16448
rect 43904 16439 43956 16448
rect 43904 16405 43913 16439
rect 43913 16405 43947 16439
rect 43947 16405 43956 16439
rect 43904 16396 43956 16405
rect 44088 16396 44140 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 25320 16192 25372 16244
rect 28356 16235 28408 16244
rect 25412 16124 25464 16176
rect 25964 16124 26016 16176
rect 28356 16201 28365 16235
rect 28365 16201 28399 16235
rect 28399 16201 28408 16235
rect 28356 16192 28408 16201
rect 28540 16192 28592 16244
rect 33600 16192 33652 16244
rect 34612 16235 34664 16244
rect 34612 16201 34621 16235
rect 34621 16201 34655 16235
rect 34655 16201 34664 16235
rect 34612 16192 34664 16201
rect 35348 16192 35400 16244
rect 37832 16192 37884 16244
rect 40500 16192 40552 16244
rect 40776 16192 40828 16244
rect 41512 16235 41564 16244
rect 41512 16201 41521 16235
rect 41521 16201 41555 16235
rect 41555 16201 41564 16235
rect 41512 16192 41564 16201
rect 43628 16192 43680 16244
rect 45468 16192 45520 16244
rect 28632 16124 28684 16176
rect 30104 16124 30156 16176
rect 25504 16099 25556 16108
rect 25504 16065 25513 16099
rect 25513 16065 25547 16099
rect 25547 16065 25556 16099
rect 25504 16056 25556 16065
rect 25872 16056 25924 16108
rect 27436 16099 27488 16108
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 24952 15988 25004 16040
rect 29092 16056 29144 16108
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 29920 16056 29972 16108
rect 30380 16099 30432 16108
rect 30380 16065 30389 16099
rect 30389 16065 30423 16099
rect 30423 16065 30432 16099
rect 30380 16056 30432 16065
rect 31116 16099 31168 16108
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 31116 16056 31168 16065
rect 31392 16056 31444 16108
rect 32496 16099 32548 16108
rect 32496 16065 32505 16099
rect 32505 16065 32539 16099
rect 32539 16065 32548 16099
rect 32496 16056 32548 16065
rect 33140 16056 33192 16108
rect 25044 15963 25096 15972
rect 25044 15929 25053 15963
rect 25053 15929 25087 15963
rect 25087 15929 25096 15963
rect 25044 15920 25096 15929
rect 26516 15852 26568 15904
rect 28816 16031 28868 16040
rect 28816 15997 28825 16031
rect 28825 15997 28859 16031
rect 28859 15997 28868 16031
rect 28816 15988 28868 15997
rect 27896 15920 27948 15972
rect 29368 15920 29420 15972
rect 33692 16056 33744 16108
rect 34428 15988 34480 16040
rect 35440 16056 35492 16108
rect 36544 16124 36596 16176
rect 40316 16124 40368 16176
rect 40868 16124 40920 16176
rect 37004 16056 37056 16108
rect 37556 16056 37608 16108
rect 37924 16099 37976 16108
rect 37924 16065 37933 16099
rect 37933 16065 37967 16099
rect 37967 16065 37976 16099
rect 37924 16056 37976 16065
rect 39304 16099 39356 16108
rect 39304 16065 39313 16099
rect 39313 16065 39347 16099
rect 39347 16065 39356 16099
rect 39304 16056 39356 16065
rect 39488 16099 39540 16108
rect 39488 16065 39497 16099
rect 39497 16065 39531 16099
rect 39531 16065 39540 16099
rect 39488 16056 39540 16065
rect 40408 16099 40460 16108
rect 40408 16065 40417 16099
rect 40417 16065 40451 16099
rect 40451 16065 40460 16099
rect 40408 16056 40460 16065
rect 41420 16056 41472 16108
rect 35808 15988 35860 16040
rect 36544 16031 36596 16040
rect 36544 15997 36553 16031
rect 36553 15997 36587 16031
rect 36587 15997 36596 16031
rect 36544 15988 36596 15997
rect 39580 16031 39632 16040
rect 39580 15997 39589 16031
rect 39589 15997 39623 16031
rect 39623 15997 39632 16031
rect 39580 15988 39632 15997
rect 40868 15988 40920 16040
rect 43812 16124 43864 16176
rect 41880 16099 41932 16108
rect 41880 16065 41889 16099
rect 41889 16065 41923 16099
rect 41923 16065 41932 16099
rect 41880 16056 41932 16065
rect 43444 16056 43496 16108
rect 43720 16056 43772 16108
rect 44272 16124 44324 16176
rect 45192 16099 45244 16108
rect 45192 16065 45201 16099
rect 45201 16065 45235 16099
rect 45235 16065 45244 16099
rect 45192 16056 45244 16065
rect 43076 15988 43128 16040
rect 28632 15852 28684 15904
rect 29184 15852 29236 15904
rect 31944 15852 31996 15904
rect 32588 15895 32640 15904
rect 32588 15861 32597 15895
rect 32597 15861 32631 15895
rect 32631 15861 32640 15895
rect 32588 15852 32640 15861
rect 33876 15852 33928 15904
rect 34336 15852 34388 15904
rect 34796 15895 34848 15904
rect 34796 15861 34805 15895
rect 34805 15861 34839 15895
rect 34839 15861 34848 15895
rect 36176 15920 36228 15972
rect 34796 15852 34848 15861
rect 35624 15852 35676 15904
rect 36728 15895 36780 15904
rect 36728 15861 36737 15895
rect 36737 15861 36771 15895
rect 36771 15861 36780 15895
rect 36728 15852 36780 15861
rect 36912 15895 36964 15904
rect 36912 15861 36921 15895
rect 36921 15861 36955 15895
rect 36955 15861 36964 15895
rect 36912 15852 36964 15861
rect 37372 15852 37424 15904
rect 37924 15852 37976 15904
rect 38108 15852 38160 15904
rect 39120 15895 39172 15904
rect 39120 15861 39129 15895
rect 39129 15861 39163 15895
rect 39163 15861 39172 15895
rect 39120 15852 39172 15861
rect 40960 15920 41012 15972
rect 44456 15988 44508 16040
rect 39764 15852 39816 15904
rect 40776 15852 40828 15904
rect 43628 15895 43680 15904
rect 43628 15861 43637 15895
rect 43637 15861 43671 15895
rect 43671 15861 43680 15895
rect 43628 15852 43680 15861
rect 45100 15895 45152 15904
rect 45100 15861 45109 15895
rect 45109 15861 45143 15895
rect 45143 15861 45152 15895
rect 45100 15852 45152 15861
rect 45652 15895 45704 15904
rect 45652 15861 45661 15895
rect 45661 15861 45695 15895
rect 45695 15861 45704 15895
rect 45652 15852 45704 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 28540 15648 28592 15700
rect 29276 15648 29328 15700
rect 31576 15691 31628 15700
rect 31576 15657 31585 15691
rect 31585 15657 31619 15691
rect 31619 15657 31628 15691
rect 31576 15648 31628 15657
rect 33232 15648 33284 15700
rect 34796 15648 34848 15700
rect 35348 15648 35400 15700
rect 40224 15691 40276 15700
rect 40224 15657 40233 15691
rect 40233 15657 40267 15691
rect 40267 15657 40276 15691
rect 40224 15648 40276 15657
rect 41144 15691 41196 15700
rect 41144 15657 41153 15691
rect 41153 15657 41187 15691
rect 41187 15657 41196 15691
rect 41144 15648 41196 15657
rect 42064 15648 42116 15700
rect 25688 15580 25740 15632
rect 34060 15580 34112 15632
rect 36452 15580 36504 15632
rect 36912 15580 36964 15632
rect 42616 15580 42668 15632
rect 26884 15512 26936 15564
rect 29368 15512 29420 15564
rect 30656 15512 30708 15564
rect 24308 15444 24360 15496
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 26424 15444 26476 15496
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 28816 15444 28868 15496
rect 29092 15487 29144 15496
rect 29092 15453 29101 15487
rect 29101 15453 29135 15487
rect 29135 15453 29144 15487
rect 32496 15512 32548 15564
rect 31944 15487 31996 15496
rect 29092 15444 29144 15453
rect 23940 15376 23992 15428
rect 26148 15376 26200 15428
rect 26884 15376 26936 15428
rect 29644 15376 29696 15428
rect 30656 15419 30708 15428
rect 23480 15351 23532 15360
rect 23480 15317 23489 15351
rect 23489 15317 23523 15351
rect 23523 15317 23532 15351
rect 23480 15308 23532 15317
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 26976 15308 27028 15317
rect 29000 15308 29052 15360
rect 30656 15385 30665 15419
rect 30665 15385 30699 15419
rect 30699 15385 30708 15419
rect 30656 15376 30708 15385
rect 31944 15453 31953 15487
rect 31953 15453 31987 15487
rect 31987 15453 31996 15487
rect 31944 15444 31996 15453
rect 32588 15487 32640 15496
rect 32588 15453 32597 15487
rect 32597 15453 32631 15487
rect 32631 15453 32640 15487
rect 32588 15444 32640 15453
rect 33140 15512 33192 15564
rect 33692 15512 33744 15564
rect 35624 15512 35676 15564
rect 33324 15444 33376 15496
rect 33968 15487 34020 15496
rect 33968 15453 33977 15487
rect 33977 15453 34011 15487
rect 34011 15453 34020 15487
rect 33968 15444 34020 15453
rect 31024 15308 31076 15360
rect 33048 15308 33100 15360
rect 34704 15376 34756 15428
rect 35992 15444 36044 15496
rect 36360 15444 36412 15496
rect 36912 15444 36964 15496
rect 40132 15512 40184 15564
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 42800 15512 42852 15564
rect 43904 15555 43956 15564
rect 43904 15521 43913 15555
rect 43913 15521 43947 15555
rect 43947 15521 43956 15555
rect 43904 15512 43956 15521
rect 45100 15512 45152 15564
rect 37280 15444 37332 15496
rect 35900 15376 35952 15428
rect 38292 15444 38344 15496
rect 41144 15444 41196 15496
rect 42524 15487 42576 15496
rect 42524 15453 42533 15487
rect 42533 15453 42567 15487
rect 42567 15453 42576 15487
rect 42524 15444 42576 15453
rect 43812 15487 43864 15496
rect 36176 15308 36228 15360
rect 36360 15308 36412 15360
rect 38108 15376 38160 15428
rect 43812 15453 43821 15487
rect 43821 15453 43855 15487
rect 43855 15453 43864 15487
rect 43812 15444 43864 15453
rect 45468 15487 45520 15496
rect 45468 15453 45477 15487
rect 45477 15453 45511 15487
rect 45511 15453 45520 15487
rect 45468 15444 45520 15453
rect 45652 15487 45704 15496
rect 45652 15453 45661 15487
rect 45661 15453 45695 15487
rect 45695 15453 45704 15487
rect 45652 15444 45704 15453
rect 45836 15487 45888 15496
rect 45836 15453 45845 15487
rect 45845 15453 45879 15487
rect 45879 15453 45888 15487
rect 45836 15444 45888 15453
rect 38844 15308 38896 15360
rect 40040 15351 40092 15360
rect 40040 15317 40049 15351
rect 40049 15317 40083 15351
rect 40083 15317 40092 15351
rect 40040 15308 40092 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 25596 15104 25648 15156
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 27252 15036 27304 15088
rect 26976 14968 27028 15020
rect 24216 14875 24268 14884
rect 24216 14841 24225 14875
rect 24225 14841 24259 14875
rect 24259 14841 24268 14875
rect 24216 14832 24268 14841
rect 26148 14900 26200 14952
rect 27160 14943 27212 14952
rect 27160 14909 27169 14943
rect 27169 14909 27203 14943
rect 27203 14909 27212 14943
rect 27160 14900 27212 14909
rect 27988 14968 28040 15020
rect 29184 15104 29236 15156
rect 30288 15104 30340 15156
rect 31300 15104 31352 15156
rect 32588 15104 32640 15156
rect 33048 15147 33100 15156
rect 33048 15113 33057 15147
rect 33057 15113 33091 15147
rect 33091 15113 33100 15147
rect 33048 15104 33100 15113
rect 33692 15147 33744 15156
rect 33692 15113 33701 15147
rect 33701 15113 33735 15147
rect 33735 15113 33744 15147
rect 33692 15104 33744 15113
rect 35256 15104 35308 15156
rect 36176 15104 36228 15156
rect 29000 15036 29052 15088
rect 27804 14900 27856 14952
rect 26424 14832 26476 14884
rect 28172 14832 28224 14884
rect 28908 15011 28960 15020
rect 28908 14977 28917 15011
rect 28917 14977 28951 15011
rect 28951 14977 28960 15011
rect 30564 15036 30616 15088
rect 28908 14968 28960 14977
rect 30656 14968 30708 15020
rect 32772 15036 32824 15088
rect 36360 15104 36412 15156
rect 36452 15104 36504 15156
rect 42432 15104 42484 15156
rect 44088 15147 44140 15156
rect 44088 15113 44097 15147
rect 44097 15113 44131 15147
rect 44131 15113 44140 15147
rect 44088 15104 44140 15113
rect 32680 15011 32732 15020
rect 32220 14900 32272 14952
rect 32680 14977 32689 15011
rect 32689 14977 32723 15011
rect 32723 14977 32732 15011
rect 32680 14968 32732 14977
rect 33048 14968 33100 15020
rect 34704 14968 34756 15020
rect 35256 15011 35308 15020
rect 35256 14977 35265 15011
rect 35265 14977 35299 15011
rect 35299 14977 35308 15011
rect 35256 14968 35308 14977
rect 35440 15011 35492 15020
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 35624 15011 35676 15020
rect 35624 14977 35633 15011
rect 35633 14977 35667 15011
rect 35667 14977 35676 15011
rect 35624 14968 35676 14977
rect 35900 14968 35952 15020
rect 36084 15011 36136 15020
rect 36084 14977 36093 15011
rect 36093 14977 36127 15011
rect 36127 14977 36136 15011
rect 36084 14968 36136 14977
rect 36268 15011 36320 15020
rect 36268 14977 36277 15011
rect 36277 14977 36311 15011
rect 36311 14977 36320 15011
rect 36268 14968 36320 14977
rect 36912 15036 36964 15088
rect 38568 15036 38620 15088
rect 37740 14968 37792 15020
rect 38476 14968 38528 15020
rect 33140 14900 33192 14952
rect 35348 14943 35400 14952
rect 35348 14909 35357 14943
rect 35357 14909 35391 14943
rect 35391 14909 35400 14943
rect 35348 14900 35400 14909
rect 39028 15011 39080 15020
rect 39028 14977 39037 15011
rect 39037 14977 39071 15011
rect 39071 14977 39080 15011
rect 39028 14968 39080 14977
rect 39304 14968 39356 15020
rect 39580 14968 39632 15020
rect 40040 15011 40092 15020
rect 40040 14977 40049 15011
rect 40049 14977 40083 15011
rect 40083 14977 40092 15011
rect 40040 14968 40092 14977
rect 40684 15011 40736 15020
rect 40684 14977 40693 15011
rect 40693 14977 40727 15011
rect 40727 14977 40736 15011
rect 40684 14968 40736 14977
rect 39672 14900 39724 14952
rect 40224 14900 40276 14952
rect 40408 14900 40460 14952
rect 32772 14875 32824 14884
rect 32772 14841 32777 14875
rect 32777 14841 32811 14875
rect 32811 14841 32824 14875
rect 32772 14832 32824 14841
rect 32956 14832 33008 14884
rect 36084 14832 36136 14884
rect 37372 14832 37424 14884
rect 38568 14875 38620 14884
rect 29644 14807 29696 14816
rect 29644 14773 29653 14807
rect 29653 14773 29687 14807
rect 29687 14773 29696 14807
rect 29644 14764 29696 14773
rect 34336 14807 34388 14816
rect 34336 14773 34345 14807
rect 34345 14773 34379 14807
rect 34379 14773 34388 14807
rect 34336 14764 34388 14773
rect 35348 14764 35400 14816
rect 38568 14841 38577 14875
rect 38577 14841 38611 14875
rect 38611 14841 38620 14875
rect 38568 14832 38620 14841
rect 41512 15036 41564 15088
rect 41604 15011 41656 15020
rect 41604 14977 41613 15011
rect 41613 14977 41647 15011
rect 41647 14977 41656 15011
rect 41604 14968 41656 14977
rect 41788 15011 41840 15020
rect 41788 14977 41797 15011
rect 41797 14977 41831 15011
rect 41831 14977 41840 15011
rect 41788 14968 41840 14977
rect 42156 14968 42208 15020
rect 42708 15011 42760 15020
rect 42708 14977 42717 15011
rect 42717 14977 42751 15011
rect 42751 14977 42760 15011
rect 42708 14968 42760 14977
rect 42800 14968 42852 15020
rect 44456 15011 44508 15020
rect 44456 14977 44465 15011
rect 44465 14977 44499 15011
rect 44499 14977 44508 15011
rect 44456 14968 44508 14977
rect 41972 14943 42024 14952
rect 41972 14909 41981 14943
rect 41981 14909 42015 14943
rect 42015 14909 42024 14943
rect 41972 14900 42024 14909
rect 42892 14900 42944 14952
rect 38936 14764 38988 14816
rect 39304 14764 39356 14816
rect 41052 14764 41104 14816
rect 42708 14832 42760 14884
rect 43352 14875 43404 14884
rect 43352 14841 43361 14875
rect 43361 14841 43395 14875
rect 43395 14841 43404 14875
rect 43352 14832 43404 14841
rect 41696 14764 41748 14816
rect 42156 14764 42208 14816
rect 43812 14764 43864 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 26148 14560 26200 14612
rect 26884 14560 26936 14612
rect 27528 14560 27580 14612
rect 27712 14560 27764 14612
rect 27988 14603 28040 14612
rect 27988 14569 27997 14603
rect 27997 14569 28031 14603
rect 28031 14569 28040 14603
rect 27988 14560 28040 14569
rect 29184 14603 29236 14612
rect 29184 14569 29193 14603
rect 29193 14569 29227 14603
rect 29227 14569 29236 14603
rect 29184 14560 29236 14569
rect 30012 14560 30064 14612
rect 31392 14603 31444 14612
rect 31392 14569 31401 14603
rect 31401 14569 31435 14603
rect 31435 14569 31444 14603
rect 31392 14560 31444 14569
rect 33968 14560 34020 14612
rect 36544 14560 36596 14612
rect 27620 14492 27672 14544
rect 34980 14492 35032 14544
rect 28172 14467 28224 14476
rect 28172 14433 28181 14467
rect 28181 14433 28215 14467
rect 28215 14433 28224 14467
rect 28172 14424 28224 14433
rect 29000 14424 29052 14476
rect 31208 14424 31260 14476
rect 35716 14424 35768 14476
rect 24216 14356 24268 14408
rect 25596 14356 25648 14408
rect 28908 14356 28960 14408
rect 30564 14399 30616 14408
rect 30564 14365 30573 14399
rect 30573 14365 30607 14399
rect 30607 14365 30616 14399
rect 30564 14356 30616 14365
rect 29184 14288 29236 14340
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 31576 14356 31628 14365
rect 34060 14399 34112 14408
rect 34060 14365 34069 14399
rect 34069 14365 34103 14399
rect 34103 14365 34112 14399
rect 34060 14356 34112 14365
rect 34336 14399 34388 14408
rect 34336 14365 34345 14399
rect 34345 14365 34379 14399
rect 34379 14365 34388 14399
rect 34336 14356 34388 14365
rect 32772 14331 32824 14340
rect 32772 14297 32781 14331
rect 32781 14297 32815 14331
rect 32815 14297 32824 14331
rect 32772 14288 32824 14297
rect 32956 14331 33008 14340
rect 32956 14297 32965 14331
rect 32965 14297 32999 14331
rect 32999 14297 33008 14331
rect 32956 14288 33008 14297
rect 35992 14492 36044 14544
rect 36268 14424 36320 14476
rect 36084 14399 36136 14408
rect 36084 14365 36093 14399
rect 36093 14365 36127 14399
rect 36127 14365 36136 14399
rect 36084 14356 36136 14365
rect 36912 14356 36964 14408
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 25412 14220 25464 14272
rect 31024 14220 31076 14272
rect 33876 14263 33928 14272
rect 33876 14229 33885 14263
rect 33885 14229 33919 14263
rect 33919 14229 33928 14263
rect 33876 14220 33928 14229
rect 36360 14288 36412 14340
rect 39304 14560 39356 14612
rect 39580 14560 39632 14612
rect 39856 14560 39908 14612
rect 43444 14560 43496 14612
rect 43812 14560 43864 14612
rect 38292 14492 38344 14544
rect 38476 14492 38528 14544
rect 43352 14492 43404 14544
rect 37556 14356 37608 14408
rect 38384 14424 38436 14476
rect 39488 14424 39540 14476
rect 40684 14467 40736 14476
rect 40684 14433 40693 14467
rect 40693 14433 40727 14467
rect 40727 14433 40736 14467
rect 40684 14424 40736 14433
rect 37832 14399 37884 14408
rect 37832 14365 37841 14399
rect 37841 14365 37875 14399
rect 37875 14365 37884 14399
rect 37832 14356 37884 14365
rect 38016 14288 38068 14340
rect 38200 14288 38252 14340
rect 38568 14288 38620 14340
rect 37648 14263 37700 14272
rect 37648 14229 37657 14263
rect 37657 14229 37691 14263
rect 37691 14229 37700 14263
rect 37648 14220 37700 14229
rect 38292 14220 38344 14272
rect 38660 14220 38712 14272
rect 38936 14288 38988 14340
rect 39212 14331 39264 14340
rect 39212 14297 39221 14331
rect 39221 14297 39255 14331
rect 39255 14297 39264 14331
rect 39212 14288 39264 14297
rect 40960 14356 41012 14408
rect 41052 14399 41104 14408
rect 41052 14365 41061 14399
rect 41061 14365 41095 14399
rect 41095 14365 41104 14399
rect 41972 14424 42024 14476
rect 42156 14467 42208 14476
rect 42156 14433 42165 14467
rect 42165 14433 42199 14467
rect 42199 14433 42208 14467
rect 42156 14424 42208 14433
rect 41052 14356 41104 14365
rect 41604 14356 41656 14408
rect 42616 14356 42668 14408
rect 43536 14356 43588 14408
rect 44456 14356 44508 14408
rect 45376 14560 45428 14612
rect 41328 14220 41380 14272
rect 44272 14220 44324 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 23756 14016 23808 14068
rect 23848 14016 23900 14068
rect 24676 13948 24728 14000
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 23480 13880 23532 13932
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 27804 14059 27856 14068
rect 25412 13948 25464 14000
rect 25504 13923 25556 13932
rect 23848 13812 23900 13864
rect 24308 13855 24360 13864
rect 24308 13821 24317 13855
rect 24317 13821 24351 13855
rect 24351 13821 24360 13855
rect 24308 13812 24360 13821
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 25504 13889 25513 13923
rect 25513 13889 25547 13923
rect 25547 13889 25556 13923
rect 25504 13880 25556 13889
rect 25780 13880 25832 13932
rect 27804 14025 27813 14059
rect 27813 14025 27847 14059
rect 27847 14025 27856 14059
rect 27804 14016 27856 14025
rect 29644 14059 29696 14068
rect 29184 13948 29236 14000
rect 27252 13880 27304 13932
rect 28540 13923 28592 13932
rect 28540 13889 28549 13923
rect 28549 13889 28583 13923
rect 28583 13889 28592 13923
rect 28540 13880 28592 13889
rect 29644 14025 29653 14059
rect 29653 14025 29687 14059
rect 29687 14025 29696 14059
rect 29644 14016 29696 14025
rect 30840 14016 30892 14068
rect 31208 14059 31260 14068
rect 31208 14025 31217 14059
rect 31217 14025 31251 14059
rect 31251 14025 31260 14059
rect 31208 14016 31260 14025
rect 32956 14016 33008 14068
rect 34428 14016 34480 14068
rect 36452 14059 36504 14068
rect 36452 14025 36461 14059
rect 36461 14025 36495 14059
rect 36495 14025 36504 14059
rect 36452 14016 36504 14025
rect 36544 14016 36596 14068
rect 40316 14016 40368 14068
rect 40776 14016 40828 14068
rect 31852 13948 31904 14000
rect 30564 13880 30616 13932
rect 31116 13880 31168 13932
rect 31300 13923 31352 13932
rect 31300 13889 31309 13923
rect 31309 13889 31343 13923
rect 31343 13889 31352 13923
rect 31300 13880 31352 13889
rect 33048 13923 33100 13932
rect 33048 13889 33057 13923
rect 33057 13889 33091 13923
rect 33091 13889 33100 13923
rect 33048 13880 33100 13889
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 33784 13880 33836 13932
rect 34980 13923 35032 13932
rect 34980 13889 34989 13923
rect 34989 13889 35023 13923
rect 35023 13889 35032 13923
rect 34980 13880 35032 13889
rect 35256 13923 35308 13932
rect 35256 13889 35265 13923
rect 35265 13889 35299 13923
rect 35299 13889 35308 13923
rect 35256 13880 35308 13889
rect 35348 13923 35400 13932
rect 35348 13889 35357 13923
rect 35357 13889 35391 13923
rect 35391 13889 35400 13923
rect 35716 13948 35768 14000
rect 37832 13948 37884 14000
rect 35348 13880 35400 13889
rect 36636 13880 36688 13932
rect 37280 13880 37332 13932
rect 37924 13923 37976 13932
rect 26792 13812 26844 13864
rect 24032 13744 24084 13796
rect 24768 13744 24820 13796
rect 27988 13812 28040 13864
rect 23388 13676 23440 13728
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 26240 13676 26292 13728
rect 32864 13812 32916 13864
rect 33140 13855 33192 13864
rect 33140 13821 33149 13855
rect 33149 13821 33183 13855
rect 33183 13821 33192 13855
rect 33140 13812 33192 13821
rect 34060 13812 34112 13864
rect 37648 13812 37700 13864
rect 37924 13889 37933 13923
rect 37933 13889 37967 13923
rect 37967 13889 37976 13923
rect 37924 13880 37976 13889
rect 38384 13948 38436 14000
rect 39212 13948 39264 14000
rect 38108 13880 38160 13932
rect 41144 13948 41196 14000
rect 41880 14016 41932 14068
rect 42064 14016 42116 14068
rect 44180 14016 44232 14068
rect 42984 13991 43036 14000
rect 42984 13957 42993 13991
rect 42993 13957 43027 13991
rect 43027 13957 43036 13991
rect 42984 13948 43036 13957
rect 44456 13948 44508 14000
rect 40684 13923 40736 13932
rect 40684 13889 40693 13923
rect 40693 13889 40727 13923
rect 40727 13889 40736 13923
rect 40684 13880 40736 13889
rect 40960 13880 41012 13932
rect 41328 13880 41380 13932
rect 41972 13880 42024 13932
rect 42616 13923 42668 13932
rect 42616 13889 42625 13923
rect 42625 13889 42659 13923
rect 42659 13889 42668 13923
rect 42616 13880 42668 13889
rect 43536 13880 43588 13932
rect 44088 13923 44140 13932
rect 44088 13889 44097 13923
rect 44097 13889 44131 13923
rect 44131 13889 44140 13923
rect 44088 13880 44140 13889
rect 44272 13923 44324 13932
rect 44272 13889 44281 13923
rect 44281 13889 44315 13923
rect 44315 13889 44324 13923
rect 44272 13880 44324 13889
rect 44364 13923 44416 13932
rect 44364 13889 44373 13923
rect 44373 13889 44407 13923
rect 44407 13889 44416 13923
rect 44364 13880 44416 13889
rect 44640 13880 44692 13932
rect 45468 13880 45520 13932
rect 40316 13812 40368 13864
rect 41144 13812 41196 13864
rect 42708 13812 42760 13864
rect 45744 13812 45796 13864
rect 30380 13744 30432 13796
rect 30656 13744 30708 13796
rect 43628 13744 43680 13796
rect 44456 13744 44508 13796
rect 45652 13787 45704 13796
rect 45652 13753 45661 13787
rect 45661 13753 45695 13787
rect 45695 13753 45704 13787
rect 45652 13744 45704 13753
rect 33876 13676 33928 13728
rect 34796 13719 34848 13728
rect 34796 13685 34805 13719
rect 34805 13685 34839 13719
rect 34839 13685 34848 13719
rect 34796 13676 34848 13685
rect 36360 13676 36412 13728
rect 37740 13719 37792 13728
rect 37740 13685 37749 13719
rect 37749 13685 37783 13719
rect 37783 13685 37792 13719
rect 37740 13676 37792 13685
rect 39304 13676 39356 13728
rect 41236 13676 41288 13728
rect 41512 13719 41564 13728
rect 41512 13685 41521 13719
rect 41521 13685 41555 13719
rect 41555 13685 41564 13719
rect 41512 13676 41564 13685
rect 42156 13676 42208 13728
rect 45008 13719 45060 13728
rect 45008 13685 45017 13719
rect 45017 13685 45051 13719
rect 45051 13685 45060 13719
rect 45008 13676 45060 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 28540 13472 28592 13524
rect 30472 13472 30524 13524
rect 31024 13515 31076 13524
rect 31024 13481 31033 13515
rect 31033 13481 31067 13515
rect 31067 13481 31076 13515
rect 31024 13472 31076 13481
rect 32772 13472 32824 13524
rect 33048 13472 33100 13524
rect 35532 13472 35584 13524
rect 36452 13515 36504 13524
rect 36452 13481 36461 13515
rect 36461 13481 36495 13515
rect 36495 13481 36504 13515
rect 36452 13472 36504 13481
rect 26792 13447 26844 13456
rect 26792 13413 26801 13447
rect 26801 13413 26835 13447
rect 26835 13413 26844 13447
rect 26792 13404 26844 13413
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 24400 13268 24452 13320
rect 25872 13268 25924 13320
rect 26240 13268 26292 13320
rect 26332 13311 26384 13320
rect 26332 13277 26341 13311
rect 26341 13277 26375 13311
rect 26375 13277 26384 13311
rect 32496 13404 32548 13456
rect 32956 13404 33008 13456
rect 35624 13404 35676 13456
rect 36268 13404 36320 13456
rect 36636 13404 36688 13456
rect 27252 13379 27304 13388
rect 27252 13345 27261 13379
rect 27261 13345 27295 13379
rect 27295 13345 27304 13379
rect 27252 13336 27304 13345
rect 27896 13336 27948 13388
rect 31024 13336 31076 13388
rect 33232 13336 33284 13388
rect 27160 13311 27212 13320
rect 26332 13268 26384 13277
rect 27160 13277 27169 13311
rect 27169 13277 27203 13311
rect 27203 13277 27212 13311
rect 27160 13268 27212 13277
rect 23572 13175 23624 13184
rect 23572 13141 23581 13175
rect 23581 13141 23615 13175
rect 23615 13141 23624 13175
rect 23572 13132 23624 13141
rect 24676 13132 24728 13184
rect 25412 13175 25464 13184
rect 25412 13141 25421 13175
rect 25421 13141 25455 13175
rect 25455 13141 25464 13175
rect 25412 13132 25464 13141
rect 27252 13200 27304 13252
rect 26424 13132 26476 13184
rect 26884 13132 26936 13184
rect 27528 13132 27580 13184
rect 29460 13268 29512 13320
rect 30196 13268 30248 13320
rect 30380 13268 30432 13320
rect 30748 13268 30800 13320
rect 31300 13311 31352 13320
rect 31300 13277 31309 13311
rect 31309 13277 31343 13311
rect 31343 13277 31352 13311
rect 31300 13268 31352 13277
rect 33048 13268 33100 13320
rect 33968 13336 34020 13388
rect 34244 13379 34296 13388
rect 34244 13345 34253 13379
rect 34253 13345 34287 13379
rect 34287 13345 34296 13379
rect 34244 13336 34296 13345
rect 36728 13379 36780 13388
rect 36728 13345 36737 13379
rect 36737 13345 36771 13379
rect 36771 13345 36780 13379
rect 36728 13336 36780 13345
rect 37740 13404 37792 13456
rect 39028 13472 39080 13524
rect 40040 13472 40092 13524
rect 40776 13472 40828 13524
rect 30564 13200 30616 13252
rect 30932 13200 30984 13252
rect 32864 13243 32916 13252
rect 32864 13209 32873 13243
rect 32873 13209 32907 13243
rect 32907 13209 32916 13243
rect 32864 13200 32916 13209
rect 34428 13268 34480 13320
rect 37464 13336 37516 13388
rect 37740 13311 37792 13320
rect 34520 13200 34572 13252
rect 28540 13132 28592 13184
rect 30840 13132 30892 13184
rect 33140 13132 33192 13184
rect 37740 13277 37749 13311
rect 37749 13277 37783 13311
rect 37783 13277 37792 13311
rect 37740 13268 37792 13277
rect 38936 13404 38988 13456
rect 39212 13404 39264 13456
rect 43260 13447 43312 13456
rect 43260 13413 43269 13447
rect 43269 13413 43303 13447
rect 43303 13413 43312 13447
rect 43260 13404 43312 13413
rect 38752 13336 38804 13388
rect 38844 13336 38896 13388
rect 40500 13336 40552 13388
rect 42064 13336 42116 13388
rect 40316 13311 40368 13320
rect 40316 13277 40325 13311
rect 40325 13277 40359 13311
rect 40359 13277 40368 13311
rect 40316 13268 40368 13277
rect 38752 13243 38804 13252
rect 38752 13209 38780 13243
rect 38780 13209 38804 13243
rect 38936 13243 38988 13252
rect 38752 13200 38804 13209
rect 38936 13209 38945 13243
rect 38945 13209 38979 13243
rect 38979 13209 38988 13243
rect 38936 13200 38988 13209
rect 40408 13243 40460 13252
rect 40408 13209 40417 13243
rect 40417 13209 40451 13243
rect 40451 13209 40460 13243
rect 40408 13200 40460 13209
rect 37740 13132 37792 13184
rect 37832 13132 37884 13184
rect 39672 13132 39724 13184
rect 40132 13132 40184 13184
rect 40500 13175 40552 13184
rect 40500 13141 40509 13175
rect 40509 13141 40543 13175
rect 40543 13141 40552 13175
rect 40500 13132 40552 13141
rect 40776 13311 40828 13320
rect 40776 13277 40785 13311
rect 40785 13277 40819 13311
rect 40819 13277 40828 13311
rect 40776 13268 40828 13277
rect 40960 13268 41012 13320
rect 41052 13200 41104 13252
rect 41880 13268 41932 13320
rect 42156 13311 42208 13320
rect 42156 13277 42165 13311
rect 42165 13277 42199 13311
rect 42199 13277 42208 13311
rect 42156 13268 42208 13277
rect 42800 13336 42852 13388
rect 42432 13311 42484 13320
rect 42432 13277 42441 13311
rect 42441 13277 42475 13311
rect 42475 13277 42484 13311
rect 42432 13268 42484 13277
rect 43444 13311 43496 13320
rect 43444 13277 43453 13311
rect 43453 13277 43487 13311
rect 43487 13277 43496 13311
rect 43444 13268 43496 13277
rect 43996 13311 44048 13320
rect 43996 13277 44005 13311
rect 44005 13277 44039 13311
rect 44039 13277 44048 13311
rect 43996 13268 44048 13277
rect 44180 13311 44232 13320
rect 44180 13277 44189 13311
rect 44189 13277 44223 13311
rect 44223 13277 44232 13311
rect 44180 13268 44232 13277
rect 42248 13132 42300 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 25872 12971 25924 12980
rect 25872 12937 25881 12971
rect 25881 12937 25915 12971
rect 25915 12937 25924 12971
rect 25872 12928 25924 12937
rect 26148 12928 26200 12980
rect 30472 12928 30524 12980
rect 33140 12928 33192 12980
rect 33508 12928 33560 12980
rect 35348 12928 35400 12980
rect 36636 12971 36688 12980
rect 36636 12937 36645 12971
rect 36645 12937 36679 12971
rect 36679 12937 36688 12971
rect 36636 12928 36688 12937
rect 38292 12971 38344 12980
rect 38292 12937 38301 12971
rect 38301 12937 38335 12971
rect 38335 12937 38344 12971
rect 38292 12928 38344 12937
rect 26424 12860 26476 12912
rect 27252 12903 27304 12912
rect 27252 12869 27261 12903
rect 27261 12869 27295 12903
rect 27295 12869 27304 12903
rect 27252 12860 27304 12869
rect 27528 12860 27580 12912
rect 23848 12792 23900 12844
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 29092 12860 29144 12912
rect 30564 12860 30616 12912
rect 30656 12860 30708 12912
rect 31116 12903 31168 12912
rect 31116 12869 31125 12903
rect 31125 12869 31159 12903
rect 31159 12869 31168 12903
rect 31116 12860 31168 12869
rect 31300 12860 31352 12912
rect 29000 12792 29052 12844
rect 29184 12792 29236 12844
rect 30748 12835 30800 12844
rect 30748 12801 30757 12835
rect 30757 12801 30791 12835
rect 30791 12801 30800 12835
rect 30748 12792 30800 12801
rect 31576 12835 31628 12844
rect 31576 12801 31585 12835
rect 31585 12801 31619 12835
rect 31619 12801 31628 12835
rect 31576 12792 31628 12801
rect 34796 12860 34848 12912
rect 28540 12724 28592 12776
rect 30196 12724 30248 12776
rect 30840 12724 30892 12776
rect 31392 12724 31444 12776
rect 32956 12792 33008 12844
rect 34428 12835 34480 12844
rect 34428 12801 34437 12835
rect 34437 12801 34471 12835
rect 34471 12801 34480 12835
rect 34428 12792 34480 12801
rect 32588 12767 32640 12776
rect 32588 12733 32597 12767
rect 32597 12733 32631 12767
rect 32631 12733 32640 12767
rect 32588 12724 32640 12733
rect 35532 12792 35584 12844
rect 35900 12860 35952 12912
rect 38752 12928 38804 12980
rect 40316 12928 40368 12980
rect 40500 12928 40552 12980
rect 44456 12928 44508 12980
rect 38936 12860 38988 12912
rect 40868 12903 40920 12912
rect 36176 12792 36228 12844
rect 36728 12835 36780 12844
rect 36728 12801 36737 12835
rect 36737 12801 36771 12835
rect 36771 12801 36780 12835
rect 36728 12792 36780 12801
rect 36912 12792 36964 12844
rect 37832 12835 37884 12844
rect 36820 12724 36872 12776
rect 37832 12801 37841 12835
rect 37841 12801 37875 12835
rect 37875 12801 37884 12835
rect 37832 12792 37884 12801
rect 39672 12835 39724 12844
rect 39672 12801 39681 12835
rect 39681 12801 39715 12835
rect 39715 12801 39724 12835
rect 39672 12792 39724 12801
rect 40868 12869 40877 12903
rect 40877 12869 40911 12903
rect 40911 12869 40920 12903
rect 40868 12860 40920 12869
rect 40960 12792 41012 12844
rect 41144 12860 41196 12912
rect 41880 12860 41932 12912
rect 41236 12835 41288 12844
rect 41236 12801 41245 12835
rect 41245 12801 41279 12835
rect 41279 12801 41288 12835
rect 41236 12792 41288 12801
rect 41512 12792 41564 12844
rect 30012 12656 30064 12708
rect 34520 12656 34572 12708
rect 35808 12699 35860 12708
rect 35808 12665 35817 12699
rect 35817 12665 35851 12699
rect 35851 12665 35860 12699
rect 35808 12656 35860 12665
rect 24952 12631 25004 12640
rect 24952 12597 24961 12631
rect 24961 12597 24995 12631
rect 24995 12597 25004 12631
rect 24952 12588 25004 12597
rect 26332 12588 26384 12640
rect 27896 12588 27948 12640
rect 29920 12588 29972 12640
rect 31300 12588 31352 12640
rect 34704 12631 34756 12640
rect 34704 12597 34713 12631
rect 34713 12597 34747 12631
rect 34747 12597 34756 12631
rect 34704 12588 34756 12597
rect 36636 12588 36688 12640
rect 45008 12656 45060 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 28540 12427 28592 12436
rect 28540 12393 28549 12427
rect 28549 12393 28583 12427
rect 28583 12393 28592 12427
rect 28540 12384 28592 12393
rect 29000 12384 29052 12436
rect 30012 12384 30064 12436
rect 30196 12427 30248 12436
rect 30196 12393 30205 12427
rect 30205 12393 30239 12427
rect 30239 12393 30248 12427
rect 30196 12384 30248 12393
rect 32588 12427 32640 12436
rect 32588 12393 32597 12427
rect 32597 12393 32631 12427
rect 32631 12393 32640 12427
rect 32588 12384 32640 12393
rect 32772 12384 32824 12436
rect 24860 12248 24912 12300
rect 27252 12248 27304 12300
rect 27896 12291 27948 12300
rect 27896 12257 27905 12291
rect 27905 12257 27939 12291
rect 27939 12257 27948 12291
rect 27896 12248 27948 12257
rect 29092 12248 29144 12300
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 25688 12180 25740 12232
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 27712 12223 27764 12232
rect 27712 12189 27721 12223
rect 27721 12189 27755 12223
rect 27755 12189 27764 12223
rect 27712 12180 27764 12189
rect 28356 12180 28408 12232
rect 29000 12180 29052 12232
rect 27436 12112 27488 12164
rect 32680 12316 32732 12368
rect 32036 12291 32088 12300
rect 30656 12180 30708 12232
rect 32036 12257 32045 12291
rect 32045 12257 32079 12291
rect 32079 12257 32088 12291
rect 32036 12248 32088 12257
rect 33140 12316 33192 12368
rect 35348 12316 35400 12368
rect 30380 12112 30432 12164
rect 31208 12189 31217 12210
rect 31217 12189 31251 12210
rect 31251 12189 31260 12210
rect 31208 12158 31260 12189
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 31484 12180 31536 12232
rect 33508 12248 33560 12300
rect 34428 12248 34480 12300
rect 34796 12248 34848 12300
rect 35532 12316 35584 12368
rect 36728 12384 36780 12436
rect 40776 12384 40828 12436
rect 41880 12384 41932 12436
rect 39120 12316 39172 12368
rect 32772 12223 32824 12232
rect 32772 12189 32781 12223
rect 32781 12189 32815 12223
rect 32815 12189 32824 12223
rect 32772 12180 32824 12189
rect 33048 12223 33100 12232
rect 33048 12189 33057 12223
rect 33057 12189 33091 12223
rect 33091 12189 33100 12223
rect 33048 12180 33100 12189
rect 33600 12180 33652 12232
rect 33876 12223 33928 12232
rect 33876 12189 33885 12223
rect 33885 12189 33919 12223
rect 33919 12189 33928 12223
rect 33876 12180 33928 12189
rect 34336 12180 34388 12232
rect 34612 12180 34664 12232
rect 36636 12248 36688 12300
rect 25504 12044 25556 12096
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 27528 12044 27580 12096
rect 30932 12044 30984 12096
rect 33508 12112 33560 12164
rect 39212 12180 39264 12232
rect 31484 12044 31536 12096
rect 32036 12044 32088 12096
rect 34244 12044 34296 12096
rect 34428 12044 34480 12096
rect 35808 12087 35860 12096
rect 35808 12053 35817 12087
rect 35817 12053 35851 12087
rect 35851 12053 35860 12087
rect 35808 12044 35860 12053
rect 36544 12087 36596 12096
rect 36544 12053 36553 12087
rect 36553 12053 36587 12087
rect 36587 12053 36596 12087
rect 36544 12044 36596 12053
rect 37188 12044 37240 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 25688 11883 25740 11892
rect 25688 11849 25697 11883
rect 25697 11849 25731 11883
rect 25731 11849 25740 11883
rect 25688 11840 25740 11849
rect 26148 11883 26200 11892
rect 26148 11849 26157 11883
rect 26157 11849 26191 11883
rect 26191 11849 26200 11883
rect 26148 11840 26200 11849
rect 27344 11840 27396 11892
rect 28816 11883 28868 11892
rect 28816 11849 28825 11883
rect 28825 11849 28859 11883
rect 28859 11849 28868 11883
rect 28816 11840 28868 11849
rect 30380 11840 30432 11892
rect 31208 11840 31260 11892
rect 31392 11840 31444 11892
rect 33140 11840 33192 11892
rect 33508 11883 33560 11892
rect 33508 11849 33517 11883
rect 33517 11849 33551 11883
rect 33551 11849 33560 11883
rect 33508 11840 33560 11849
rect 34244 11840 34296 11892
rect 18604 11704 18656 11756
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 27528 11747 27580 11756
rect 25228 11636 25280 11688
rect 26240 11636 26292 11688
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 27528 11713 27537 11747
rect 27537 11713 27571 11747
rect 27571 11713 27580 11747
rect 27528 11704 27580 11713
rect 29092 11772 29144 11824
rect 30012 11772 30064 11824
rect 33048 11772 33100 11824
rect 34428 11815 34480 11824
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 30472 11747 30524 11756
rect 30472 11713 30481 11747
rect 30481 11713 30515 11747
rect 30515 11713 30524 11747
rect 30472 11704 30524 11713
rect 31116 11704 31168 11756
rect 29184 11679 29236 11688
rect 29184 11645 29193 11679
rect 29193 11645 29227 11679
rect 29227 11645 29236 11679
rect 29184 11636 29236 11645
rect 31576 11747 31628 11756
rect 31576 11713 31585 11747
rect 31585 11713 31619 11747
rect 31619 11713 31628 11747
rect 31576 11704 31628 11713
rect 32772 11704 32824 11756
rect 34428 11781 34437 11815
rect 34437 11781 34471 11815
rect 34471 11781 34480 11815
rect 34428 11772 34480 11781
rect 34704 11772 34756 11824
rect 35532 11815 35584 11824
rect 35532 11781 35541 11815
rect 35541 11781 35575 11815
rect 35575 11781 35584 11815
rect 35532 11772 35584 11781
rect 35808 11772 35860 11824
rect 30656 11568 30708 11620
rect 32680 11636 32732 11688
rect 36268 11704 36320 11756
rect 36728 11747 36780 11756
rect 36728 11713 36737 11747
rect 36737 11713 36771 11747
rect 36771 11713 36780 11747
rect 36728 11704 36780 11713
rect 36912 11704 36964 11756
rect 38200 11747 38252 11756
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 40592 11772 40644 11824
rect 28448 11500 28500 11552
rect 34796 11543 34848 11552
rect 34796 11509 34805 11543
rect 34805 11509 34839 11543
rect 34839 11509 34848 11543
rect 34796 11500 34848 11509
rect 36544 11568 36596 11620
rect 39212 11704 39264 11756
rect 39304 11747 39356 11756
rect 39304 11713 39313 11747
rect 39313 11713 39347 11747
rect 39347 11713 39356 11747
rect 39304 11704 39356 11713
rect 35900 11543 35952 11552
rect 35900 11509 35909 11543
rect 35909 11509 35943 11543
rect 35943 11509 35952 11543
rect 35900 11500 35952 11509
rect 36360 11543 36412 11552
rect 36360 11509 36369 11543
rect 36369 11509 36403 11543
rect 36403 11509 36412 11543
rect 36360 11500 36412 11509
rect 39120 11500 39172 11552
rect 39764 11543 39816 11552
rect 39764 11509 39773 11543
rect 39773 11509 39807 11543
rect 39807 11509 39816 11543
rect 39764 11500 39816 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 24860 11296 24912 11348
rect 27436 11339 27488 11348
rect 26240 11271 26292 11280
rect 26240 11237 26249 11271
rect 26249 11237 26283 11271
rect 26283 11237 26292 11271
rect 26240 11228 26292 11237
rect 27436 11305 27445 11339
rect 27445 11305 27479 11339
rect 27479 11305 27488 11339
rect 27436 11296 27488 11305
rect 29276 11296 29328 11348
rect 30564 11296 30616 11348
rect 33232 11296 33284 11348
rect 33876 11296 33928 11348
rect 35532 11296 35584 11348
rect 29000 11228 29052 11280
rect 36360 11228 36412 11280
rect 36728 11296 36780 11348
rect 37004 11296 37056 11348
rect 37740 11296 37792 11348
rect 38200 11296 38252 11348
rect 58164 11339 58216 11348
rect 58164 11305 58173 11339
rect 58173 11305 58207 11339
rect 58207 11305 58216 11339
rect 58164 11296 58216 11305
rect 39304 11228 39356 11280
rect 29184 11160 29236 11212
rect 32312 11160 32364 11212
rect 33232 11160 33284 11212
rect 33968 11160 34020 11212
rect 37004 11203 37056 11212
rect 37004 11169 37013 11203
rect 37013 11169 37047 11203
rect 37047 11169 37056 11203
rect 37004 11160 37056 11169
rect 37372 11160 37424 11212
rect 29736 11135 29788 11144
rect 28724 10956 28776 11008
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 33508 11092 33560 11144
rect 33048 11024 33100 11076
rect 33692 11135 33744 11144
rect 33692 11101 33701 11135
rect 33701 11101 33735 11135
rect 33735 11101 33744 11135
rect 33692 11092 33744 11101
rect 34428 11092 34480 11144
rect 35716 11135 35768 11144
rect 35716 11101 35725 11135
rect 35725 11101 35759 11135
rect 35759 11101 35768 11135
rect 35716 11092 35768 11101
rect 36452 11092 36504 11144
rect 36912 11092 36964 11144
rect 37280 11135 37332 11144
rect 37280 11101 37289 11135
rect 37289 11101 37323 11135
rect 37323 11101 37332 11135
rect 37280 11092 37332 11101
rect 33876 11067 33928 11076
rect 33876 11033 33885 11067
rect 33885 11033 33919 11067
rect 33919 11033 33928 11067
rect 33876 11024 33928 11033
rect 38568 11024 38620 11076
rect 58256 11067 58308 11076
rect 58256 11033 58265 11067
rect 58265 11033 58299 11067
rect 58299 11033 58308 11067
rect 58256 11024 58308 11033
rect 32496 10956 32548 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 32312 10795 32364 10804
rect 27712 10684 27764 10736
rect 28724 10684 28776 10736
rect 32312 10761 32321 10795
rect 32321 10761 32355 10795
rect 32355 10761 32364 10795
rect 32312 10752 32364 10761
rect 33692 10752 33744 10804
rect 37280 10752 37332 10804
rect 30012 10727 30064 10736
rect 30012 10693 30021 10727
rect 30021 10693 30055 10727
rect 30055 10693 30064 10727
rect 30012 10684 30064 10693
rect 31024 10684 31076 10736
rect 31300 10684 31352 10736
rect 34428 10684 34480 10736
rect 34704 10684 34756 10736
rect 27068 10616 27120 10668
rect 33048 10616 33100 10668
rect 33508 10659 33560 10668
rect 33508 10625 33517 10659
rect 33517 10625 33551 10659
rect 33551 10625 33560 10659
rect 33508 10616 33560 10625
rect 29092 10548 29144 10600
rect 34612 10659 34664 10668
rect 34612 10625 34621 10659
rect 34621 10625 34655 10659
rect 34655 10625 34664 10659
rect 35716 10684 35768 10736
rect 36268 10727 36320 10736
rect 36268 10693 36277 10727
rect 36277 10693 36311 10727
rect 36311 10693 36320 10727
rect 36268 10684 36320 10693
rect 36452 10727 36504 10736
rect 36452 10693 36461 10727
rect 36461 10693 36495 10727
rect 36495 10693 36504 10727
rect 36452 10684 36504 10693
rect 39764 10684 39816 10736
rect 34612 10616 34664 10625
rect 34704 10591 34756 10600
rect 34704 10557 34713 10591
rect 34713 10557 34747 10591
rect 34747 10557 34756 10591
rect 34704 10548 34756 10557
rect 33968 10480 34020 10532
rect 39120 10523 39172 10532
rect 39120 10489 39129 10523
rect 39129 10489 39163 10523
rect 39163 10489 39172 10523
rect 39120 10480 39172 10489
rect 26424 10455 26476 10464
rect 26424 10421 26433 10455
rect 26433 10421 26467 10455
rect 26467 10421 26476 10455
rect 26424 10412 26476 10421
rect 32496 10455 32548 10464
rect 32496 10421 32505 10455
rect 32505 10421 32539 10455
rect 32539 10421 32548 10455
rect 32496 10412 32548 10421
rect 33232 10412 33284 10464
rect 36084 10455 36136 10464
rect 36084 10421 36093 10455
rect 36093 10421 36127 10455
rect 36127 10421 36136 10455
rect 36084 10412 36136 10421
rect 38292 10412 38344 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 27068 10208 27120 10260
rect 29092 10251 29144 10260
rect 29092 10217 29101 10251
rect 29101 10217 29135 10251
rect 29135 10217 29144 10251
rect 29092 10208 29144 10217
rect 30288 10208 30340 10260
rect 32496 10208 32548 10260
rect 33232 10251 33284 10260
rect 33232 10217 33241 10251
rect 33241 10217 33275 10251
rect 33275 10217 33284 10251
rect 33232 10208 33284 10217
rect 33692 10208 33744 10260
rect 29920 10140 29972 10192
rect 34520 10140 34572 10192
rect 31024 10072 31076 10124
rect 36084 10115 36136 10124
rect 36084 10081 36093 10115
rect 36093 10081 36127 10115
rect 36127 10081 36136 10115
rect 36084 10072 36136 10081
rect 37464 10072 37516 10124
rect 39120 10072 39172 10124
rect 28908 10004 28960 10056
rect 29736 10004 29788 10056
rect 31300 10004 31352 10056
rect 33048 10004 33100 10056
rect 33968 10004 34020 10056
rect 37188 10047 37240 10056
rect 37188 10013 37197 10047
rect 37197 10013 37231 10047
rect 37231 10013 37240 10047
rect 37188 10004 37240 10013
rect 38292 10047 38344 10056
rect 38292 10013 38301 10047
rect 38301 10013 38335 10047
rect 38335 10013 38344 10047
rect 38292 10004 38344 10013
rect 38568 10047 38620 10056
rect 38568 10013 38577 10047
rect 38577 10013 38611 10047
rect 38611 10013 38620 10047
rect 38568 10004 38620 10013
rect 37740 9936 37792 9988
rect 38384 9936 38436 9988
rect 39764 10004 39816 10056
rect 27896 9911 27948 9920
rect 27896 9877 27905 9911
rect 27905 9877 27939 9911
rect 27939 9877 27948 9911
rect 27896 9868 27948 9877
rect 28724 9868 28776 9920
rect 33692 9911 33744 9920
rect 33692 9877 33701 9911
rect 33701 9877 33735 9911
rect 33735 9877 33744 9911
rect 33692 9868 33744 9877
rect 35716 9868 35768 9920
rect 37648 9868 37700 9920
rect 57520 9868 57572 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 28908 9707 28960 9716
rect 28908 9673 28917 9707
rect 28917 9673 28951 9707
rect 28951 9673 28960 9707
rect 28908 9664 28960 9673
rect 36912 9664 36964 9716
rect 28724 9596 28776 9648
rect 30380 9596 30432 9648
rect 31300 9596 31352 9648
rect 32496 9639 32548 9648
rect 32496 9605 32505 9639
rect 32505 9605 32539 9639
rect 32539 9605 32548 9639
rect 33048 9639 33100 9648
rect 32496 9596 32548 9605
rect 33048 9605 33057 9639
rect 33057 9605 33091 9639
rect 33091 9605 33100 9639
rect 38384 9664 38436 9716
rect 33048 9596 33100 9605
rect 27068 9528 27120 9580
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 33692 9571 33744 9580
rect 33692 9537 33701 9571
rect 33701 9537 33735 9571
rect 33735 9537 33744 9571
rect 33692 9528 33744 9537
rect 33876 9571 33928 9580
rect 33876 9537 33885 9571
rect 33885 9537 33919 9571
rect 33919 9537 33928 9571
rect 33876 9528 33928 9537
rect 34520 9528 34572 9580
rect 34796 9528 34848 9580
rect 35532 9571 35584 9580
rect 27436 9503 27488 9512
rect 27436 9469 27445 9503
rect 27445 9469 27479 9503
rect 27479 9469 27488 9503
rect 27436 9460 27488 9469
rect 30564 9503 30616 9512
rect 30564 9469 30573 9503
rect 30573 9469 30607 9503
rect 30607 9469 30616 9503
rect 30564 9460 30616 9469
rect 30932 9460 30984 9512
rect 31208 9460 31260 9512
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 35716 9571 35768 9580
rect 35716 9537 35725 9571
rect 35725 9537 35759 9571
rect 35759 9537 35768 9571
rect 35716 9528 35768 9537
rect 37280 9528 37332 9580
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 38476 9503 38528 9512
rect 38476 9469 38485 9503
rect 38485 9469 38519 9503
rect 38519 9469 38528 9503
rect 38476 9460 38528 9469
rect 39120 9460 39172 9512
rect 32956 9392 33008 9444
rect 37464 9435 37516 9444
rect 37464 9401 37473 9435
rect 37473 9401 37507 9435
rect 37507 9401 37516 9435
rect 37464 9392 37516 9401
rect 30012 9367 30064 9376
rect 30012 9333 30021 9367
rect 30021 9333 30055 9367
rect 30055 9333 30064 9367
rect 30012 9324 30064 9333
rect 31116 9367 31168 9376
rect 31116 9333 31125 9367
rect 31125 9333 31159 9367
rect 31159 9333 31168 9367
rect 31116 9324 31168 9333
rect 31392 9367 31444 9376
rect 31392 9333 31401 9367
rect 31401 9333 31435 9367
rect 31435 9333 31444 9367
rect 31392 9324 31444 9333
rect 34796 9324 34848 9376
rect 35624 9367 35676 9376
rect 35624 9333 35633 9367
rect 35633 9333 35667 9367
rect 35667 9333 35676 9367
rect 35624 9324 35676 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 27436 9120 27488 9172
rect 28172 9120 28224 9172
rect 28724 9120 28776 9172
rect 30564 9120 30616 9172
rect 31116 9120 31168 9172
rect 32956 9163 33008 9172
rect 32956 9129 32965 9163
rect 32965 9129 32999 9163
rect 32999 9129 33008 9163
rect 32956 9120 33008 9129
rect 30656 9052 30708 9104
rect 26424 8916 26476 8968
rect 27160 8916 27212 8968
rect 27896 8916 27948 8968
rect 30012 8959 30064 8968
rect 30012 8925 30021 8959
rect 30021 8925 30055 8959
rect 30055 8925 30064 8959
rect 30012 8916 30064 8925
rect 31024 8984 31076 9036
rect 31208 8916 31260 8968
rect 32772 8984 32824 9036
rect 32956 8984 33008 9036
rect 33692 8984 33744 9036
rect 33876 8959 33928 8968
rect 27344 8848 27396 8900
rect 31484 8848 31536 8900
rect 33876 8925 33885 8959
rect 33885 8925 33919 8959
rect 33919 8925 33928 8959
rect 33876 8916 33928 8925
rect 35716 8984 35768 9036
rect 34520 8916 34572 8968
rect 35532 8959 35584 8968
rect 35532 8925 35541 8959
rect 35541 8925 35575 8959
rect 35575 8925 35584 8959
rect 35532 8916 35584 8925
rect 37648 8959 37700 8968
rect 37648 8925 37657 8959
rect 37657 8925 37691 8959
rect 37691 8925 37700 8959
rect 37648 8916 37700 8925
rect 37832 8916 37884 8968
rect 33048 8848 33100 8900
rect 57704 8848 57756 8900
rect 30472 8823 30524 8832
rect 30472 8789 30481 8823
rect 30481 8789 30515 8823
rect 30515 8789 30524 8823
rect 30472 8780 30524 8789
rect 33876 8780 33928 8832
rect 36084 8780 36136 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 27068 8576 27120 8628
rect 30380 8576 30432 8628
rect 31392 8576 31444 8628
rect 34060 8576 34112 8628
rect 35624 8576 35676 8628
rect 30564 8508 30616 8560
rect 30472 8440 30524 8492
rect 31024 8440 31076 8492
rect 31208 8483 31260 8492
rect 31208 8449 31217 8483
rect 31217 8449 31251 8483
rect 31251 8449 31260 8483
rect 31208 8440 31260 8449
rect 31484 8440 31536 8492
rect 32864 8508 32916 8560
rect 37648 8508 37700 8560
rect 32956 8483 33008 8492
rect 32956 8449 32965 8483
rect 32965 8449 32999 8483
rect 32999 8449 33008 8483
rect 32956 8440 33008 8449
rect 27160 8372 27212 8424
rect 27344 8347 27396 8356
rect 27344 8313 27353 8347
rect 27353 8313 27387 8347
rect 27387 8313 27396 8347
rect 27344 8304 27396 8313
rect 30104 8372 30156 8424
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 34796 8440 34848 8492
rect 35900 8483 35952 8492
rect 35900 8449 35909 8483
rect 35909 8449 35943 8483
rect 35943 8449 35952 8483
rect 35900 8440 35952 8449
rect 36084 8483 36136 8492
rect 36084 8449 36093 8483
rect 36093 8449 36127 8483
rect 36127 8449 36136 8483
rect 36084 8440 36136 8449
rect 33968 8372 34020 8424
rect 30656 8304 30708 8356
rect 37832 8304 37884 8356
rect 33232 8236 33284 8288
rect 37556 8279 37608 8288
rect 37556 8245 37565 8279
rect 37565 8245 37599 8279
rect 37599 8245 37608 8279
rect 37556 8236 37608 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 28172 8075 28224 8084
rect 28172 8041 28181 8075
rect 28181 8041 28215 8075
rect 28215 8041 28224 8075
rect 28172 8032 28224 8041
rect 30656 8032 30708 8084
rect 33876 8032 33928 8084
rect 31392 8007 31444 8016
rect 31392 7973 31401 8007
rect 31401 7973 31435 8007
rect 31435 7973 31444 8007
rect 31392 7964 31444 7973
rect 31024 7939 31076 7948
rect 31024 7905 31033 7939
rect 31033 7905 31067 7939
rect 31067 7905 31076 7939
rect 31024 7896 31076 7905
rect 31208 7828 31260 7880
rect 33232 7871 33284 7880
rect 33232 7837 33241 7871
rect 33241 7837 33275 7871
rect 33275 7837 33284 7871
rect 33232 7828 33284 7837
rect 33784 7828 33836 7880
rect 37556 7828 37608 7880
rect 33140 7760 33192 7812
rect 33968 7803 34020 7812
rect 31392 7692 31444 7744
rect 33968 7769 33995 7803
rect 33995 7769 34020 7803
rect 33968 7760 34020 7769
rect 34060 7760 34112 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 33692 7395 33744 7404
rect 33692 7361 33701 7395
rect 33701 7361 33735 7395
rect 33735 7361 33744 7395
rect 33692 7352 33744 7361
rect 31208 7284 31260 7336
rect 33784 7327 33836 7336
rect 33784 7293 33793 7327
rect 33793 7293 33827 7327
rect 33827 7293 33836 7327
rect 33784 7284 33836 7293
rect 22284 7148 22336 7200
rect 32956 7148 33008 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 33692 6987 33744 6996
rect 33692 6953 33701 6987
rect 33701 6953 33735 6987
rect 33735 6953 33744 6987
rect 33692 6944 33744 6953
rect 24952 6876 25004 6928
rect 27712 6876 27764 6928
rect 33232 6876 33284 6928
rect 33140 6740 33192 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 57520 5899 57572 5908
rect 57520 5865 57529 5899
rect 57529 5865 57563 5899
rect 57563 5865 57572 5899
rect 57520 5856 57572 5865
rect 20444 5652 20496 5704
rect 57520 5652 57572 5704
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 58256 5559 58308 5568
rect 58256 5525 58265 5559
rect 58265 5525 58299 5559
rect 58299 5525 58308 5559
rect 58256 5516 58308 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 27344 2524 27396 2576
rect 5540 2388 5592 2440
rect 14648 2456 14700 2508
rect 17684 2499 17736 2508
rect 17684 2465 17693 2499
rect 17693 2465 17727 2499
rect 17727 2465 17736 2499
rect 17684 2456 17736 2465
rect 31668 2592 31720 2644
rect 37096 2592 37148 2644
rect 44088 2635 44140 2644
rect 44088 2601 44097 2635
rect 44097 2601 44131 2635
rect 44131 2601 44140 2635
rect 44088 2592 44140 2601
rect 44180 2592 44232 2644
rect 34428 2524 34480 2576
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 25412 2388 25464 2440
rect 22192 2320 22244 2372
rect 20 2252 72 2304
rect 10968 2252 11020 2304
rect 16120 2252 16172 2304
rect 21916 2252 21968 2304
rect 27068 2252 27120 2304
rect 27712 2388 27764 2440
rect 43996 2456 44048 2508
rect 32956 2431 33008 2440
rect 32956 2397 32965 2431
rect 32965 2397 32999 2431
rect 32999 2397 33008 2431
rect 32956 2388 33008 2397
rect 37096 2388 37148 2440
rect 43812 2388 43864 2440
rect 32864 2252 32916 2304
rect 38016 2252 38068 2304
rect 48964 2252 49016 2304
rect 55128 2252 55180 2304
rect 59912 2252 59964 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 2594 59200 2650 59800
rect 8390 59200 8446 59800
rect 13542 59200 13598 59800
rect 19338 59200 19394 59800
rect 24490 59200 24546 59800
rect 30286 59200 30342 59800
rect 35438 59200 35494 59800
rect 41234 59200 41290 59800
rect 46386 59200 46442 59800
rect 52182 59200 52238 59800
rect 57334 59200 57390 59800
rect 1674 57896 1730 57905
rect 1674 57831 1730 57840
rect 1688 57594 1716 57831
rect 1676 57588 1728 57594
rect 1676 57530 1728 57536
rect 2608 57526 2636 59200
rect 8404 57594 8432 59200
rect 13556 57594 13584 59200
rect 19352 57594 19380 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 24504 57594 24532 59200
rect 8392 57588 8444 57594
rect 8392 57530 8444 57536
rect 13544 57588 13596 57594
rect 13544 57530 13596 57536
rect 19340 57588 19392 57594
rect 19340 57530 19392 57536
rect 24492 57588 24544 57594
rect 24492 57530 24544 57536
rect 30300 57526 30328 59200
rect 35452 57594 35480 59200
rect 35440 57588 35492 57594
rect 41248 57576 41276 59200
rect 46400 57594 46428 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 52196 57594 52224 59200
rect 57348 57594 57376 59200
rect 41420 57588 41472 57594
rect 41248 57548 41420 57576
rect 35440 57530 35492 57536
rect 41420 57530 41472 57536
rect 46388 57588 46440 57594
rect 46388 57530 46440 57536
rect 52184 57588 52236 57594
rect 52184 57530 52236 57536
rect 57336 57588 57388 57594
rect 57336 57530 57388 57536
rect 2596 57520 2648 57526
rect 2596 57462 2648 57468
rect 30288 57520 30340 57526
rect 30288 57462 30340 57468
rect 1860 57452 1912 57458
rect 1860 57394 1912 57400
rect 1872 56710 1900 57394
rect 2608 57050 2636 57462
rect 9864 57452 9916 57458
rect 9864 57394 9916 57400
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 25320 57452 25372 57458
rect 25320 57394 25372 57400
rect 35532 57452 35584 57458
rect 35532 57394 35584 57400
rect 41328 57452 41380 57458
rect 41328 57394 41380 57400
rect 46480 57452 46532 57458
rect 46480 57394 46532 57400
rect 52276 57452 52328 57458
rect 52276 57394 52328 57400
rect 9876 57254 9904 57394
rect 2872 57248 2924 57254
rect 2872 57190 2924 57196
rect 9864 57248 9916 57254
rect 9864 57190 9916 57196
rect 2596 57044 2648 57050
rect 2596 56986 2648 56992
rect 1860 56704 1912 56710
rect 1860 56646 1912 56652
rect 1676 51808 1728 51814
rect 1674 51776 1676 51785
rect 1728 51776 1730 51785
rect 1674 51711 1730 51720
rect 1676 46368 1728 46374
rect 1674 46336 1676 46345
rect 1728 46336 1730 46345
rect 1674 46271 1730 46280
rect 1872 45830 1900 56646
rect 2136 52012 2188 52018
rect 2136 51954 2188 51960
rect 2148 51814 2176 51954
rect 2136 51808 2188 51814
rect 2136 51750 2188 51756
rect 1860 45824 1912 45830
rect 1860 45766 1912 45772
rect 1952 40520 2004 40526
rect 1952 40462 2004 40468
rect 1676 40384 1728 40390
rect 1676 40326 1728 40332
rect 1688 40225 1716 40326
rect 1674 40216 1730 40225
rect 1674 40151 1730 40160
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1688 34785 1716 34886
rect 1674 34776 1730 34785
rect 1674 34711 1730 34720
rect 1676 29028 1728 29034
rect 1676 28970 1728 28976
rect 1688 28665 1716 28970
rect 1674 28656 1730 28665
rect 1674 28591 1730 28600
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23225 1716 23462
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1964 21962 1992 40462
rect 2044 34944 2096 34950
rect 2044 34886 2096 34892
rect 2056 24750 2084 34886
rect 2148 27441 2176 51750
rect 2320 46572 2372 46578
rect 2320 46514 2372 46520
rect 2332 46374 2360 46514
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2134 27432 2190 27441
rect 2134 27367 2190 27376
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 1952 21956 2004 21962
rect 1952 21898 2004 21904
rect 1674 17096 1730 17105
rect 1674 17031 1676 17040
rect 1728 17031 1730 17040
rect 1676 17002 1728 17008
rect 2332 16998 2360 46310
rect 2884 27606 2912 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 9876 28082 9904 57190
rect 14292 35834 14320 57394
rect 25332 57254 25360 57394
rect 32404 57384 32456 57390
rect 32404 57326 32456 57332
rect 25320 57248 25372 57254
rect 25320 57190 25372 57196
rect 30564 57248 30616 57254
rect 30564 57190 30616 57196
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 25332 55214 25360 57190
rect 30576 56681 30604 57190
rect 30562 56672 30618 56681
rect 30562 56607 30618 56616
rect 25332 55186 25452 55214
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 22376 47456 22428 47462
rect 22376 47398 22428 47404
rect 23204 47456 23256 47462
rect 23204 47398 23256 47404
rect 24676 47456 24728 47462
rect 24676 47398 24728 47404
rect 21272 47116 21324 47122
rect 21272 47058 21324 47064
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 21284 46578 21312 47058
rect 22098 47016 22154 47025
rect 22098 46951 22100 46960
rect 22152 46951 22154 46960
rect 22100 46922 22152 46928
rect 22388 46578 22416 47398
rect 23020 47048 23072 47054
rect 23020 46990 23072 46996
rect 23032 46578 23060 46990
rect 21272 46572 21324 46578
rect 21272 46514 21324 46520
rect 21548 46572 21600 46578
rect 21548 46514 21600 46520
rect 22376 46572 22428 46578
rect 22376 46514 22428 46520
rect 23020 46572 23072 46578
rect 23020 46514 23072 46520
rect 20812 46368 20864 46374
rect 20812 46310 20864 46316
rect 20444 45824 20496 45830
rect 20444 45766 20496 45772
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 20456 44470 20484 45766
rect 20720 45484 20772 45490
rect 20720 45426 20772 45432
rect 20536 44736 20588 44742
rect 20536 44678 20588 44684
rect 20628 44736 20680 44742
rect 20628 44678 20680 44684
rect 20444 44464 20496 44470
rect 20442 44432 20444 44441
rect 20496 44432 20498 44441
rect 18696 44396 18748 44402
rect 20442 44367 20498 44376
rect 18696 44338 18748 44344
rect 18708 43790 18736 44338
rect 20548 44334 20576 44678
rect 19432 44328 19484 44334
rect 19432 44270 19484 44276
rect 20536 44328 20588 44334
rect 20536 44270 20588 44276
rect 19156 44192 19208 44198
rect 19156 44134 19208 44140
rect 18696 43784 18748 43790
rect 18696 43726 18748 43732
rect 18604 43648 18656 43654
rect 18604 43590 18656 43596
rect 18616 43382 18644 43590
rect 18604 43376 18656 43382
rect 18604 43318 18656 43324
rect 19168 43246 19196 44134
rect 19444 43858 19472 44270
rect 20536 43988 20588 43994
rect 20536 43930 20588 43936
rect 19432 43852 19484 43858
rect 19432 43794 19484 43800
rect 20352 43784 20404 43790
rect 20352 43726 20404 43732
rect 19340 43648 19392 43654
rect 19340 43590 19392 43596
rect 19156 43240 19208 43246
rect 19156 43182 19208 43188
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18340 40050 18368 40462
rect 18512 40384 18564 40390
rect 18512 40326 18564 40332
rect 17776 40044 17828 40050
rect 17776 39986 17828 39992
rect 17960 40044 18012 40050
rect 17960 39986 18012 39992
rect 18328 40044 18380 40050
rect 18328 39986 18380 39992
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 17316 39296 17368 39302
rect 17316 39238 17368 39244
rect 16592 38962 16620 39238
rect 16580 38956 16632 38962
rect 16580 38898 16632 38904
rect 17040 38956 17092 38962
rect 17040 38898 17092 38904
rect 17224 38956 17276 38962
rect 17224 38898 17276 38904
rect 17052 38758 17080 38898
rect 17132 38820 17184 38826
rect 17132 38762 17184 38768
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 17040 38752 17092 38758
rect 17144 38729 17172 38762
rect 17040 38694 17092 38700
rect 17130 38720 17186 38729
rect 16592 38418 16620 38694
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16224 38270 16436 38298
rect 17052 38282 17080 38694
rect 17130 38655 17186 38664
rect 17144 38554 17172 38655
rect 17132 38548 17184 38554
rect 17132 38490 17184 38496
rect 15568 37868 15620 37874
rect 15568 37810 15620 37816
rect 15580 37262 15608 37810
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 15384 37188 15436 37194
rect 15384 37130 15436 37136
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 15396 35766 15424 37130
rect 15580 36718 15608 37198
rect 16120 36780 16172 36786
rect 16120 36722 16172 36728
rect 15568 36712 15620 36718
rect 15568 36654 15620 36660
rect 16132 36650 16160 36722
rect 16120 36644 16172 36650
rect 16120 36586 16172 36592
rect 15568 36576 15620 36582
rect 15568 36518 15620 36524
rect 15580 35834 15608 36518
rect 16132 35834 16160 36586
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 16120 35828 16172 35834
rect 16120 35770 16172 35776
rect 15200 35760 15252 35766
rect 15200 35702 15252 35708
rect 15384 35760 15436 35766
rect 15384 35702 15436 35708
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 15016 35692 15068 35698
rect 15016 35634 15068 35640
rect 14108 35290 14136 35634
rect 14096 35284 14148 35290
rect 14096 35226 14148 35232
rect 14936 35018 14964 35634
rect 15028 35290 15056 35634
rect 15016 35284 15068 35290
rect 15068 35244 15148 35272
rect 15016 35226 15068 35232
rect 14924 35012 14976 35018
rect 14924 34954 14976 34960
rect 14936 34746 14964 34954
rect 14924 34740 14976 34746
rect 14924 34682 14976 34688
rect 15120 34542 15148 35244
rect 15212 34950 15240 35702
rect 15580 35086 15608 35770
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15764 35154 15792 35634
rect 15752 35148 15804 35154
rect 15752 35090 15804 35096
rect 15568 35080 15620 35086
rect 15568 35022 15620 35028
rect 15948 34950 15976 35634
rect 15200 34944 15252 34950
rect 15200 34886 15252 34892
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15212 34678 15240 34886
rect 15200 34672 15252 34678
rect 15200 34614 15252 34620
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 15304 33454 15332 33934
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15212 33046 15240 33390
rect 15200 33040 15252 33046
rect 15200 32982 15252 32988
rect 15396 32586 15424 34342
rect 15672 34202 15700 34886
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 16224 34066 16252 38270
rect 16408 38214 16436 38270
rect 17040 38276 17092 38282
rect 17040 38218 17092 38224
rect 16304 38208 16356 38214
rect 16304 38150 16356 38156
rect 16396 38208 16448 38214
rect 16396 38150 16448 38156
rect 16316 36854 16344 38150
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16396 37664 16448 37670
rect 16396 37606 16448 37612
rect 16408 37262 16436 37606
rect 16592 37330 16620 37810
rect 16580 37324 16632 37330
rect 16580 37266 16632 37272
rect 17144 37262 17172 38490
rect 17236 38350 17264 38898
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 17236 38010 17264 38286
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 17224 37664 17276 37670
rect 17328 37652 17356 39238
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17696 37738 17724 38286
rect 17788 38214 17816 39986
rect 17972 39098 18000 39986
rect 18524 39642 18552 40326
rect 18604 39840 18656 39846
rect 18604 39782 18656 39788
rect 18512 39636 18564 39642
rect 18512 39578 18564 39584
rect 18616 39370 18644 39782
rect 18708 39642 18736 40870
rect 18880 40452 18932 40458
rect 18880 40394 18932 40400
rect 18788 40384 18840 40390
rect 18788 40326 18840 40332
rect 18696 39636 18748 39642
rect 18696 39578 18748 39584
rect 18604 39364 18656 39370
rect 18604 39306 18656 39312
rect 18052 39296 18104 39302
rect 18052 39238 18104 39244
rect 17960 39092 18012 39098
rect 17960 39034 18012 39040
rect 17868 38752 17920 38758
rect 17868 38694 17920 38700
rect 17880 38486 17908 38694
rect 17868 38480 17920 38486
rect 17868 38422 17920 38428
rect 17868 38344 17920 38350
rect 17868 38286 17920 38292
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 17788 37942 17816 38150
rect 17776 37936 17828 37942
rect 17776 37878 17828 37884
rect 17684 37732 17736 37738
rect 17684 37674 17736 37680
rect 17276 37624 17356 37652
rect 17224 37606 17276 37612
rect 17236 37262 17264 37606
rect 17592 37324 17644 37330
rect 17592 37266 17644 37272
rect 16396 37256 16448 37262
rect 17132 37256 17184 37262
rect 16396 37198 16448 37204
rect 16486 37224 16542 37233
rect 17132 37198 17184 37204
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 16486 37159 16542 37168
rect 16500 37126 16528 37159
rect 16488 37120 16540 37126
rect 16488 37062 16540 37068
rect 17500 37120 17552 37126
rect 17500 37062 17552 37068
rect 16304 36848 16356 36854
rect 16304 36790 16356 36796
rect 17512 36786 17540 37062
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16224 33522 16252 34002
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 15660 33380 15712 33386
rect 15660 33322 15712 33328
rect 15672 32978 15700 33322
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15304 32558 15424 32586
rect 15200 32292 15252 32298
rect 15200 32234 15252 32240
rect 14648 31748 14700 31754
rect 14648 31690 14700 31696
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 2872 27600 2924 27606
rect 2872 27542 2924 27548
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2516 17270 2544 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 1674 11656 1730 11665
rect 1674 11591 1676 11600
rect 1728 11591 1730 11600
rect 1676 11562 1728 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1676 5568 1728 5574
rect 1674 5536 1676 5545
rect 1728 5536 1730 5545
rect 1674 5471 1730 5480
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 14660 2514 14688 31690
rect 15212 31346 15240 32234
rect 15304 31822 15332 32558
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 15384 32224 15436 32230
rect 15384 32166 15436 32172
rect 15396 31822 15424 32166
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15212 30938 15240 31282
rect 15304 31278 15332 31758
rect 15856 31482 15884 32302
rect 15844 31476 15896 31482
rect 15844 31418 15896 31424
rect 15948 31346 15976 33254
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16132 31346 16160 32710
rect 16672 31884 16724 31890
rect 16672 31826 16724 31832
rect 16684 31414 16712 31826
rect 16672 31408 16724 31414
rect 16672 31350 16724 31356
rect 15936 31340 15988 31346
rect 15936 31282 15988 31288
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 15948 30938 15976 31282
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 16132 30802 16160 31282
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16684 30734 16712 31350
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16868 17202 16896 36654
rect 17224 36644 17276 36650
rect 17224 36586 17276 36592
rect 17236 36174 17264 36586
rect 17512 36378 17540 36722
rect 17604 36378 17632 37266
rect 17880 37210 17908 38286
rect 17972 37874 18000 39034
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 17788 37182 17908 37210
rect 17788 37126 17816 37182
rect 17776 37120 17828 37126
rect 17776 37062 17828 37068
rect 17500 36372 17552 36378
rect 17500 36314 17552 36320
rect 17592 36372 17644 36378
rect 17592 36314 17644 36320
rect 17224 36168 17276 36174
rect 17224 36110 17276 36116
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 17052 35086 17080 35634
rect 17132 35624 17184 35630
rect 17132 35566 17184 35572
rect 17144 35086 17172 35566
rect 17040 35080 17092 35086
rect 17040 35022 17092 35028
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17408 34128 17460 34134
rect 17408 34070 17460 34076
rect 17420 32910 17448 34070
rect 17788 32910 17816 37062
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 17972 33522 18000 33798
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 18064 31958 18092 39238
rect 18708 39098 18736 39578
rect 18512 39092 18564 39098
rect 18512 39034 18564 39040
rect 18696 39092 18748 39098
rect 18696 39034 18748 39040
rect 18524 38554 18552 39034
rect 18602 38720 18658 38729
rect 18602 38655 18658 38664
rect 18616 38554 18644 38655
rect 18512 38548 18564 38554
rect 18512 38490 18564 38496
rect 18604 38548 18656 38554
rect 18604 38490 18656 38496
rect 18696 38276 18748 38282
rect 18696 38218 18748 38224
rect 18708 38010 18736 38218
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18800 36786 18828 40326
rect 18892 40050 18920 40394
rect 18880 40044 18932 40050
rect 18880 39986 18932 39992
rect 18892 37874 18920 39986
rect 19260 38418 19288 43046
rect 19352 41313 19380 43590
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19984 43308 20036 43314
rect 20260 43308 20312 43314
rect 20036 43268 20260 43296
rect 19984 43250 20036 43256
rect 20260 43250 20312 43256
rect 19432 43104 19484 43110
rect 19432 43046 19484 43052
rect 19338 41304 19394 41313
rect 19338 41239 19394 41248
rect 19340 41132 19392 41138
rect 19340 41074 19392 41080
rect 19352 40050 19380 41074
rect 19444 40594 19472 43046
rect 20272 42906 20300 43250
rect 20364 43178 20392 43726
rect 20444 43716 20496 43722
rect 20444 43658 20496 43664
rect 20352 43172 20404 43178
rect 20352 43114 20404 43120
rect 20260 42900 20312 42906
rect 20260 42842 20312 42848
rect 20352 42628 20404 42634
rect 20352 42570 20404 42576
rect 20260 42560 20312 42566
rect 20260 42502 20312 42508
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 20168 42288 20220 42294
rect 20168 42230 20220 42236
rect 20076 42016 20128 42022
rect 20076 41958 20128 41964
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19982 41168 20038 41177
rect 20088 41138 20116 41958
rect 19982 41103 20038 41112
rect 20076 41132 20128 41138
rect 19432 40588 19484 40594
rect 19432 40530 19484 40536
rect 19340 40044 19392 40050
rect 19340 39986 19392 39992
rect 19444 39914 19472 40530
rect 19996 40474 20024 41103
rect 20076 41074 20128 41080
rect 19996 40446 20116 40474
rect 19984 40384 20036 40390
rect 19984 40326 20036 40332
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19892 40180 19944 40186
rect 19996 40168 20024 40326
rect 19944 40140 20024 40168
rect 19892 40122 19944 40128
rect 19432 39908 19484 39914
rect 19432 39850 19484 39856
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19248 38412 19300 38418
rect 19248 38354 19300 38360
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 19800 37868 19852 37874
rect 19800 37810 19852 37816
rect 18892 37330 18920 37810
rect 19812 37466 19840 37810
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 18880 37324 18932 37330
rect 18880 37266 18932 37272
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19444 36786 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19616 36780 19668 36786
rect 19616 36722 19668 36728
rect 18800 36174 18828 36722
rect 19444 36310 19472 36722
rect 19628 36378 19656 36722
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 19432 36304 19484 36310
rect 19432 36246 19484 36252
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18788 36168 18840 36174
rect 18788 36110 18840 36116
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 18524 35494 18552 36110
rect 18512 35488 18564 35494
rect 18512 35430 18564 35436
rect 18236 35148 18288 35154
rect 18236 35090 18288 35096
rect 18248 34746 18276 35090
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 18800 34678 18828 36110
rect 19352 35086 19380 36110
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 19444 35494 19472 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19524 35692 19576 35698
rect 19524 35634 19576 35640
rect 19708 35692 19760 35698
rect 19708 35634 19760 35640
rect 19432 35488 19484 35494
rect 19432 35430 19484 35436
rect 19536 35290 19564 35634
rect 19524 35284 19576 35290
rect 19524 35226 19576 35232
rect 19432 35216 19484 35222
rect 19432 35158 19484 35164
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 18512 34672 18564 34678
rect 18512 34614 18564 34620
rect 18788 34672 18840 34678
rect 18788 34614 18840 34620
rect 18524 34134 18552 34614
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 18512 34128 18564 34134
rect 18512 34070 18564 34076
rect 18524 33998 18552 34070
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18604 33992 18656 33998
rect 18604 33934 18656 33940
rect 18340 33862 18368 33934
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 18340 32978 18368 33798
rect 18524 33522 18552 33934
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18420 33312 18472 33318
rect 18420 33254 18472 33260
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 18432 32434 18460 33254
rect 18616 32774 18644 33934
rect 19260 32842 19288 34478
rect 19444 34066 19472 35158
rect 19720 35154 19748 35634
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34060 19484 34066
rect 19432 34002 19484 34008
rect 19444 33658 19472 34002
rect 19996 33998 20024 38354
rect 20088 35698 20116 40446
rect 20180 40118 20208 42230
rect 20272 40730 20300 42502
rect 20364 41682 20392 42570
rect 20456 42226 20484 43658
rect 20444 42220 20496 42226
rect 20444 42162 20496 42168
rect 20352 41676 20404 41682
rect 20352 41618 20404 41624
rect 20260 40724 20312 40730
rect 20260 40666 20312 40672
rect 20168 40112 20220 40118
rect 20168 40054 20220 40060
rect 20364 39506 20392 41618
rect 20444 41472 20496 41478
rect 20444 41414 20496 41420
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20168 39432 20220 39438
rect 20168 39374 20220 39380
rect 20260 39432 20312 39438
rect 20260 39374 20312 39380
rect 20180 39098 20208 39374
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20180 36786 20208 37198
rect 20168 36780 20220 36786
rect 20168 36722 20220 36728
rect 20180 36174 20208 36722
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 20180 35630 20208 36110
rect 20168 35624 20220 35630
rect 20168 35566 20220 35572
rect 20076 35556 20128 35562
rect 20076 35498 20128 35504
rect 20088 34678 20116 35498
rect 20076 34672 20128 34678
rect 20076 34614 20128 34620
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 20272 33862 20300 39374
rect 20456 39098 20484 41414
rect 20444 39092 20496 39098
rect 20444 39034 20496 39040
rect 20444 38820 20496 38826
rect 20444 38762 20496 38768
rect 20456 38729 20484 38762
rect 20442 38720 20498 38729
rect 20442 38655 20498 38664
rect 20548 38350 20576 43930
rect 20640 43858 20668 44678
rect 20628 43852 20680 43858
rect 20628 43794 20680 43800
rect 20626 43752 20682 43761
rect 20626 43687 20628 43696
rect 20680 43687 20682 43696
rect 20628 43658 20680 43664
rect 20732 43330 20760 45426
rect 20640 43302 20760 43330
rect 20640 42770 20668 43302
rect 20718 42936 20774 42945
rect 20718 42871 20774 42880
rect 20628 42764 20680 42770
rect 20628 42706 20680 42712
rect 20640 42362 20668 42706
rect 20732 42702 20760 42871
rect 20720 42696 20772 42702
rect 20720 42638 20772 42644
rect 20628 42356 20680 42362
rect 20628 42298 20680 42304
rect 20720 42220 20772 42226
rect 20720 42162 20772 42168
rect 20626 41304 20682 41313
rect 20626 41239 20682 41248
rect 20640 41206 20668 41239
rect 20628 41200 20680 41206
rect 20628 41142 20680 41148
rect 20732 41070 20760 42162
rect 20720 41064 20772 41070
rect 20720 41006 20772 41012
rect 20628 40928 20680 40934
rect 20628 40870 20680 40876
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20548 38214 20576 38286
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 20352 36304 20404 36310
rect 20352 36246 20404 36252
rect 20364 35698 20392 36246
rect 20548 36174 20576 37062
rect 20640 36802 20668 40870
rect 20720 39296 20772 39302
rect 20720 39238 20772 39244
rect 20732 38894 20760 39238
rect 20824 39030 20852 46310
rect 21088 45824 21140 45830
rect 21088 45766 21140 45772
rect 20902 45520 20958 45529
rect 20902 45455 20904 45464
rect 20956 45455 20958 45464
rect 20904 45426 20956 45432
rect 21100 45422 21128 45766
rect 21456 45552 21508 45558
rect 21456 45494 21508 45500
rect 21364 45484 21416 45490
rect 21364 45426 21416 45432
rect 21088 45416 21140 45422
rect 21088 45358 21140 45364
rect 21100 44946 21128 45358
rect 21180 45280 21232 45286
rect 21180 45222 21232 45228
rect 21088 44940 21140 44946
rect 21088 44882 21140 44888
rect 20996 44872 21048 44878
rect 20996 44814 21048 44820
rect 21008 43314 21036 44814
rect 21100 44470 21128 44882
rect 21088 44464 21140 44470
rect 21088 44406 21140 44412
rect 21192 43314 21220 45222
rect 21376 44520 21404 45426
rect 21468 44985 21496 45494
rect 21454 44976 21510 44985
rect 21454 44911 21510 44920
rect 21468 44878 21496 44911
rect 21456 44872 21508 44878
rect 21456 44814 21508 44820
rect 21456 44532 21508 44538
rect 21376 44492 21456 44520
rect 21456 44474 21508 44480
rect 21362 43888 21418 43897
rect 21362 43823 21418 43832
rect 21376 43790 21404 43823
rect 21364 43784 21416 43790
rect 21364 43726 21416 43732
rect 20996 43308 21048 43314
rect 20996 43250 21048 43256
rect 21180 43308 21232 43314
rect 21180 43250 21232 43256
rect 20904 42764 20956 42770
rect 20904 42706 20956 42712
rect 20916 42294 20944 42706
rect 21008 42634 21036 43250
rect 21088 42696 21140 42702
rect 21088 42638 21140 42644
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 20904 42288 20956 42294
rect 20904 42230 20956 42236
rect 20904 41472 20956 41478
rect 20904 41414 20956 41420
rect 20916 40050 20944 41414
rect 21100 41138 21128 42638
rect 21272 42016 21324 42022
rect 21272 41958 21324 41964
rect 21180 41268 21232 41274
rect 21180 41210 21232 41216
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 21100 40474 21128 41074
rect 21192 40594 21220 41210
rect 21180 40588 21232 40594
rect 21180 40530 21232 40536
rect 21100 40446 21220 40474
rect 21192 40390 21220 40446
rect 21088 40384 21140 40390
rect 21088 40326 21140 40332
rect 21180 40384 21232 40390
rect 21180 40326 21232 40332
rect 20904 40044 20956 40050
rect 20904 39986 20956 39992
rect 20996 39840 21048 39846
rect 20996 39782 21048 39788
rect 20904 39568 20956 39574
rect 20904 39510 20956 39516
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 20720 38888 20772 38894
rect 20720 38830 20772 38836
rect 20732 38010 20760 38830
rect 20824 38554 20852 38966
rect 20812 38548 20864 38554
rect 20812 38490 20864 38496
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20916 37874 20944 39510
rect 20904 37868 20956 37874
rect 20904 37810 20956 37816
rect 21008 37466 21036 39782
rect 21100 38010 21128 40326
rect 21180 39432 21232 39438
rect 21180 39374 21232 39380
rect 21192 39030 21220 39374
rect 21180 39024 21232 39030
rect 21180 38966 21232 38972
rect 21180 38344 21232 38350
rect 21178 38312 21180 38321
rect 21232 38312 21234 38321
rect 21178 38247 21234 38256
rect 21088 38004 21140 38010
rect 21088 37946 21140 37952
rect 21100 37466 21128 37946
rect 21284 37874 21312 41958
rect 21376 41002 21404 43726
rect 21468 42702 21496 44474
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 21468 41818 21496 42638
rect 21456 41812 21508 41818
rect 21456 41754 21508 41760
rect 21560 41750 21588 46514
rect 22100 46368 22152 46374
rect 22100 46310 22152 46316
rect 22112 44810 22140 46310
rect 22388 46102 22416 46514
rect 22376 46096 22428 46102
rect 22376 46038 22428 46044
rect 23216 45966 23244 47398
rect 24688 46986 24716 47398
rect 25228 47184 25280 47190
rect 25228 47126 25280 47132
rect 24768 47048 24820 47054
rect 24768 46990 24820 46996
rect 25136 47048 25188 47054
rect 25136 46990 25188 46996
rect 24676 46980 24728 46986
rect 24676 46922 24728 46928
rect 23296 46912 23348 46918
rect 23296 46854 23348 46860
rect 22560 45960 22612 45966
rect 22560 45902 22612 45908
rect 23204 45960 23256 45966
rect 23204 45902 23256 45908
rect 22284 45892 22336 45898
rect 22284 45834 22336 45840
rect 22192 45484 22244 45490
rect 22296 45472 22324 45834
rect 22376 45824 22428 45830
rect 22376 45766 22428 45772
rect 22388 45626 22416 45766
rect 22572 45626 22600 45902
rect 22744 45824 22796 45830
rect 22742 45792 22744 45801
rect 22796 45792 22798 45801
rect 22742 45727 22798 45736
rect 22376 45620 22428 45626
rect 22376 45562 22428 45568
rect 22560 45620 22612 45626
rect 22560 45562 22612 45568
rect 22376 45484 22428 45490
rect 22296 45444 22376 45472
rect 22192 45426 22244 45432
rect 22376 45426 22428 45432
rect 22204 45082 22232 45426
rect 22192 45076 22244 45082
rect 22192 45018 22244 45024
rect 22388 45014 22416 45426
rect 22376 45008 22428 45014
rect 22376 44950 22428 44956
rect 22192 44940 22244 44946
rect 22192 44882 22244 44888
rect 22008 44804 22060 44810
rect 22008 44746 22060 44752
rect 22100 44804 22152 44810
rect 22100 44746 22152 44752
rect 22020 44402 22048 44746
rect 22204 44402 22232 44882
rect 22008 44396 22060 44402
rect 22008 44338 22060 44344
rect 22192 44396 22244 44402
rect 22192 44338 22244 44344
rect 21732 44328 21784 44334
rect 21732 44270 21784 44276
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 21744 43602 21772 44270
rect 22008 44260 22060 44266
rect 22008 44202 22060 44208
rect 21916 43852 21968 43858
rect 21916 43794 21968 43800
rect 21822 43752 21878 43761
rect 21822 43687 21824 43696
rect 21876 43687 21878 43696
rect 21824 43658 21876 43664
rect 21744 43574 21864 43602
rect 21836 42838 21864 43574
rect 21824 42832 21876 42838
rect 21824 42774 21876 42780
rect 21732 42696 21784 42702
rect 21732 42638 21784 42644
rect 21640 42560 21692 42566
rect 21640 42502 21692 42508
rect 21548 41744 21600 41750
rect 21548 41686 21600 41692
rect 21456 41132 21508 41138
rect 21456 41074 21508 41080
rect 21364 40996 21416 41002
rect 21364 40938 21416 40944
rect 21362 39536 21418 39545
rect 21362 39471 21418 39480
rect 21376 39438 21404 39471
rect 21364 39432 21416 39438
rect 21364 39374 21416 39380
rect 21468 39302 21496 41074
rect 21560 41002 21588 41686
rect 21548 40996 21600 41002
rect 21548 40938 21600 40944
rect 21652 40882 21680 42502
rect 21744 42362 21772 42638
rect 21732 42356 21784 42362
rect 21732 42298 21784 42304
rect 21836 42294 21864 42774
rect 21928 42770 21956 43794
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 21824 42288 21876 42294
rect 21824 42230 21876 42236
rect 22020 42226 22048 44202
rect 22192 44192 22244 44198
rect 22192 44134 22244 44140
rect 22204 43994 22232 44134
rect 22192 43988 22244 43994
rect 22192 43930 22244 43936
rect 22296 43382 22324 44270
rect 22388 43722 22416 44950
rect 22468 44872 22520 44878
rect 22466 44840 22468 44849
rect 22520 44840 22522 44849
rect 22466 44775 22522 44784
rect 22468 44736 22520 44742
rect 22468 44678 22520 44684
rect 22376 43716 22428 43722
rect 22376 43658 22428 43664
rect 22100 43376 22152 43382
rect 22100 43318 22152 43324
rect 22284 43376 22336 43382
rect 22284 43318 22336 43324
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 21916 42084 21968 42090
rect 21916 42026 21968 42032
rect 21824 42016 21876 42022
rect 21824 41958 21876 41964
rect 21836 41070 21864 41958
rect 21928 41614 21956 42026
rect 21916 41608 21968 41614
rect 21916 41550 21968 41556
rect 21916 41472 21968 41478
rect 21916 41414 21968 41420
rect 21824 41064 21876 41070
rect 21824 41006 21876 41012
rect 21560 40854 21680 40882
rect 21560 39438 21588 40854
rect 21640 40724 21692 40730
rect 21640 40666 21692 40672
rect 21652 39574 21680 40666
rect 21732 40520 21784 40526
rect 21730 40488 21732 40497
rect 21784 40488 21786 40497
rect 21730 40423 21786 40432
rect 21732 40384 21784 40390
rect 21732 40326 21784 40332
rect 21640 39568 21692 39574
rect 21640 39510 21692 39516
rect 21548 39432 21600 39438
rect 21744 39409 21772 40326
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21836 39574 21864 39782
rect 21824 39568 21876 39574
rect 21824 39510 21876 39516
rect 21548 39374 21600 39380
rect 21730 39400 21786 39409
rect 21730 39335 21786 39344
rect 21456 39296 21508 39302
rect 21456 39238 21508 39244
rect 21468 38400 21496 39238
rect 21640 39024 21692 39030
rect 21640 38966 21692 38972
rect 21548 38412 21600 38418
rect 21468 38372 21548 38400
rect 21548 38354 21600 38360
rect 21272 37868 21324 37874
rect 21272 37810 21324 37816
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 21088 37460 21140 37466
rect 21088 37402 21140 37408
rect 21454 37360 21510 37369
rect 21454 37295 21510 37304
rect 21548 37324 21600 37330
rect 21364 37256 21416 37262
rect 21364 37198 21416 37204
rect 20640 36786 20760 36802
rect 20640 36780 20772 36786
rect 20640 36774 20720 36780
rect 20720 36722 20772 36728
rect 20628 36644 20680 36650
rect 20628 36586 20680 36592
rect 20640 36242 20668 36586
rect 20732 36310 20760 36722
rect 20996 36576 21048 36582
rect 20996 36518 21048 36524
rect 20720 36304 20772 36310
rect 20720 36246 20772 36252
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20548 35698 20576 36110
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20364 35154 20392 35634
rect 20352 35148 20404 35154
rect 20352 35090 20404 35096
rect 20548 35086 20576 35634
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20364 34202 20392 34342
rect 20352 34196 20404 34202
rect 20352 34138 20404 34144
rect 20536 34060 20588 34066
rect 20536 34002 20588 34008
rect 20260 33856 20312 33862
rect 20260 33798 20312 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 20272 33522 20300 33798
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20456 33046 20484 33254
rect 20444 33040 20496 33046
rect 20444 32982 20496 32988
rect 19248 32836 19300 32842
rect 19248 32778 19300 32784
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 19260 32570 19288 32778
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 20456 32434 20484 32982
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 18248 32026 18276 32302
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17696 31278 17724 31826
rect 18064 31822 18092 31894
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 18248 31346 18276 31962
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18432 31278 18460 32370
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 18616 31890 18644 32166
rect 19996 31890 20024 32166
rect 18604 31884 18656 31890
rect 18604 31826 18656 31832
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 20444 31884 20496 31890
rect 20444 31826 20496 31832
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 29238 16988 31078
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17972 30394 18000 30738
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 18524 30258 18552 31622
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 18880 31204 18932 31210
rect 18880 31146 18932 31152
rect 18892 30734 18920 31146
rect 20456 30938 20484 31826
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 20168 30728 20220 30734
rect 20168 30670 20220 30676
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 30258 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 16948 29232 17000 29238
rect 16948 29174 17000 29180
rect 16960 28694 16988 29174
rect 18064 29102 18092 30194
rect 18524 29782 18552 30194
rect 18512 29776 18564 29782
rect 18512 29718 18564 29724
rect 18524 29238 18552 29718
rect 19444 29646 19472 30194
rect 20180 30122 20208 30670
rect 20168 30116 20220 30122
rect 20168 30058 20220 30064
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18052 29096 18104 29102
rect 18052 29038 18104 29044
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 17868 28960 17920 28966
rect 17868 28902 17920 28908
rect 16948 28688 17000 28694
rect 16948 28630 17000 28636
rect 17880 28490 17908 28902
rect 18892 28558 18920 28970
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 17868 28484 17920 28490
rect 17868 28426 17920 28432
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 18616 11762 18644 28358
rect 19260 28014 19288 28494
rect 19352 28150 19380 29446
rect 19444 29102 19472 29582
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19996 29170 20024 29446
rect 20088 29170 20116 29582
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 20272 29034 20300 30738
rect 20456 30394 20484 30874
rect 20548 30666 20576 34002
rect 20732 33522 20760 35974
rect 20904 35624 20956 35630
rect 20904 35566 20956 35572
rect 20916 35086 20944 35566
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20916 34746 20944 35022
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 21008 33522 21036 36518
rect 21376 36174 21404 37198
rect 21364 36168 21416 36174
rect 21364 36110 21416 36116
rect 21468 35766 21496 37295
rect 21652 37312 21680 38966
rect 21744 37806 21772 39335
rect 21928 39114 21956 41414
rect 22020 39488 22048 42162
rect 22112 40186 22140 43318
rect 22388 43228 22416 43658
rect 22480 43314 22508 44678
rect 22572 43654 22600 45562
rect 22652 45280 22704 45286
rect 22652 45222 22704 45228
rect 22664 44305 22692 45222
rect 22756 44742 22784 45727
rect 23216 45286 23244 45902
rect 23308 45490 23336 46854
rect 24688 46578 24716 46922
rect 24676 46572 24728 46578
rect 24676 46514 24728 46520
rect 24780 46510 24808 46990
rect 25148 46646 25176 46990
rect 25136 46640 25188 46646
rect 25136 46582 25188 46588
rect 25240 46578 25268 47126
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25228 46572 25280 46578
rect 25228 46514 25280 46520
rect 24308 46504 24360 46510
rect 24308 46446 24360 46452
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 24032 46436 24084 46442
rect 24032 46378 24084 46384
rect 23664 46368 23716 46374
rect 23848 46368 23900 46374
rect 23716 46328 23796 46356
rect 23664 46310 23716 46316
rect 23572 45892 23624 45898
rect 23572 45834 23624 45840
rect 23480 45824 23532 45830
rect 23480 45766 23532 45772
rect 23296 45484 23348 45490
rect 23296 45426 23348 45432
rect 23308 45393 23336 45426
rect 23492 45422 23520 45766
rect 23480 45416 23532 45422
rect 23294 45384 23350 45393
rect 23480 45358 23532 45364
rect 23294 45319 23350 45328
rect 23112 45280 23164 45286
rect 23112 45222 23164 45228
rect 23204 45280 23256 45286
rect 23204 45222 23256 45228
rect 22836 44872 22888 44878
rect 22836 44814 22888 44820
rect 22744 44736 22796 44742
rect 22744 44678 22796 44684
rect 22848 44538 22876 44814
rect 23020 44736 23072 44742
rect 23020 44678 23072 44684
rect 22836 44532 22888 44538
rect 22836 44474 22888 44480
rect 22834 44432 22890 44441
rect 22834 44367 22836 44376
rect 22888 44367 22890 44376
rect 22836 44338 22888 44344
rect 22650 44296 22706 44305
rect 22650 44231 22706 44240
rect 22560 43648 22612 43654
rect 22560 43590 22612 43596
rect 22468 43308 22520 43314
rect 22468 43250 22520 43256
rect 22296 43200 22416 43228
rect 22192 43172 22244 43178
rect 22192 43114 22244 43120
rect 22204 42566 22232 43114
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22190 41848 22246 41857
rect 22190 41783 22246 41792
rect 22204 41750 22232 41783
rect 22192 41744 22244 41750
rect 22192 41686 22244 41692
rect 22192 41132 22244 41138
rect 22192 41074 22244 41080
rect 22100 40180 22152 40186
rect 22100 40122 22152 40128
rect 22204 40066 22232 41074
rect 22296 40526 22324 43200
rect 22480 42673 22508 43250
rect 22560 43104 22612 43110
rect 22560 43046 22612 43052
rect 22466 42664 22522 42673
rect 22466 42599 22522 42608
rect 22376 42084 22428 42090
rect 22376 42026 22428 42032
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 22296 40361 22324 40462
rect 22282 40352 22338 40361
rect 22282 40287 22338 40296
rect 22112 40050 22232 40066
rect 22100 40044 22232 40050
rect 22152 40038 22232 40044
rect 22284 40044 22336 40050
rect 22100 39986 22152 39992
rect 22284 39986 22336 39992
rect 22112 39914 22140 39986
rect 22190 39944 22246 39953
rect 22100 39908 22152 39914
rect 22190 39879 22246 39888
rect 22100 39850 22152 39856
rect 22100 39500 22152 39506
rect 22020 39460 22100 39488
rect 22100 39442 22152 39448
rect 22006 39264 22062 39273
rect 22006 39199 22062 39208
rect 21836 39086 21956 39114
rect 21732 37800 21784 37806
rect 21732 37742 21784 37748
rect 21652 37284 21772 37312
rect 21548 37266 21600 37272
rect 21560 37210 21588 37266
rect 21560 37182 21680 37210
rect 21744 37194 21772 37284
rect 21548 37120 21600 37126
rect 21548 37062 21600 37068
rect 21560 36582 21588 37062
rect 21548 36576 21600 36582
rect 21548 36518 21600 36524
rect 21560 36242 21588 36518
rect 21548 36236 21600 36242
rect 21548 36178 21600 36184
rect 21456 35760 21508 35766
rect 21456 35702 21508 35708
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 21100 34542 21128 34886
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21100 33658 21128 34342
rect 21468 34202 21496 35702
rect 21652 34950 21680 37182
rect 21732 37188 21784 37194
rect 21732 37130 21784 37136
rect 21836 36650 21864 39086
rect 22020 38962 22048 39199
rect 22112 39098 22140 39442
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22008 38956 22060 38962
rect 22008 38898 22060 38904
rect 22204 38826 22232 39879
rect 22192 38820 22244 38826
rect 22192 38762 22244 38768
rect 22008 38752 22060 38758
rect 22296 38729 22324 39986
rect 22388 39846 22416 42026
rect 22468 41608 22520 41614
rect 22468 41550 22520 41556
rect 22480 41449 22508 41550
rect 22466 41440 22522 41449
rect 22466 41375 22522 41384
rect 22466 41168 22522 41177
rect 22466 41103 22468 41112
rect 22520 41103 22522 41112
rect 22468 41074 22520 41080
rect 22376 39840 22428 39846
rect 22376 39782 22428 39788
rect 22468 39840 22520 39846
rect 22468 39782 22520 39788
rect 22388 39681 22416 39782
rect 22374 39672 22430 39681
rect 22374 39607 22430 39616
rect 22480 38962 22508 39782
rect 22468 38956 22520 38962
rect 22468 38898 22520 38904
rect 22008 38694 22060 38700
rect 22282 38720 22338 38729
rect 21916 38208 21968 38214
rect 21916 38150 21968 38156
rect 21928 37806 21956 38150
rect 21916 37800 21968 37806
rect 21916 37742 21968 37748
rect 21824 36644 21876 36650
rect 21824 36586 21876 36592
rect 21928 36106 21956 37742
rect 22020 37262 22048 38694
rect 22282 38655 22338 38664
rect 22296 38350 22324 38655
rect 22480 38570 22508 38898
rect 22388 38542 22508 38570
rect 22284 38344 22336 38350
rect 22284 38286 22336 38292
rect 22100 37936 22152 37942
rect 22100 37878 22152 37884
rect 22112 37398 22140 37878
rect 22284 37664 22336 37670
rect 22284 37606 22336 37612
rect 22100 37392 22152 37398
rect 22100 37334 22152 37340
rect 22192 37324 22244 37330
rect 22192 37266 22244 37272
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 22100 37120 22152 37126
rect 22100 37062 22152 37068
rect 22112 36854 22140 37062
rect 22204 36854 22232 37266
rect 22296 37262 22324 37606
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22100 36848 22152 36854
rect 22100 36790 22152 36796
rect 22192 36848 22244 36854
rect 22192 36790 22244 36796
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 22100 36032 22152 36038
rect 22100 35974 22152 35980
rect 21640 34944 21692 34950
rect 21640 34886 21692 34892
rect 21732 34944 21784 34950
rect 21732 34886 21784 34892
rect 21456 34196 21508 34202
rect 21456 34138 21508 34144
rect 21468 33930 21496 34138
rect 21652 33998 21680 34886
rect 21744 34610 21772 34886
rect 21732 34604 21784 34610
rect 21732 34546 21784 34552
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 21732 34468 21784 34474
rect 21732 34410 21784 34416
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21284 33114 21312 33798
rect 21640 33380 21692 33386
rect 21640 33322 21692 33328
rect 21272 33108 21324 33114
rect 21272 33050 21324 33056
rect 21284 32910 21312 33050
rect 21272 32904 21324 32910
rect 21272 32846 21324 32852
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 21364 32768 21416 32774
rect 21364 32710 21416 32716
rect 20640 32434 20668 32710
rect 20628 32428 20680 32434
rect 20628 32370 20680 32376
rect 21376 32230 21404 32710
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20548 30258 20576 30602
rect 20732 30326 20760 30602
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20916 30258 20944 31758
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 21008 30258 21036 30534
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 20824 29646 20852 30126
rect 20916 29714 20944 30194
rect 21008 29850 21036 30194
rect 21088 30048 21140 30054
rect 21088 29990 21140 29996
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20640 29034 20668 29514
rect 20824 29510 20852 29582
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20824 29170 20852 29446
rect 20916 29238 20944 29650
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 21008 29102 21036 29786
rect 21100 29782 21128 29990
rect 21088 29776 21140 29782
rect 21088 29718 21140 29724
rect 21376 29170 21404 32166
rect 21468 31822 21496 32166
rect 21456 31816 21508 31822
rect 21456 31758 21508 31764
rect 21652 31754 21680 33322
rect 21744 31822 21772 34410
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21640 31748 21692 31754
rect 21640 31690 21692 31696
rect 21652 31482 21680 31690
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21836 30734 21864 32710
rect 22020 31346 22048 34478
rect 22112 33930 22140 35974
rect 22296 35698 22324 37198
rect 22388 36242 22416 38542
rect 22468 38412 22520 38418
rect 22468 38354 22520 38360
rect 22480 37262 22508 38354
rect 22572 37874 22600 43046
rect 22652 42764 22704 42770
rect 22652 42706 22704 42712
rect 22664 39420 22692 42706
rect 22744 42696 22796 42702
rect 22742 42664 22744 42673
rect 22796 42664 22798 42673
rect 22742 42599 22798 42608
rect 22848 42566 22876 44338
rect 22836 42560 22888 42566
rect 22836 42502 22888 42508
rect 22744 42220 22796 42226
rect 22744 42162 22796 42168
rect 22756 41546 22784 42162
rect 23032 42090 23060 44678
rect 23020 42084 23072 42090
rect 23020 42026 23072 42032
rect 22744 41540 22796 41546
rect 22796 41500 22876 41528
rect 22744 41482 22796 41488
rect 22848 40458 22876 41500
rect 23124 41070 23152 45222
rect 23216 42770 23244 45222
rect 23388 44940 23440 44946
rect 23388 44882 23440 44888
rect 23296 43784 23348 43790
rect 23296 43726 23348 43732
rect 23204 42764 23256 42770
rect 23204 42706 23256 42712
rect 23308 41138 23336 43726
rect 23400 42702 23428 44882
rect 23480 44872 23532 44878
rect 23480 44814 23532 44820
rect 23492 44538 23520 44814
rect 23480 44532 23532 44538
rect 23480 44474 23532 44480
rect 23480 43648 23532 43654
rect 23480 43590 23532 43596
rect 23492 43314 23520 43590
rect 23480 43308 23532 43314
rect 23480 43250 23532 43256
rect 23584 43178 23612 45834
rect 23768 44402 23796 46328
rect 23848 46310 23900 46316
rect 23756 44396 23808 44402
rect 23756 44338 23808 44344
rect 23664 44328 23716 44334
rect 23664 44270 23716 44276
rect 23676 44198 23704 44270
rect 23664 44192 23716 44198
rect 23664 44134 23716 44140
rect 23860 43994 23888 46310
rect 24044 46034 24072 46378
rect 24032 46028 24084 46034
rect 24032 45970 24084 45976
rect 24320 45966 24348 46446
rect 24780 46374 24808 46446
rect 25136 46436 25188 46442
rect 25136 46378 25188 46384
rect 24768 46368 24820 46374
rect 24768 46310 24820 46316
rect 24584 46028 24636 46034
rect 24584 45970 24636 45976
rect 24308 45960 24360 45966
rect 24308 45902 24360 45908
rect 24032 45824 24084 45830
rect 24032 45766 24084 45772
rect 24044 44985 24072 45766
rect 24320 45422 24348 45902
rect 24308 45416 24360 45422
rect 24308 45358 24360 45364
rect 24400 45280 24452 45286
rect 24400 45222 24452 45228
rect 24030 44976 24086 44985
rect 24030 44911 24086 44920
rect 23940 44872 23992 44878
rect 23940 44814 23992 44820
rect 23952 44266 23980 44814
rect 23940 44260 23992 44266
rect 23940 44202 23992 44208
rect 23848 43988 23900 43994
rect 23848 43930 23900 43936
rect 23756 43308 23808 43314
rect 23756 43250 23808 43256
rect 23572 43172 23624 43178
rect 23572 43114 23624 43120
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 23480 42288 23532 42294
rect 23480 42230 23532 42236
rect 23388 41200 23440 41206
rect 23388 41142 23440 41148
rect 23296 41132 23348 41138
rect 23296 41074 23348 41080
rect 22928 41064 22980 41070
rect 22928 41006 22980 41012
rect 23112 41064 23164 41070
rect 23112 41006 23164 41012
rect 22940 40934 22968 41006
rect 22928 40928 22980 40934
rect 22928 40870 22980 40876
rect 22940 40526 22968 40870
rect 23308 40769 23336 41074
rect 23294 40760 23350 40769
rect 23124 40718 23294 40746
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22836 40452 22888 40458
rect 22836 40394 22888 40400
rect 23020 40384 23072 40390
rect 23020 40326 23072 40332
rect 22928 40044 22980 40050
rect 22928 39986 22980 39992
rect 22940 39438 22968 39986
rect 22744 39432 22796 39438
rect 22664 39392 22744 39420
rect 22744 39374 22796 39380
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22836 39296 22888 39302
rect 22836 39238 22888 39244
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22652 38208 22704 38214
rect 22652 38150 22704 38156
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22664 37806 22692 38150
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 22560 37664 22612 37670
rect 22560 37606 22612 37612
rect 22652 37664 22704 37670
rect 22652 37606 22704 37612
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22480 37126 22508 37198
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 22480 36786 22508 36858
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22376 36236 22428 36242
rect 22376 36178 22428 36184
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22572 34746 22600 37606
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 22100 33924 22152 33930
rect 22100 33866 22152 33872
rect 22112 32978 22140 33866
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 22204 33658 22232 33798
rect 22192 33652 22244 33658
rect 22192 33594 22244 33600
rect 22388 33522 22416 34614
rect 22664 34542 22692 37606
rect 22756 37244 22784 38490
rect 22848 38026 22876 39238
rect 22940 38214 22968 39374
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22848 37998 22968 38026
rect 22836 37256 22888 37262
rect 22756 37216 22836 37244
rect 22756 36922 22784 37216
rect 22836 37198 22888 37204
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 22848 36718 22876 37062
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22940 36242 22968 37998
rect 22928 36236 22980 36242
rect 22928 36178 22980 36184
rect 22834 35864 22890 35873
rect 22834 35799 22890 35808
rect 22848 35766 22876 35799
rect 22836 35760 22888 35766
rect 22836 35702 22888 35708
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22756 35290 22784 35634
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 22848 35086 22876 35702
rect 23032 35698 23060 40326
rect 23124 38418 23152 40718
rect 23294 40695 23350 40704
rect 23308 40635 23336 40695
rect 23400 40458 23428 41142
rect 23492 40934 23520 42230
rect 23480 40928 23532 40934
rect 23480 40870 23532 40876
rect 23388 40452 23440 40458
rect 23388 40394 23440 40400
rect 23400 40118 23428 40394
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 23492 40050 23520 40870
rect 23480 40044 23532 40050
rect 23480 39986 23532 39992
rect 23388 39976 23440 39982
rect 23388 39918 23440 39924
rect 23294 39808 23350 39817
rect 23294 39743 23350 39752
rect 23308 39030 23336 39743
rect 23400 39642 23428 39918
rect 23480 39908 23532 39914
rect 23480 39850 23532 39856
rect 23388 39636 23440 39642
rect 23388 39578 23440 39584
rect 23400 39438 23428 39578
rect 23388 39432 23440 39438
rect 23388 39374 23440 39380
rect 23388 39296 23440 39302
rect 23386 39264 23388 39273
rect 23440 39264 23442 39273
rect 23386 39199 23442 39208
rect 23400 39030 23428 39199
rect 23492 39137 23520 39850
rect 23478 39128 23534 39137
rect 23478 39063 23534 39072
rect 23296 39024 23348 39030
rect 23296 38966 23348 38972
rect 23388 39024 23440 39030
rect 23388 38966 23440 38972
rect 23492 38962 23520 39063
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23112 38412 23164 38418
rect 23164 38372 23244 38400
rect 23112 38354 23164 38360
rect 23112 38208 23164 38214
rect 23112 38150 23164 38156
rect 23124 37398 23152 38150
rect 23112 37392 23164 37398
rect 23112 37334 23164 37340
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 23124 35766 23152 37198
rect 23216 36310 23244 38372
rect 23296 38276 23348 38282
rect 23296 38218 23348 38224
rect 23308 37738 23336 38218
rect 23296 37732 23348 37738
rect 23296 37674 23348 37680
rect 23400 37330 23428 38830
rect 23584 38350 23612 43114
rect 23768 42702 23796 43250
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23756 42696 23808 42702
rect 23756 42638 23808 42644
rect 23676 42362 23704 42638
rect 23664 42356 23716 42362
rect 23664 42298 23716 42304
rect 23676 42226 23704 42298
rect 23664 42220 23716 42226
rect 23664 42162 23716 42168
rect 23676 41818 23704 42162
rect 23768 41818 23796 42638
rect 23860 42294 23888 43930
rect 23952 43314 23980 44202
rect 24044 43654 24072 44911
rect 24308 44532 24360 44538
rect 24308 44474 24360 44480
rect 24216 44396 24268 44402
rect 24216 44338 24268 44344
rect 24124 44192 24176 44198
rect 24124 44134 24176 44140
rect 24136 43722 24164 44134
rect 24124 43716 24176 43722
rect 24124 43658 24176 43664
rect 24032 43648 24084 43654
rect 24032 43590 24084 43596
rect 23940 43308 23992 43314
rect 23940 43250 23992 43256
rect 23848 42288 23900 42294
rect 23848 42230 23900 42236
rect 23952 42090 23980 43250
rect 23940 42084 23992 42090
rect 23940 42026 23992 42032
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23756 41812 23808 41818
rect 23756 41754 23808 41760
rect 23676 40526 23704 41754
rect 23940 41064 23992 41070
rect 23940 41006 23992 41012
rect 23952 40730 23980 41006
rect 23940 40724 23992 40730
rect 23940 40666 23992 40672
rect 24044 40610 24072 43590
rect 24136 43450 24164 43658
rect 24124 43444 24176 43450
rect 24124 43386 24176 43392
rect 24136 43314 24164 43386
rect 24228 43314 24256 44338
rect 24320 43994 24348 44474
rect 24412 44305 24440 45222
rect 24596 44402 24624 45970
rect 24952 45960 25004 45966
rect 24952 45902 25004 45908
rect 24860 45552 24912 45558
rect 24860 45494 24912 45500
rect 24676 45348 24728 45354
rect 24676 45290 24728 45296
rect 24688 44985 24716 45290
rect 24674 44976 24730 44985
rect 24872 44946 24900 45494
rect 24964 45422 24992 45902
rect 25148 45626 25176 46378
rect 25136 45620 25188 45626
rect 25136 45562 25188 45568
rect 24952 45416 25004 45422
rect 24952 45358 25004 45364
rect 24674 44911 24730 44920
rect 24860 44940 24912 44946
rect 24584 44396 24636 44402
rect 24584 44338 24636 44344
rect 24398 44296 24454 44305
rect 24398 44231 24454 44240
rect 24308 43988 24360 43994
rect 24308 43930 24360 43936
rect 24320 43790 24348 43930
rect 24308 43784 24360 43790
rect 24308 43726 24360 43732
rect 24124 43308 24176 43314
rect 24124 43250 24176 43256
rect 24216 43308 24268 43314
rect 24216 43250 24268 43256
rect 24124 42628 24176 42634
rect 24124 42570 24176 42576
rect 23860 40582 24072 40610
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23860 39370 23888 40582
rect 24032 40520 24084 40526
rect 24032 40462 24084 40468
rect 23940 39840 23992 39846
rect 23940 39782 23992 39788
rect 23848 39364 23900 39370
rect 23848 39306 23900 39312
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23662 38992 23718 39001
rect 23662 38927 23718 38936
rect 23676 38894 23704 38927
rect 23664 38888 23716 38894
rect 23664 38830 23716 38836
rect 23664 38752 23716 38758
rect 23664 38694 23716 38700
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23480 38004 23532 38010
rect 23480 37946 23532 37952
rect 23388 37324 23440 37330
rect 23388 37266 23440 37272
rect 23492 37194 23520 37946
rect 23676 37670 23704 38694
rect 23768 37874 23796 39238
rect 23756 37868 23808 37874
rect 23756 37810 23808 37816
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23676 37466 23704 37606
rect 23664 37460 23716 37466
rect 23664 37402 23716 37408
rect 23768 37330 23796 37810
rect 23860 37466 23888 39306
rect 23952 38729 23980 39782
rect 24044 39302 24072 40462
rect 24136 40050 24164 42570
rect 24228 42158 24256 43250
rect 24216 42152 24268 42158
rect 24216 42094 24268 42100
rect 24228 40526 24256 42094
rect 24320 41546 24348 43726
rect 24688 43314 24716 44911
rect 24860 44882 24912 44888
rect 24964 44826 24992 45358
rect 24872 44798 24992 44826
rect 24768 43376 24820 43382
rect 24768 43318 24820 43324
rect 24676 43308 24728 43314
rect 24676 43250 24728 43256
rect 24780 43110 24808 43318
rect 24768 43104 24820 43110
rect 24768 43046 24820 43052
rect 24676 42900 24728 42906
rect 24676 42842 24728 42848
rect 24688 42770 24716 42842
rect 24676 42764 24728 42770
rect 24676 42706 24728 42712
rect 24398 42528 24454 42537
rect 24398 42463 24454 42472
rect 24308 41540 24360 41546
rect 24308 41482 24360 41488
rect 24308 41064 24360 41070
rect 24308 41006 24360 41012
rect 24320 40730 24348 41006
rect 24308 40724 24360 40730
rect 24308 40666 24360 40672
rect 24216 40520 24268 40526
rect 24412 40497 24440 42463
rect 24490 42392 24546 42401
rect 24490 42327 24546 42336
rect 24504 42090 24532 42327
rect 24676 42220 24728 42226
rect 24676 42162 24728 42168
rect 24492 42084 24544 42090
rect 24492 42026 24544 42032
rect 24584 42016 24636 42022
rect 24584 41958 24636 41964
rect 24596 41682 24624 41958
rect 24584 41676 24636 41682
rect 24584 41618 24636 41624
rect 24492 41200 24544 41206
rect 24492 41142 24544 41148
rect 24216 40462 24268 40468
rect 24398 40488 24454 40497
rect 24398 40423 24454 40432
rect 24412 40338 24440 40423
rect 24228 40310 24440 40338
rect 24124 40044 24176 40050
rect 24124 39986 24176 39992
rect 24032 39296 24084 39302
rect 24032 39238 24084 39244
rect 24032 38956 24084 38962
rect 24228 38944 24256 40310
rect 24400 39976 24452 39982
rect 24504 39964 24532 41142
rect 24584 40384 24636 40390
rect 24584 40326 24636 40332
rect 24452 39936 24532 39964
rect 24400 39918 24452 39924
rect 24084 38916 24256 38944
rect 24032 38898 24084 38904
rect 24124 38752 24176 38758
rect 23938 38720 23994 38729
rect 24124 38694 24176 38700
rect 23938 38655 23994 38664
rect 24136 38486 24164 38694
rect 24124 38480 24176 38486
rect 24124 38422 24176 38428
rect 24032 38208 24084 38214
rect 24032 38150 24084 38156
rect 24044 37942 24072 38150
rect 24032 37936 24084 37942
rect 24032 37878 24084 37884
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23756 37324 23808 37330
rect 23756 37266 23808 37272
rect 23480 37188 23532 37194
rect 23480 37130 23532 37136
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23204 36304 23256 36310
rect 23204 36246 23256 36252
rect 23112 35760 23164 35766
rect 23112 35702 23164 35708
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 23032 35170 23060 35634
rect 23204 35488 23256 35494
rect 23204 35430 23256 35436
rect 22940 35154 23060 35170
rect 22928 35148 23060 35154
rect 22980 35142 23060 35148
rect 22928 35090 22980 35096
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 23020 34740 23072 34746
rect 23020 34682 23072 34688
rect 22652 34536 22704 34542
rect 22652 34478 22704 34484
rect 22744 34468 22796 34474
rect 22744 34410 22796 34416
rect 22756 33998 22784 34410
rect 23032 33998 23060 34682
rect 23216 34678 23244 35430
rect 23400 35018 23428 36722
rect 23388 35012 23440 35018
rect 23388 34954 23440 34960
rect 23676 34950 23704 37062
rect 24044 36786 24072 37878
rect 24124 37664 24176 37670
rect 24124 37606 24176 37612
rect 24216 37664 24268 37670
rect 24216 37606 24268 37612
rect 24136 37466 24164 37606
rect 24124 37460 24176 37466
rect 24124 37402 24176 37408
rect 24124 37120 24176 37126
rect 24124 37062 24176 37068
rect 24136 36922 24164 37062
rect 24124 36916 24176 36922
rect 24124 36858 24176 36864
rect 24228 36786 24256 37606
rect 24412 36854 24440 39918
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 24504 37874 24532 39034
rect 24596 38350 24624 40326
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 24688 37874 24716 42162
rect 24780 41274 24808 43046
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24780 40526 24808 41210
rect 24872 41138 24900 44798
rect 25148 44402 25176 45562
rect 25228 45348 25280 45354
rect 25332 45336 25360 46854
rect 25280 45308 25360 45336
rect 25228 45290 25280 45296
rect 25240 44946 25268 45290
rect 25228 44940 25280 44946
rect 25228 44882 25280 44888
rect 25136 44396 25188 44402
rect 25136 44338 25188 44344
rect 25240 44198 25268 44882
rect 25320 44736 25372 44742
rect 25320 44678 25372 44684
rect 25332 44305 25360 44678
rect 25318 44296 25374 44305
rect 25318 44231 25374 44240
rect 24952 44192 25004 44198
rect 24952 44134 25004 44140
rect 25228 44192 25280 44198
rect 25228 44134 25280 44140
rect 24860 41132 24912 41138
rect 24860 41074 24912 41080
rect 24768 40520 24820 40526
rect 24768 40462 24820 40468
rect 24964 40066 24992 44134
rect 25044 43648 25096 43654
rect 25044 43590 25096 43596
rect 25056 42702 25084 43590
rect 25044 42696 25096 42702
rect 25044 42638 25096 42644
rect 25056 42226 25084 42638
rect 25044 42220 25096 42226
rect 25044 42162 25096 42168
rect 25044 42084 25096 42090
rect 25044 42026 25096 42032
rect 25056 41614 25084 42026
rect 25044 41608 25096 41614
rect 25044 41550 25096 41556
rect 25136 41472 25188 41478
rect 25136 41414 25188 41420
rect 25148 41138 25176 41414
rect 25136 41132 25188 41138
rect 25136 41074 25188 41080
rect 24780 40050 24992 40066
rect 24768 40044 24992 40050
rect 24820 40038 24992 40044
rect 24768 39986 24820 39992
rect 25136 39976 25188 39982
rect 25240 39964 25268 44134
rect 25424 43353 25452 55186
rect 32416 48314 32444 57326
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 35544 57050 35572 57394
rect 35532 57044 35584 57050
rect 35532 56986 35584 56992
rect 35624 56704 35676 56710
rect 35624 56646 35676 56652
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 32416 48286 32628 48314
rect 29736 48000 29788 48006
rect 29736 47942 29788 47948
rect 25964 47796 26016 47802
rect 25964 47738 26016 47744
rect 25780 47592 25832 47598
rect 25780 47534 25832 47540
rect 25792 46986 25820 47534
rect 25976 47122 26004 47738
rect 27252 47728 27304 47734
rect 27252 47670 27304 47676
rect 26976 47184 27028 47190
rect 26976 47126 27028 47132
rect 25964 47116 26016 47122
rect 25964 47058 26016 47064
rect 25780 46980 25832 46986
rect 25780 46922 25832 46928
rect 25872 46368 25924 46374
rect 25872 46310 25924 46316
rect 25502 45792 25558 45801
rect 25502 45727 25558 45736
rect 25516 45490 25544 45727
rect 25504 45484 25556 45490
rect 25504 45426 25556 45432
rect 25688 45348 25740 45354
rect 25688 45290 25740 45296
rect 25594 44976 25650 44985
rect 25594 44911 25650 44920
rect 25608 44878 25636 44911
rect 25596 44872 25648 44878
rect 25596 44814 25648 44820
rect 25504 44804 25556 44810
rect 25504 44746 25556 44752
rect 25410 43344 25466 43353
rect 25516 43314 25544 44746
rect 25700 44742 25728 45290
rect 25780 45280 25832 45286
rect 25780 45222 25832 45228
rect 25792 44878 25820 45222
rect 25780 44872 25832 44878
rect 25780 44814 25832 44820
rect 25688 44736 25740 44742
rect 25688 44678 25740 44684
rect 25688 44532 25740 44538
rect 25688 44474 25740 44480
rect 25596 43784 25648 43790
rect 25596 43726 25648 43732
rect 25608 43450 25636 43726
rect 25596 43444 25648 43450
rect 25596 43386 25648 43392
rect 25700 43330 25728 44474
rect 25792 43790 25820 44814
rect 25780 43784 25832 43790
rect 25780 43726 25832 43732
rect 25700 43314 25820 43330
rect 25410 43279 25466 43288
rect 25504 43308 25556 43314
rect 25504 43250 25556 43256
rect 25700 43308 25832 43314
rect 25700 43302 25780 43308
rect 25516 42906 25544 43250
rect 25596 43172 25648 43178
rect 25596 43114 25648 43120
rect 25504 42900 25556 42906
rect 25504 42842 25556 42848
rect 25320 42016 25372 42022
rect 25320 41958 25372 41964
rect 25332 41614 25360 41958
rect 25320 41608 25372 41614
rect 25318 41576 25320 41585
rect 25372 41576 25374 41585
rect 25318 41511 25374 41520
rect 25320 40996 25372 41002
rect 25320 40938 25372 40944
rect 25188 39936 25268 39964
rect 25136 39918 25188 39924
rect 25044 39908 25096 39914
rect 25044 39850 25096 39856
rect 24952 39840 25004 39846
rect 24952 39782 25004 39788
rect 24858 39672 24914 39681
rect 24858 39607 24914 39616
rect 24872 39438 24900 39607
rect 24860 39432 24912 39438
rect 24860 39374 24912 39380
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 24676 37868 24728 37874
rect 24676 37810 24728 37816
rect 24688 37194 24716 37810
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24032 36780 24084 36786
rect 24032 36722 24084 36728
rect 24216 36780 24268 36786
rect 24216 36722 24268 36728
rect 24228 36106 24256 36722
rect 24780 36718 24808 37198
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 24780 36378 24808 36654
rect 24768 36372 24820 36378
rect 24768 36314 24820 36320
rect 24596 36242 24900 36258
rect 24584 36236 24900 36242
rect 24636 36230 24900 36236
rect 24584 36178 24636 36184
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 24216 36100 24268 36106
rect 24216 36042 24268 36048
rect 23756 35828 23808 35834
rect 23756 35770 23808 35776
rect 23664 34944 23716 34950
rect 23664 34886 23716 34892
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23032 33658 23060 33934
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 23216 33590 23244 34614
rect 23676 34610 23704 34886
rect 23480 34604 23532 34610
rect 23664 34604 23716 34610
rect 23532 34564 23612 34592
rect 23480 34546 23532 34552
rect 23584 34202 23612 34564
rect 23664 34546 23716 34552
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23480 34128 23532 34134
rect 23480 34070 23532 34076
rect 23204 33584 23256 33590
rect 23204 33526 23256 33532
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22848 32910 22876 33050
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22848 32434 22876 32846
rect 22940 32434 22968 33390
rect 23124 32774 23152 33458
rect 23388 33040 23440 33046
rect 23388 32982 23440 32988
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23020 32768 23072 32774
rect 23020 32710 23072 32716
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 23032 31822 23060 32710
rect 23308 32366 23336 32846
rect 23400 32774 23428 32982
rect 23388 32768 23440 32774
rect 23388 32710 23440 32716
rect 23492 32434 23520 34070
rect 23584 33522 23612 34138
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23676 33454 23704 34546
rect 23768 33930 23796 35770
rect 23860 35698 23888 36042
rect 24214 35864 24270 35873
rect 24504 35834 24532 36110
rect 24872 36038 24900 36230
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24214 35799 24270 35808
rect 24492 35828 24544 35834
rect 24228 35766 24256 35799
rect 24492 35770 24544 35776
rect 24216 35760 24268 35766
rect 24216 35702 24268 35708
rect 23848 35692 23900 35698
rect 23848 35634 23900 35640
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23756 33924 23808 33930
rect 23756 33866 23808 33872
rect 23768 33538 23796 33866
rect 23768 33522 23888 33538
rect 23768 33516 23900 33522
rect 23768 33510 23848 33516
rect 23848 33458 23900 33464
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23584 32366 23612 33254
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23296 32360 23348 32366
rect 23296 32302 23348 32308
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23676 32026 23704 32370
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 22284 31816 22336 31822
rect 22284 31758 22336 31764
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 22296 31346 22324 31758
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22284 30864 22336 30870
rect 22284 30806 22336 30812
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21744 29646 21772 29990
rect 21836 29714 21864 30670
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22112 29850 22140 30602
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 20996 29096 21048 29102
rect 20996 29038 21048 29044
rect 19616 29028 19668 29034
rect 19616 28970 19668 28976
rect 20260 29028 20312 29034
rect 20260 28970 20312 28976
rect 20628 29028 20680 29034
rect 20628 28970 20680 28976
rect 19432 28960 19484 28966
rect 19432 28902 19484 28908
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19352 27402 19380 28086
rect 19444 28014 19472 28902
rect 19628 28762 19656 28970
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 20628 28620 20680 28626
rect 20628 28562 20680 28568
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 20640 27470 20668 28562
rect 22296 28558 22324 30806
rect 22572 30734 22600 31078
rect 22756 30734 22784 31622
rect 22560 30728 22612 30734
rect 22744 30728 22796 30734
rect 22560 30670 22612 30676
rect 22664 30688 22744 30716
rect 22572 30258 22600 30670
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22468 29640 22520 29646
rect 22572 29628 22600 30194
rect 22664 30190 22692 30688
rect 22744 30670 22796 30676
rect 23952 30258 23980 35566
rect 24780 35086 24808 35974
rect 24964 35154 24992 39782
rect 25056 39556 25084 39850
rect 25136 39568 25188 39574
rect 25056 39528 25136 39556
rect 25136 39510 25188 39516
rect 25148 39273 25176 39510
rect 25240 39438 25268 39936
rect 25228 39432 25280 39438
rect 25228 39374 25280 39380
rect 25134 39264 25190 39273
rect 25134 39199 25190 39208
rect 25136 38888 25188 38894
rect 25136 38830 25188 38836
rect 25148 38486 25176 38830
rect 25136 38480 25188 38486
rect 25136 38422 25188 38428
rect 25226 38312 25282 38321
rect 25226 38247 25282 38256
rect 25136 38208 25188 38214
rect 25136 38150 25188 38156
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 25056 37262 25084 37606
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 25042 37088 25098 37097
rect 25042 37023 25098 37032
rect 25056 36174 25084 37023
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 24952 35148 25004 35154
rect 24952 35090 25004 35096
rect 24768 35080 24820 35086
rect 24768 35022 24820 35028
rect 25044 35080 25096 35086
rect 25148 35068 25176 38150
rect 25240 37738 25268 38247
rect 25228 37732 25280 37738
rect 25228 37674 25280 37680
rect 25096 35040 25176 35068
rect 25044 35022 25096 35028
rect 24584 34944 24636 34950
rect 24584 34886 24636 34892
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 24044 33590 24072 33798
rect 24596 33590 24624 34886
rect 25056 34746 25084 35022
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 24964 34066 24992 34682
rect 25228 34672 25280 34678
rect 25228 34614 25280 34620
rect 25240 34066 25268 34614
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24032 33584 24084 33590
rect 24032 33526 24084 33532
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 24688 32910 24716 33798
rect 24780 33590 24808 33866
rect 24952 33856 25004 33862
rect 24952 33798 25004 33804
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24964 33454 24992 33798
rect 25056 33590 25084 33798
rect 25044 33584 25096 33590
rect 25044 33526 25096 33532
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 24676 32904 24728 32910
rect 24676 32846 24728 32852
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24492 32768 24544 32774
rect 24492 32710 24544 32716
rect 24504 32366 24532 32710
rect 24688 32434 24716 32846
rect 24872 32502 24900 32846
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24492 32360 24544 32366
rect 24492 32302 24544 32308
rect 24504 31754 24532 32302
rect 24688 32026 24716 32370
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24676 32020 24728 32026
rect 24676 31962 24728 31968
rect 24780 31822 24808 32302
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24492 31748 24544 31754
rect 24492 31690 24544 31696
rect 24504 31482 24532 31690
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 24768 31340 24820 31346
rect 24872 31328 24900 32438
rect 25332 31822 25360 40938
rect 25516 40390 25544 42842
rect 25608 42838 25636 43114
rect 25596 42832 25648 42838
rect 25596 42774 25648 42780
rect 25700 42226 25728 43302
rect 25780 43250 25832 43256
rect 25780 42696 25832 42702
rect 25780 42638 25832 42644
rect 25792 42537 25820 42638
rect 25778 42528 25834 42537
rect 25778 42463 25834 42472
rect 25884 42226 25912 46310
rect 25976 44402 26004 47058
rect 26516 47048 26568 47054
rect 26516 46990 26568 46996
rect 26792 47048 26844 47054
rect 26792 46990 26844 46996
rect 26056 46912 26108 46918
rect 26056 46854 26108 46860
rect 26332 46912 26384 46918
rect 26332 46854 26384 46860
rect 26068 46578 26096 46854
rect 26056 46572 26108 46578
rect 26056 46514 26108 46520
rect 26068 44860 26096 46514
rect 26148 45960 26200 45966
rect 26148 45902 26200 45908
rect 26160 45490 26188 45902
rect 26148 45484 26200 45490
rect 26148 45426 26200 45432
rect 26160 45014 26188 45426
rect 26148 45008 26200 45014
rect 26148 44950 26200 44956
rect 26068 44832 26188 44860
rect 25964 44396 26016 44402
rect 25964 44338 26016 44344
rect 25964 43784 26016 43790
rect 25964 43726 26016 43732
rect 25976 43314 26004 43726
rect 25964 43308 26016 43314
rect 25964 43250 26016 43256
rect 26056 43104 26108 43110
rect 26056 43046 26108 43052
rect 26068 42702 26096 43046
rect 26056 42696 26108 42702
rect 26056 42638 26108 42644
rect 26068 42362 26096 42638
rect 26160 42566 26188 44832
rect 26240 43988 26292 43994
rect 26240 43930 26292 43936
rect 26252 43790 26280 43930
rect 26240 43784 26292 43790
rect 26240 43726 26292 43732
rect 26344 43382 26372 46854
rect 26528 46646 26556 46990
rect 26516 46640 26568 46646
rect 26516 46582 26568 46588
rect 26700 46572 26752 46578
rect 26700 46514 26752 46520
rect 26712 45966 26740 46514
rect 26804 46442 26832 46990
rect 26792 46436 26844 46442
rect 26792 46378 26844 46384
rect 26988 45966 27016 47126
rect 26700 45960 26752 45966
rect 26700 45902 26752 45908
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 26608 45892 26660 45898
rect 26608 45834 26660 45840
rect 26620 45490 26648 45834
rect 27264 45558 27292 47670
rect 28264 47660 28316 47666
rect 28264 47602 28316 47608
rect 28448 47660 28500 47666
rect 28448 47602 28500 47608
rect 27620 46912 27672 46918
rect 27620 46854 27672 46860
rect 27436 46368 27488 46374
rect 27436 46310 27488 46316
rect 27344 46096 27396 46102
rect 27344 46038 27396 46044
rect 27356 45830 27384 46038
rect 27448 46034 27476 46310
rect 27436 46028 27488 46034
rect 27436 45970 27488 45976
rect 27344 45824 27396 45830
rect 27344 45766 27396 45772
rect 27252 45552 27304 45558
rect 27252 45494 27304 45500
rect 26424 45484 26476 45490
rect 26424 45426 26476 45432
rect 26608 45484 26660 45490
rect 26608 45426 26660 45432
rect 26436 44946 26464 45426
rect 27448 45422 27476 45970
rect 27436 45416 27488 45422
rect 27436 45358 27488 45364
rect 26884 45348 26936 45354
rect 26884 45290 26936 45296
rect 26516 45280 26568 45286
rect 26516 45222 26568 45228
rect 26424 44940 26476 44946
rect 26424 44882 26476 44888
rect 26528 44305 26556 45222
rect 26896 45082 26924 45290
rect 26884 45076 26936 45082
rect 26884 45018 26936 45024
rect 27448 44810 27476 45358
rect 27528 45280 27580 45286
rect 27528 45222 27580 45228
rect 27540 44878 27568 45222
rect 27528 44872 27580 44878
rect 27526 44840 27528 44849
rect 27580 44840 27582 44849
rect 27436 44804 27488 44810
rect 27526 44775 27582 44784
rect 27436 44746 27488 44752
rect 26700 44396 26752 44402
rect 26700 44338 26752 44344
rect 26514 44296 26570 44305
rect 26514 44231 26570 44240
rect 26424 44192 26476 44198
rect 26424 44134 26476 44140
rect 26332 43376 26384 43382
rect 26332 43318 26384 43324
rect 26344 42838 26372 43318
rect 26332 42832 26384 42838
rect 26332 42774 26384 42780
rect 26344 42650 26372 42774
rect 26436 42770 26464 44134
rect 26516 43784 26568 43790
rect 26516 43726 26568 43732
rect 26528 43450 26556 43726
rect 26516 43444 26568 43450
rect 26516 43386 26568 43392
rect 26608 43172 26660 43178
rect 26608 43114 26660 43120
rect 26424 42764 26476 42770
rect 26424 42706 26476 42712
rect 26344 42622 26464 42650
rect 26148 42560 26200 42566
rect 26148 42502 26200 42508
rect 26056 42356 26108 42362
rect 26056 42298 26108 42304
rect 25688 42220 25740 42226
rect 25688 42162 25740 42168
rect 25872 42220 25924 42226
rect 25872 42162 25924 42168
rect 25884 42106 25912 42162
rect 25792 42078 25912 42106
rect 25688 42016 25740 42022
rect 25688 41958 25740 41964
rect 25596 41608 25648 41614
rect 25596 41550 25648 41556
rect 25608 41274 25636 41550
rect 25596 41268 25648 41274
rect 25596 41210 25648 41216
rect 25700 41138 25728 41958
rect 25688 41132 25740 41138
rect 25688 41074 25740 41080
rect 25688 40656 25740 40662
rect 25688 40598 25740 40604
rect 25504 40384 25556 40390
rect 25504 40326 25556 40332
rect 25412 39364 25464 39370
rect 25412 39306 25464 39312
rect 25424 38729 25452 39306
rect 25410 38720 25466 38729
rect 25410 38655 25466 38664
rect 25412 37936 25464 37942
rect 25412 37878 25464 37884
rect 25424 36922 25452 37878
rect 25516 37466 25544 40326
rect 25700 39982 25728 40598
rect 25792 40458 25820 42078
rect 25872 41608 25924 41614
rect 25872 41550 25924 41556
rect 25780 40452 25832 40458
rect 25780 40394 25832 40400
rect 25884 40050 25912 41550
rect 26068 41041 26096 42298
rect 26240 42220 26292 42226
rect 26240 42162 26292 42168
rect 26148 41540 26200 41546
rect 26148 41482 26200 41488
rect 26160 41206 26188 41482
rect 26252 41274 26280 42162
rect 26332 42152 26384 42158
rect 26332 42094 26384 42100
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 26148 41200 26200 41206
rect 26148 41142 26200 41148
rect 26054 41032 26110 41041
rect 26054 40967 26110 40976
rect 26240 40724 26292 40730
rect 26240 40666 26292 40672
rect 25964 40452 26016 40458
rect 25964 40394 26016 40400
rect 25872 40044 25924 40050
rect 25872 39986 25924 39992
rect 25688 39976 25740 39982
rect 25688 39918 25740 39924
rect 25700 39828 25728 39918
rect 25700 39800 25820 39828
rect 25688 39364 25740 39370
rect 25688 39306 25740 39312
rect 25596 38208 25648 38214
rect 25596 38150 25648 38156
rect 25504 37460 25556 37466
rect 25504 37402 25556 37408
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 25412 36780 25464 36786
rect 25412 36722 25464 36728
rect 25424 35630 25452 36722
rect 25608 36106 25636 38150
rect 25700 36378 25728 39306
rect 25792 37738 25820 39800
rect 25780 37732 25832 37738
rect 25780 37674 25832 37680
rect 25780 37460 25832 37466
rect 25780 37402 25832 37408
rect 25792 36666 25820 37402
rect 25884 37244 25912 39986
rect 25976 38486 26004 40394
rect 26252 40202 26280 40666
rect 26160 40174 26280 40202
rect 26056 39636 26108 39642
rect 26056 39578 26108 39584
rect 26068 39420 26096 39578
rect 26160 39438 26188 40174
rect 26240 40044 26292 40050
rect 26240 39986 26292 39992
rect 26148 39432 26200 39438
rect 26068 39392 26148 39420
rect 26148 39374 26200 39380
rect 26160 38826 26188 39374
rect 26148 38820 26200 38826
rect 26148 38762 26200 38768
rect 26056 38752 26108 38758
rect 26056 38694 26108 38700
rect 25964 38480 26016 38486
rect 25964 38422 26016 38428
rect 26068 38350 26096 38694
rect 26056 38344 26108 38350
rect 26056 38286 26108 38292
rect 26160 38214 26188 38762
rect 26252 38418 26280 39986
rect 26344 39098 26372 42094
rect 26436 40934 26464 42622
rect 26620 42022 26648 43114
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 26620 41478 26648 41958
rect 26516 41472 26568 41478
rect 26516 41414 26568 41420
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26528 41313 26556 41414
rect 26514 41304 26570 41313
rect 26514 41239 26570 41248
rect 26516 41200 26568 41206
rect 26516 41142 26568 41148
rect 26528 41041 26556 41142
rect 26514 41032 26570 41041
rect 26514 40967 26570 40976
rect 26424 40928 26476 40934
rect 26424 40870 26476 40876
rect 26528 40662 26556 40967
rect 26620 40730 26648 41414
rect 26608 40724 26660 40730
rect 26608 40666 26660 40672
rect 26516 40656 26568 40662
rect 26516 40598 26568 40604
rect 26712 39488 26740 44338
rect 27160 44328 27212 44334
rect 27528 44328 27580 44334
rect 27212 44288 27292 44316
rect 27160 44270 27212 44276
rect 27160 44192 27212 44198
rect 27160 44134 27212 44140
rect 27172 43790 27200 44134
rect 27160 43784 27212 43790
rect 27160 43726 27212 43732
rect 27068 43240 27120 43246
rect 27068 43182 27120 43188
rect 26976 42832 27028 42838
rect 26976 42774 27028 42780
rect 26792 42764 26844 42770
rect 26792 42706 26844 42712
rect 26436 39460 26740 39488
rect 26332 39092 26384 39098
rect 26332 39034 26384 39040
rect 26240 38412 26292 38418
rect 26240 38354 26292 38360
rect 26332 38344 26384 38350
rect 26332 38286 26384 38292
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 26146 38040 26202 38049
rect 26146 37975 26202 37984
rect 26160 37942 26188 37975
rect 26148 37936 26200 37942
rect 26148 37878 26200 37884
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 26160 37466 26188 37742
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 26252 37262 26280 37334
rect 25964 37256 26016 37262
rect 25884 37216 25964 37244
rect 26240 37256 26292 37262
rect 26016 37204 26188 37210
rect 25964 37198 26188 37204
rect 26240 37198 26292 37204
rect 25976 37182 26188 37198
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 25884 36854 25912 37062
rect 25872 36848 25924 36854
rect 25872 36790 25924 36796
rect 25792 36638 25912 36666
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25688 36372 25740 36378
rect 25688 36314 25740 36320
rect 25596 36100 25648 36106
rect 25596 36042 25648 36048
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25608 35562 25636 36042
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25700 35601 25728 35634
rect 25686 35592 25742 35601
rect 25596 35556 25648 35562
rect 25686 35527 25742 35536
rect 25596 35498 25648 35504
rect 25700 35018 25728 35527
rect 25688 35012 25740 35018
rect 25688 34954 25740 34960
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 25516 33504 25544 34478
rect 25608 33658 25636 34546
rect 25688 33924 25740 33930
rect 25688 33866 25740 33872
rect 25596 33652 25648 33658
rect 25596 33594 25648 33600
rect 25596 33516 25648 33522
rect 25516 33476 25596 33504
rect 25596 33458 25648 33464
rect 25504 32564 25556 32570
rect 25504 32506 25556 32512
rect 25516 32473 25544 32506
rect 25502 32464 25558 32473
rect 25502 32399 25558 32408
rect 25608 31822 25636 33458
rect 25700 32978 25728 33866
rect 25792 33862 25820 36518
rect 25884 35698 25912 36638
rect 26160 36582 26188 37182
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 26160 35766 26188 36518
rect 26148 35760 26200 35766
rect 26148 35702 26200 35708
rect 25872 35692 25924 35698
rect 25872 35634 25924 35640
rect 25884 35290 25912 35634
rect 26160 35494 26188 35702
rect 26344 35630 26372 38286
rect 26436 37194 26464 39460
rect 26514 39400 26570 39409
rect 26514 39335 26516 39344
rect 26568 39335 26570 39344
rect 26516 39306 26568 39312
rect 26804 39302 26832 42706
rect 26988 42090 27016 42774
rect 26976 42084 27028 42090
rect 26976 42026 27028 42032
rect 26884 42016 26936 42022
rect 26884 41958 26936 41964
rect 26896 39545 26924 41958
rect 26988 41818 27016 42026
rect 26976 41812 27028 41818
rect 26976 41754 27028 41760
rect 27080 41614 27108 43182
rect 27264 43178 27292 44288
rect 27528 44270 27580 44276
rect 27540 43382 27568 44270
rect 27528 43376 27580 43382
rect 27528 43318 27580 43324
rect 27160 43172 27212 43178
rect 27160 43114 27212 43120
rect 27252 43172 27304 43178
rect 27252 43114 27304 43120
rect 27172 42945 27200 43114
rect 27158 42936 27214 42945
rect 27158 42871 27214 42880
rect 27436 42764 27488 42770
rect 27436 42706 27488 42712
rect 27252 42696 27304 42702
rect 27252 42638 27304 42644
rect 27344 42696 27396 42702
rect 27344 42638 27396 42644
rect 27160 42560 27212 42566
rect 27160 42502 27212 42508
rect 27068 41608 27120 41614
rect 27068 41550 27120 41556
rect 26974 41440 27030 41449
rect 26974 41375 27030 41384
rect 26988 41274 27016 41375
rect 26976 41268 27028 41274
rect 26976 41210 27028 41216
rect 27172 41070 27200 42502
rect 27160 41064 27212 41070
rect 27158 41032 27160 41041
rect 27212 41032 27214 41041
rect 27158 40967 27214 40976
rect 27068 40928 27120 40934
rect 27264 40916 27292 42638
rect 27356 41614 27384 42638
rect 27448 41614 27476 42706
rect 27528 42560 27580 42566
rect 27528 42502 27580 42508
rect 27540 41993 27568 42502
rect 27526 41984 27582 41993
rect 27526 41919 27582 41928
rect 27632 41857 27660 46854
rect 27712 46708 27764 46714
rect 27712 46650 27764 46656
rect 27724 46578 27752 46650
rect 27896 46640 27948 46646
rect 27896 46582 27948 46588
rect 27712 46572 27764 46578
rect 27712 46514 27764 46520
rect 27724 45966 27752 46514
rect 27804 46028 27856 46034
rect 27804 45970 27856 45976
rect 27712 45960 27764 45966
rect 27712 45902 27764 45908
rect 27816 45354 27844 45970
rect 27908 45966 27936 46582
rect 28276 46442 28304 47602
rect 28264 46436 28316 46442
rect 28264 46378 28316 46384
rect 27988 46096 28040 46102
rect 27988 46038 28040 46044
rect 27896 45960 27948 45966
rect 27896 45902 27948 45908
rect 27804 45348 27856 45354
rect 27804 45290 27856 45296
rect 27804 44940 27856 44946
rect 27804 44882 27856 44888
rect 27816 43092 27844 44882
rect 27896 44872 27948 44878
rect 27896 44814 27948 44820
rect 27908 44402 27936 44814
rect 27896 44396 27948 44402
rect 27896 44338 27948 44344
rect 28000 43790 28028 46038
rect 28276 46034 28304 46378
rect 28460 46374 28488 47602
rect 29368 47592 29420 47598
rect 29368 47534 29420 47540
rect 28632 47184 28684 47190
rect 28632 47126 28684 47132
rect 28540 47048 28592 47054
rect 28540 46990 28592 46996
rect 28552 46578 28580 46990
rect 28540 46572 28592 46578
rect 28540 46514 28592 46520
rect 28448 46368 28500 46374
rect 28448 46310 28500 46316
rect 28540 46368 28592 46374
rect 28540 46310 28592 46316
rect 28264 46028 28316 46034
rect 28264 45970 28316 45976
rect 28080 45348 28132 45354
rect 28080 45290 28132 45296
rect 28092 44878 28120 45290
rect 28356 45280 28408 45286
rect 28356 45222 28408 45228
rect 28080 44872 28132 44878
rect 28080 44814 28132 44820
rect 28080 44192 28132 44198
rect 28080 44134 28132 44140
rect 27988 43784 28040 43790
rect 27988 43726 28040 43732
rect 27896 43104 27948 43110
rect 27816 43064 27896 43092
rect 27896 43046 27948 43052
rect 27804 42288 27856 42294
rect 27804 42230 27856 42236
rect 27618 41848 27674 41857
rect 27618 41783 27674 41792
rect 27632 41614 27660 41783
rect 27344 41608 27396 41614
rect 27342 41576 27344 41585
rect 27436 41608 27488 41614
rect 27396 41576 27398 41585
rect 27620 41608 27672 41614
rect 27488 41568 27568 41596
rect 27436 41550 27488 41556
rect 27342 41511 27398 41520
rect 27344 41200 27396 41206
rect 27344 41142 27396 41148
rect 27356 41070 27384 41142
rect 27344 41064 27396 41070
rect 27344 41006 27396 41012
rect 27264 40888 27384 40916
rect 27068 40870 27120 40876
rect 27080 40594 27108 40870
rect 27252 40724 27304 40730
rect 27252 40666 27304 40672
rect 27068 40588 27120 40594
rect 27068 40530 27120 40536
rect 27080 40050 27108 40530
rect 27160 40520 27212 40526
rect 27160 40462 27212 40468
rect 27172 40390 27200 40462
rect 27160 40384 27212 40390
rect 27160 40326 27212 40332
rect 27160 40112 27212 40118
rect 27264 40100 27292 40666
rect 27356 40594 27384 40888
rect 27344 40588 27396 40594
rect 27344 40530 27396 40536
rect 27356 40186 27384 40530
rect 27436 40384 27488 40390
rect 27436 40326 27488 40332
rect 27344 40180 27396 40186
rect 27344 40122 27396 40128
rect 27212 40072 27292 40100
rect 27160 40054 27212 40060
rect 27068 40044 27120 40050
rect 27068 39986 27120 39992
rect 26976 39976 27028 39982
rect 26976 39918 27028 39924
rect 26988 39681 27016 39918
rect 26974 39672 27030 39681
rect 26974 39607 27030 39616
rect 26882 39536 26938 39545
rect 26882 39471 26938 39480
rect 26988 39420 27016 39607
rect 27068 39500 27120 39506
rect 27068 39442 27120 39448
rect 26896 39392 27016 39420
rect 26700 39296 26752 39302
rect 26700 39238 26752 39244
rect 26792 39296 26844 39302
rect 26792 39238 26844 39244
rect 26514 39128 26570 39137
rect 26514 39063 26570 39072
rect 26424 37188 26476 37194
rect 26424 37130 26476 37136
rect 26436 36174 26464 37130
rect 26528 36786 26556 39063
rect 26712 39030 26740 39238
rect 26792 39092 26844 39098
rect 26792 39034 26844 39040
rect 26700 39024 26752 39030
rect 26700 38966 26752 38972
rect 26606 38856 26662 38865
rect 26606 38791 26662 38800
rect 26620 38758 26648 38791
rect 26608 38752 26660 38758
rect 26608 38694 26660 38700
rect 26608 38412 26660 38418
rect 26608 38354 26660 38360
rect 26620 36854 26648 38354
rect 26804 37262 26832 39034
rect 26896 38962 26924 39392
rect 26976 39296 27028 39302
rect 26976 39238 27028 39244
rect 26884 38956 26936 38962
rect 26884 38898 26936 38904
rect 26884 37460 26936 37466
rect 26884 37402 26936 37408
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26804 37126 26832 37198
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26608 36848 26660 36854
rect 26608 36790 26660 36796
rect 26516 36780 26568 36786
rect 26516 36722 26568 36728
rect 26792 36576 26844 36582
rect 26792 36518 26844 36524
rect 26516 36304 26568 36310
rect 26516 36246 26568 36252
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 25872 35284 25924 35290
rect 25872 35226 25924 35232
rect 26344 35018 26372 35566
rect 26528 35018 26556 36246
rect 26804 36174 26832 36518
rect 26896 36174 26924 37402
rect 26988 36786 27016 39238
rect 27080 38418 27108 39442
rect 27264 38894 27292 40072
rect 27448 39982 27476 40326
rect 27540 40100 27568 41568
rect 27620 41550 27672 41556
rect 27618 41304 27674 41313
rect 27816 41274 27844 42230
rect 27908 41682 27936 43046
rect 28000 42362 28028 43726
rect 27988 42356 28040 42362
rect 27988 42298 28040 42304
rect 28092 42226 28120 44134
rect 28264 43784 28316 43790
rect 28184 43744 28264 43772
rect 28184 42770 28212 43744
rect 28264 43726 28316 43732
rect 28264 43648 28316 43654
rect 28264 43590 28316 43596
rect 28276 43314 28304 43590
rect 28264 43308 28316 43314
rect 28264 43250 28316 43256
rect 28264 43172 28316 43178
rect 28264 43114 28316 43120
rect 28172 42764 28224 42770
rect 28172 42706 28224 42712
rect 28276 42650 28304 43114
rect 28184 42622 28304 42650
rect 28080 42220 28132 42226
rect 28080 42162 28132 42168
rect 27988 42016 28040 42022
rect 27988 41958 28040 41964
rect 27896 41676 27948 41682
rect 27896 41618 27948 41624
rect 27618 41239 27674 41248
rect 27804 41268 27856 41274
rect 27632 41138 27660 41239
rect 27804 41210 27856 41216
rect 27620 41132 27672 41138
rect 27620 41074 27672 41080
rect 27804 40928 27856 40934
rect 27804 40870 27856 40876
rect 27712 40520 27764 40526
rect 27712 40462 27764 40468
rect 27620 40112 27672 40118
rect 27540 40072 27620 40100
rect 27344 39976 27396 39982
rect 27344 39918 27396 39924
rect 27436 39976 27488 39982
rect 27540 39953 27568 40072
rect 27620 40054 27672 40060
rect 27620 39976 27672 39982
rect 27436 39918 27488 39924
rect 27526 39944 27582 39953
rect 27356 39642 27384 39918
rect 27620 39918 27672 39924
rect 27526 39879 27582 39888
rect 27436 39840 27488 39846
rect 27528 39840 27580 39846
rect 27436 39782 27488 39788
rect 27526 39808 27528 39817
rect 27580 39808 27582 39817
rect 27344 39636 27396 39642
rect 27344 39578 27396 39584
rect 27448 39556 27476 39782
rect 27526 39743 27582 39752
rect 27632 39642 27660 39918
rect 27724 39681 27752 40462
rect 27816 39982 27844 40870
rect 27804 39976 27856 39982
rect 27804 39918 27856 39924
rect 27802 39808 27858 39817
rect 27802 39743 27858 39752
rect 27710 39672 27766 39681
rect 27620 39636 27672 39642
rect 27710 39607 27766 39616
rect 27620 39578 27672 39584
rect 27448 39528 27568 39556
rect 27436 39092 27488 39098
rect 27436 39034 27488 39040
rect 27344 39024 27396 39030
rect 27344 38966 27396 38972
rect 27160 38888 27212 38894
rect 27160 38830 27212 38836
rect 27252 38888 27304 38894
rect 27252 38830 27304 38836
rect 27356 38842 27384 38966
rect 27448 38962 27476 39034
rect 27436 38956 27488 38962
rect 27436 38898 27488 38904
rect 27172 38758 27200 38830
rect 27356 38814 27476 38842
rect 27160 38752 27212 38758
rect 27160 38694 27212 38700
rect 27344 38752 27396 38758
rect 27344 38694 27396 38700
rect 27068 38412 27120 38418
rect 27068 38354 27120 38360
rect 27252 37868 27304 37874
rect 27252 37810 27304 37816
rect 27264 37194 27292 37810
rect 27252 37188 27304 37194
rect 27252 37130 27304 37136
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26792 36168 26844 36174
rect 26792 36110 26844 36116
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 26608 35556 26660 35562
rect 26608 35498 26660 35504
rect 26620 35086 26648 35498
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26332 35012 26384 35018
rect 26332 34954 26384 34960
rect 26516 35012 26568 35018
rect 26516 34954 26568 34960
rect 26056 34944 26108 34950
rect 26344 34921 26372 34954
rect 26056 34886 26108 34892
rect 26330 34912 26386 34921
rect 26068 34678 26096 34886
rect 26330 34847 26386 34856
rect 26804 34678 26832 36110
rect 26896 35698 26924 36110
rect 26988 36106 27016 36722
rect 27068 36304 27120 36310
rect 27068 36246 27120 36252
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 27080 35766 27108 36246
rect 27356 35766 27384 38694
rect 27448 38350 27476 38814
rect 27436 38344 27488 38350
rect 27436 38286 27488 38292
rect 27068 35760 27120 35766
rect 27068 35702 27120 35708
rect 27344 35760 27396 35766
rect 27344 35702 27396 35708
rect 26884 35692 26936 35698
rect 26884 35634 26936 35640
rect 27066 35592 27122 35601
rect 27066 35527 27122 35536
rect 27080 35086 27108 35527
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 26056 34672 26108 34678
rect 26056 34614 26108 34620
rect 26792 34672 26844 34678
rect 26792 34614 26844 34620
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 25780 33856 25832 33862
rect 25780 33798 25832 33804
rect 25688 32972 25740 32978
rect 25688 32914 25740 32920
rect 25700 32502 25728 32914
rect 25688 32496 25740 32502
rect 25688 32438 25740 32444
rect 25792 32434 25820 33798
rect 25872 32972 25924 32978
rect 25872 32914 25924 32920
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25688 32292 25740 32298
rect 25688 32234 25740 32240
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25596 31816 25648 31822
rect 25596 31758 25648 31764
rect 24820 31300 24900 31328
rect 24768 31282 24820 31288
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24308 30796 24360 30802
rect 24308 30738 24360 30744
rect 23940 30252 23992 30258
rect 23940 30194 23992 30200
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22664 29646 22692 30126
rect 23756 30116 23808 30122
rect 23756 30058 23808 30064
rect 22520 29600 22600 29628
rect 22652 29640 22704 29646
rect 22468 29582 22520 29588
rect 22652 29582 22704 29588
rect 23768 29170 23796 30058
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 24124 29504 24176 29510
rect 24124 29446 24176 29452
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23860 29034 23888 29446
rect 24136 29306 24164 29446
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 23848 29028 23900 29034
rect 23848 28970 23900 28976
rect 23572 28960 23624 28966
rect 23572 28902 23624 28908
rect 23584 28626 23612 28902
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 22284 28552 22336 28558
rect 22204 28500 22284 28506
rect 22204 28494 22336 28500
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20996 28484 21048 28490
rect 20996 28426 21048 28432
rect 22204 28478 22324 28494
rect 20916 28082 20944 28426
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 20916 27334 20944 28018
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 21008 27062 21036 28426
rect 22204 28150 22232 28478
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 21364 27872 21416 27878
rect 21364 27814 21416 27820
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 21376 26994 21404 27814
rect 22204 27538 22232 28086
rect 22296 28082 22324 28358
rect 22480 28150 22508 28494
rect 22468 28144 22520 28150
rect 22468 28086 22520 28092
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22192 27532 22244 27538
rect 22192 27474 22244 27480
rect 22480 27470 22508 28086
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20456 5710 20484 26862
rect 23400 26586 23428 26998
rect 23860 26586 23888 27270
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23848 23248 23900 23254
rect 23848 23190 23900 23196
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21744 22030 21772 22918
rect 22296 22030 22324 22986
rect 22848 22778 22876 23054
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22848 22098 22876 22714
rect 23584 22642 23612 23054
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22848 21486 22876 22034
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23308 21622 23336 21830
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 17682 2544 17738 2553
rect 14648 2508 14700 2514
rect 17682 2479 17684 2488
rect 14648 2450 14700 2456
rect 17736 2479 17738 2488
rect 17684 2450 17736 2456
rect 5540 2440 5592 2446
rect 5460 2388 5540 2394
rect 5460 2382 5592 2388
rect 5460 2366 5580 2382
rect 22204 2378 22232 21422
rect 23400 21146 23428 21898
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21554 23520 21830
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23584 20534 23612 22578
rect 23676 21690 23704 22918
rect 23860 22642 23888 23190
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23768 21690 23796 21898
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23768 20942 23796 21422
rect 23860 20942 23888 21490
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22848 19922 22876 20334
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23032 19854 23060 20402
rect 23768 20058 23796 20878
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 19310 23520 19790
rect 23676 19378 23704 19994
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23768 19378 23796 19790
rect 23860 19514 23888 20878
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18970 23520 19246
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23584 18290 23612 18770
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18290 23888 18566
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23952 17202 23980 21558
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23492 13938 23520 15302
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23400 13818 23428 13874
rect 23676 13818 23704 17138
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 14074 23796 14214
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23400 13790 23704 13818
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 13326 23428 13670
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23584 13190 23612 13790
rect 23768 13394 23796 14010
rect 23860 13870 23888 14010
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 24044 13802 24072 27406
rect 24228 26790 24256 30194
rect 24320 29102 24348 30738
rect 24596 30258 24624 31078
rect 24768 30864 24820 30870
rect 24674 30832 24730 30841
rect 24768 30806 24820 30812
rect 24674 30767 24730 30776
rect 24688 30734 24716 30767
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24780 30258 24808 30806
rect 25332 30734 25360 31758
rect 25700 30802 25728 32234
rect 25792 31958 25820 32370
rect 25780 31952 25832 31958
rect 25780 31894 25832 31900
rect 25884 31890 25912 32914
rect 25976 32774 26004 33934
rect 26436 33590 26464 34478
rect 26792 34468 26844 34474
rect 26792 34410 26844 34416
rect 26608 33992 26660 33998
rect 26608 33934 26660 33940
rect 26620 33658 26648 33934
rect 26608 33652 26660 33658
rect 26608 33594 26660 33600
rect 26424 33584 26476 33590
rect 26476 33532 26556 33538
rect 26424 33526 26556 33532
rect 26436 33510 26556 33526
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26056 33040 26108 33046
rect 26056 32982 26108 32988
rect 25964 32768 26016 32774
rect 25964 32710 26016 32716
rect 25976 32570 26004 32710
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 26068 32450 26096 32982
rect 26344 32910 26372 33254
rect 26528 33046 26556 33510
rect 26620 33114 26648 33594
rect 26700 33380 26752 33386
rect 26700 33322 26752 33328
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 26516 33040 26568 33046
rect 26516 32982 26568 32988
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26344 32450 26372 32506
rect 26068 32422 26372 32450
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 25884 31754 25912 31826
rect 26332 31816 26384 31822
rect 26252 31776 26332 31804
rect 25872 31748 25924 31754
rect 25872 31690 25924 31696
rect 25884 31346 25912 31690
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 26068 31346 26096 31622
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 25964 31272 26016 31278
rect 25964 31214 26016 31220
rect 25976 30938 26004 31214
rect 25964 30932 26016 30938
rect 25964 30874 26016 30880
rect 25688 30796 25740 30802
rect 25688 30738 25740 30744
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 26252 30433 26280 31776
rect 26332 31758 26384 31764
rect 26528 31686 26556 32982
rect 26620 32434 26648 33050
rect 26712 32978 26740 33322
rect 26804 33114 26832 34410
rect 27172 34066 27200 35430
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 27264 34610 27292 34886
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 27160 34060 27212 34066
rect 27160 34002 27212 34008
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26792 33108 26844 33114
rect 26792 33050 26844 33056
rect 26700 32972 26752 32978
rect 26700 32914 26752 32920
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 26332 30592 26384 30598
rect 26332 30534 26384 30540
rect 26238 30424 26294 30433
rect 26238 30359 26240 30368
rect 26292 30359 26294 30368
rect 26240 30330 26292 30336
rect 26344 30258 26372 30534
rect 26436 30394 26464 30670
rect 26528 30666 26556 31622
rect 26516 30660 26568 30666
rect 26516 30602 26568 30608
rect 26424 30388 26476 30394
rect 26424 30330 26476 30336
rect 26620 30258 26648 32370
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24768 30252 24820 30258
rect 24768 30194 24820 30200
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 24596 29646 24624 30194
rect 24780 29782 24808 30194
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 25056 29220 25084 29650
rect 25136 29232 25188 29238
rect 25056 29192 25136 29220
rect 24308 29096 24360 29102
rect 24308 29038 24360 29044
rect 25056 28558 25084 29192
rect 25136 29174 25188 29180
rect 25332 29170 25360 29990
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25976 29306 26004 29582
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 26240 29028 26292 29034
rect 26240 28970 26292 28976
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 25148 28490 25176 28902
rect 25596 28688 25648 28694
rect 25596 28630 25648 28636
rect 25136 28484 25188 28490
rect 25136 28426 25188 28432
rect 25148 28082 25176 28426
rect 25412 28416 25464 28422
rect 25412 28358 25464 28364
rect 25424 28082 25452 28358
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25148 27470 25176 28018
rect 25608 27878 25636 28630
rect 26252 28626 26280 28970
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25608 27470 25636 27814
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24596 27130 24624 27338
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24136 26042 24164 26318
rect 24228 26314 24256 26726
rect 24596 26450 24624 26862
rect 26804 26450 26832 33050
rect 26988 32230 27016 33934
rect 27172 33522 27200 34002
rect 27264 33658 27292 34546
rect 27540 34456 27568 39528
rect 27620 39432 27672 39438
rect 27620 39374 27672 39380
rect 27632 39137 27660 39374
rect 27816 39302 27844 39743
rect 27712 39296 27764 39302
rect 27712 39238 27764 39244
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27618 39128 27674 39137
rect 27618 39063 27620 39072
rect 27672 39063 27674 39072
rect 27620 39034 27672 39040
rect 27632 39003 27660 39034
rect 27724 38944 27752 39238
rect 27816 39030 27844 39238
rect 27804 39024 27856 39030
rect 27804 38966 27856 38972
rect 27632 38916 27752 38944
rect 27632 38758 27660 38916
rect 27804 38888 27856 38894
rect 27802 38856 27804 38865
rect 27856 38856 27858 38865
rect 27712 38820 27764 38826
rect 27802 38791 27858 38800
rect 27712 38762 27764 38768
rect 27620 38752 27672 38758
rect 27620 38694 27672 38700
rect 27724 38654 27752 38762
rect 27632 38626 27752 38654
rect 27632 37244 27660 38626
rect 27908 38486 27936 41618
rect 28000 40118 28028 41958
rect 28080 41472 28132 41478
rect 28078 41440 28080 41449
rect 28132 41440 28134 41449
rect 28078 41375 28134 41384
rect 28080 40996 28132 41002
rect 28080 40938 28132 40944
rect 27988 40112 28040 40118
rect 27988 40054 28040 40060
rect 27988 39976 28040 39982
rect 27988 39918 28040 39924
rect 28000 38978 28028 39918
rect 28092 39420 28120 40938
rect 28184 40769 28212 42622
rect 28264 42560 28316 42566
rect 28264 42502 28316 42508
rect 28276 41993 28304 42502
rect 28262 41984 28318 41993
rect 28262 41919 28318 41928
rect 28262 41304 28318 41313
rect 28262 41239 28318 41248
rect 28170 40760 28226 40769
rect 28170 40695 28172 40704
rect 28224 40695 28226 40704
rect 28172 40666 28224 40672
rect 28170 40080 28226 40089
rect 28170 40015 28226 40024
rect 28184 39574 28212 40015
rect 28172 39568 28224 39574
rect 28172 39510 28224 39516
rect 28172 39432 28224 39438
rect 28092 39392 28172 39420
rect 28172 39374 28224 39380
rect 28170 39264 28226 39273
rect 28170 39199 28226 39208
rect 28078 38992 28134 39001
rect 28000 38950 28078 38978
rect 28078 38927 28134 38936
rect 27988 38752 28040 38758
rect 27988 38694 28040 38700
rect 27896 38480 27948 38486
rect 27896 38422 27948 38428
rect 27804 37936 27856 37942
rect 27804 37878 27856 37884
rect 27816 37670 27844 37878
rect 27908 37806 27936 38422
rect 27896 37800 27948 37806
rect 27896 37742 27948 37748
rect 27804 37664 27856 37670
rect 27804 37606 27856 37612
rect 27816 37330 27844 37606
rect 27804 37324 27856 37330
rect 27804 37266 27856 37272
rect 27712 37256 27764 37262
rect 27632 37216 27712 37244
rect 27712 37198 27764 37204
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27632 34678 27660 36178
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27804 35012 27856 35018
rect 27804 34954 27856 34960
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 27816 34610 27844 34954
rect 27908 34678 27936 35974
rect 27896 34672 27948 34678
rect 27896 34614 27948 34620
rect 27804 34604 27856 34610
rect 27804 34546 27856 34552
rect 27448 34428 27568 34456
rect 27710 34504 27766 34513
rect 27710 34439 27766 34448
rect 27448 33862 27476 34428
rect 27526 34368 27582 34377
rect 27526 34303 27582 34312
rect 27540 34066 27568 34303
rect 27724 34066 27752 34439
rect 28000 34406 28028 38694
rect 28092 36582 28120 38927
rect 28184 36786 28212 39199
rect 28276 37942 28304 41239
rect 28368 39642 28396 45222
rect 28460 43246 28488 46310
rect 28448 43240 28500 43246
rect 28448 43182 28500 43188
rect 28448 42560 28500 42566
rect 28448 42502 28500 42508
rect 28460 42401 28488 42502
rect 28446 42392 28502 42401
rect 28446 42327 28502 42336
rect 28552 40458 28580 46310
rect 28644 45529 28672 47126
rect 28908 47116 28960 47122
rect 28908 47058 28960 47064
rect 28920 46918 28948 47058
rect 28724 46912 28776 46918
rect 28724 46854 28776 46860
rect 28908 46912 28960 46918
rect 28908 46854 28960 46860
rect 28736 46714 28764 46854
rect 28724 46708 28776 46714
rect 28724 46650 28776 46656
rect 29184 46572 29236 46578
rect 29184 46514 29236 46520
rect 28908 46436 28960 46442
rect 28908 46378 28960 46384
rect 28920 45966 28948 46378
rect 28908 45960 28960 45966
rect 28908 45902 28960 45908
rect 29196 45898 29224 46514
rect 29276 46368 29328 46374
rect 29276 46310 29328 46316
rect 29288 46170 29316 46310
rect 29276 46164 29328 46170
rect 29276 46106 29328 46112
rect 29184 45892 29236 45898
rect 29184 45834 29236 45840
rect 29092 45552 29144 45558
rect 28630 45520 28686 45529
rect 29092 45494 29144 45500
rect 28908 45484 28960 45490
rect 28630 45455 28686 45464
rect 28644 43790 28672 45455
rect 28736 45444 28908 45472
rect 28736 45014 28764 45444
rect 28908 45426 28960 45432
rect 28724 45008 28776 45014
rect 28724 44950 28776 44956
rect 28632 43784 28684 43790
rect 28632 43726 28684 43732
rect 28632 42288 28684 42294
rect 28632 42230 28684 42236
rect 28540 40452 28592 40458
rect 28540 40394 28592 40400
rect 28644 40225 28672 42230
rect 28736 41478 28764 44950
rect 29104 44878 29132 45494
rect 29092 44872 29144 44878
rect 29092 44814 29144 44820
rect 28908 44736 28960 44742
rect 28908 44678 28960 44684
rect 28920 44402 28948 44678
rect 28908 44396 28960 44402
rect 28908 44338 28960 44344
rect 29092 44192 29144 44198
rect 29092 44134 29144 44140
rect 29104 43926 29132 44134
rect 29092 43920 29144 43926
rect 29092 43862 29144 43868
rect 29184 43852 29236 43858
rect 29184 43794 29236 43800
rect 28908 43648 28960 43654
rect 28908 43590 28960 43596
rect 28816 42356 28868 42362
rect 28816 42298 28868 42304
rect 28828 42226 28856 42298
rect 28816 42220 28868 42226
rect 28816 42162 28868 42168
rect 28816 41540 28868 41546
rect 28816 41482 28868 41488
rect 28724 41472 28776 41478
rect 28828 41449 28856 41482
rect 28724 41414 28776 41420
rect 28814 41440 28870 41449
rect 28736 41313 28764 41414
rect 28814 41375 28870 41384
rect 28722 41304 28778 41313
rect 28722 41239 28778 41248
rect 28816 41268 28868 41274
rect 28816 41210 28868 41216
rect 28828 40934 28856 41210
rect 28816 40928 28868 40934
rect 28816 40870 28868 40876
rect 28724 40520 28776 40526
rect 28724 40462 28776 40468
rect 28630 40216 28686 40225
rect 28630 40151 28686 40160
rect 28736 40118 28764 40462
rect 28540 40112 28592 40118
rect 28540 40054 28592 40060
rect 28724 40112 28776 40118
rect 28724 40054 28776 40060
rect 28356 39636 28408 39642
rect 28356 39578 28408 39584
rect 28446 38992 28502 39001
rect 28446 38927 28448 38936
rect 28500 38927 28502 38936
rect 28448 38898 28500 38904
rect 28356 38888 28408 38894
rect 28356 38830 28408 38836
rect 28264 37936 28316 37942
rect 28264 37878 28316 37884
rect 28368 37466 28396 38830
rect 28446 38720 28502 38729
rect 28446 38655 28502 38664
rect 28460 37874 28488 38655
rect 28448 37868 28500 37874
rect 28448 37810 28500 37816
rect 28448 37732 28500 37738
rect 28448 37674 28500 37680
rect 28356 37460 28408 37466
rect 28356 37402 28408 37408
rect 28460 37262 28488 37674
rect 28552 37369 28580 40054
rect 28816 40044 28868 40050
rect 28816 39986 28868 39992
rect 28632 39840 28684 39846
rect 28632 39782 28684 39788
rect 28644 38758 28672 39782
rect 28828 39642 28856 39986
rect 28816 39636 28868 39642
rect 28816 39578 28868 39584
rect 28920 39488 28948 43590
rect 29196 43450 29224 43794
rect 29184 43444 29236 43450
rect 29184 43386 29236 43392
rect 29092 42832 29144 42838
rect 29092 42774 29144 42780
rect 29104 42226 29132 42774
rect 29288 42702 29316 46106
rect 29380 45898 29408 47534
rect 29748 47462 29776 47942
rect 31760 47728 31812 47734
rect 31760 47670 31812 47676
rect 31024 47524 31076 47530
rect 31024 47466 31076 47472
rect 29736 47456 29788 47462
rect 29736 47398 29788 47404
rect 29748 46578 29776 47398
rect 31036 47054 31064 47466
rect 31300 47456 31352 47462
rect 31300 47398 31352 47404
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 31024 47048 31076 47054
rect 31024 46990 31076 46996
rect 30104 46980 30156 46986
rect 30104 46922 30156 46928
rect 29736 46572 29788 46578
rect 29736 46514 29788 46520
rect 29736 46368 29788 46374
rect 29736 46310 29788 46316
rect 29748 45966 29776 46310
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29368 45892 29420 45898
rect 29368 45834 29420 45840
rect 29380 44878 29408 45834
rect 29748 45558 29776 45902
rect 29736 45552 29788 45558
rect 29736 45494 29788 45500
rect 30116 45286 30144 46922
rect 30656 46640 30708 46646
rect 30656 46582 30708 46588
rect 30288 46436 30340 46442
rect 30288 46378 30340 46384
rect 30300 45966 30328 46378
rect 30668 46374 30696 46582
rect 30656 46368 30708 46374
rect 30656 46310 30708 46316
rect 30668 46034 30696 46310
rect 30748 46096 30800 46102
rect 30748 46038 30800 46044
rect 30656 46028 30708 46034
rect 30656 45970 30708 45976
rect 30288 45960 30340 45966
rect 30288 45902 30340 45908
rect 30668 45490 30696 45970
rect 30656 45484 30708 45490
rect 30656 45426 30708 45432
rect 29736 45280 29788 45286
rect 29736 45222 29788 45228
rect 30104 45280 30156 45286
rect 30104 45222 30156 45228
rect 29368 44872 29420 44878
rect 29368 44814 29420 44820
rect 29644 44804 29696 44810
rect 29644 44746 29696 44752
rect 29656 44470 29684 44746
rect 29644 44464 29696 44470
rect 29644 44406 29696 44412
rect 29552 44396 29604 44402
rect 29552 44338 29604 44344
rect 29368 44192 29420 44198
rect 29368 44134 29420 44140
rect 29458 44160 29514 44169
rect 29380 43314 29408 44134
rect 29458 44095 29514 44104
rect 29472 43722 29500 44095
rect 29460 43716 29512 43722
rect 29460 43658 29512 43664
rect 29368 43308 29420 43314
rect 29368 43250 29420 43256
rect 29460 43308 29512 43314
rect 29460 43250 29512 43256
rect 29276 42696 29328 42702
rect 29276 42638 29328 42644
rect 29092 42220 29144 42226
rect 29092 42162 29144 42168
rect 29288 41682 29316 42638
rect 29276 41676 29328 41682
rect 29276 41618 29328 41624
rect 29274 41168 29330 41177
rect 29274 41103 29276 41112
rect 29328 41103 29330 41112
rect 29276 41074 29328 41080
rect 29184 40384 29236 40390
rect 29184 40326 29236 40332
rect 28998 40080 29054 40089
rect 29196 40050 29224 40326
rect 28998 40015 29000 40024
rect 29052 40015 29054 40024
rect 29184 40044 29236 40050
rect 29000 39986 29052 39992
rect 29184 39986 29236 39992
rect 28828 39460 28948 39488
rect 28722 38856 28778 38865
rect 28722 38791 28778 38800
rect 28632 38752 28684 38758
rect 28632 38694 28684 38700
rect 28736 38418 28764 38791
rect 28828 38468 28856 39460
rect 29092 39432 29144 39438
rect 29092 39374 29144 39380
rect 29276 39432 29328 39438
rect 29276 39374 29328 39380
rect 29104 39302 29132 39374
rect 29092 39296 29144 39302
rect 29092 39238 29144 39244
rect 29090 39128 29146 39137
rect 29090 39063 29146 39072
rect 29000 39024 29052 39030
rect 29000 38966 29052 38972
rect 28908 38480 28960 38486
rect 28828 38440 28908 38468
rect 28908 38422 28960 38428
rect 28724 38412 28776 38418
rect 28724 38354 28776 38360
rect 28632 37868 28684 37874
rect 28632 37810 28684 37816
rect 28538 37360 28594 37369
rect 28538 37295 28594 37304
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 28080 36576 28132 36582
rect 28080 36518 28132 36524
rect 28276 36174 28304 37198
rect 28644 36938 28672 37810
rect 28736 37738 28764 38354
rect 28816 38208 28868 38214
rect 28816 38150 28868 38156
rect 28724 37732 28776 37738
rect 28724 37674 28776 37680
rect 28828 37194 28856 38150
rect 28920 37670 28948 38422
rect 29012 38282 29040 38966
rect 29104 38350 29132 39063
rect 29184 38956 29236 38962
rect 29184 38898 29236 38904
rect 29092 38344 29144 38350
rect 29092 38286 29144 38292
rect 29000 38276 29052 38282
rect 29000 38218 29052 38224
rect 28908 37664 28960 37670
rect 28908 37606 28960 37612
rect 28908 37392 28960 37398
rect 28908 37334 28960 37340
rect 28816 37188 28868 37194
rect 28816 37130 28868 37136
rect 28552 36910 28764 36938
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 28080 35828 28132 35834
rect 28080 35770 28132 35776
rect 28092 34610 28120 35770
rect 28276 34626 28304 36110
rect 28460 35698 28488 36518
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28552 35086 28580 36910
rect 28736 36854 28764 36910
rect 28632 36848 28684 36854
rect 28632 36790 28684 36796
rect 28724 36848 28776 36854
rect 28724 36790 28776 36796
rect 28644 36310 28672 36790
rect 28724 36712 28776 36718
rect 28724 36654 28776 36660
rect 28632 36304 28684 36310
rect 28632 36246 28684 36252
rect 28736 36106 28764 36654
rect 28724 36100 28776 36106
rect 28724 36042 28776 36048
rect 28540 35080 28592 35086
rect 28540 35022 28592 35028
rect 28736 35018 28764 36042
rect 28828 35154 28856 37130
rect 28920 36378 28948 37334
rect 29012 36922 29040 38218
rect 29196 37670 29224 38898
rect 29288 38865 29316 39374
rect 29274 38856 29330 38865
rect 29274 38791 29330 38800
rect 29288 37874 29316 38791
rect 29276 37868 29328 37874
rect 29276 37810 29328 37816
rect 29184 37664 29236 37670
rect 29184 37606 29236 37612
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 29012 36378 29040 36722
rect 28908 36372 28960 36378
rect 28908 36314 28960 36320
rect 29000 36372 29052 36378
rect 29000 36314 29052 36320
rect 29012 35834 29040 36314
rect 29196 36174 29224 37606
rect 29184 36168 29236 36174
rect 29184 36110 29236 36116
rect 29000 35828 29052 35834
rect 29196 35816 29224 36110
rect 29000 35770 29052 35776
rect 29104 35788 29224 35816
rect 28908 35692 28960 35698
rect 28908 35634 28960 35640
rect 28816 35148 28868 35154
rect 28816 35090 28868 35096
rect 28920 35086 28948 35634
rect 29104 35630 29132 35788
rect 29182 35728 29238 35737
rect 29182 35663 29184 35672
rect 29236 35663 29238 35672
rect 29184 35634 29236 35640
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29092 35488 29144 35494
rect 29092 35430 29144 35436
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 28724 35012 28776 35018
rect 28724 34954 28776 34960
rect 29000 34944 29052 34950
rect 28814 34912 28870 34921
rect 29000 34886 29052 34892
rect 28814 34847 28870 34856
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28184 34598 28304 34626
rect 28828 34610 28856 34847
rect 29012 34746 29040 34886
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 28816 34604 28868 34610
rect 27988 34400 28040 34406
rect 27988 34342 28040 34348
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27712 34060 27764 34066
rect 27712 34002 27764 34008
rect 27436 33856 27488 33862
rect 27436 33798 27488 33804
rect 28184 33658 28212 34598
rect 28816 34546 28868 34552
rect 28264 34400 28316 34406
rect 28264 34342 28316 34348
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 28172 33652 28224 33658
rect 28172 33594 28224 33600
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 28276 32978 28304 34342
rect 29012 34066 29040 34342
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 29104 33998 29132 35430
rect 29196 35170 29224 35634
rect 29380 35222 29408 43250
rect 29472 42770 29500 43250
rect 29460 42764 29512 42770
rect 29460 42706 29512 42712
rect 29472 42226 29500 42706
rect 29460 42220 29512 42226
rect 29460 42162 29512 42168
rect 29472 42090 29500 42162
rect 29460 42084 29512 42090
rect 29460 42026 29512 42032
rect 29564 41614 29592 44338
rect 29748 44266 29776 45222
rect 30564 44940 30616 44946
rect 30564 44882 30616 44888
rect 29828 44872 29880 44878
rect 29828 44814 29880 44820
rect 30288 44872 30340 44878
rect 30288 44814 30340 44820
rect 29840 44538 29868 44814
rect 30012 44736 30064 44742
rect 30012 44678 30064 44684
rect 29828 44532 29880 44538
rect 29828 44474 29880 44480
rect 29736 44260 29788 44266
rect 29656 44220 29736 44248
rect 29656 42362 29684 44220
rect 29736 44202 29788 44208
rect 29920 43988 29972 43994
rect 29920 43930 29972 43936
rect 29828 43784 29880 43790
rect 29828 43726 29880 43732
rect 29736 43648 29788 43654
rect 29736 43590 29788 43596
rect 29748 42945 29776 43590
rect 29840 43178 29868 43726
rect 29828 43172 29880 43178
rect 29828 43114 29880 43120
rect 29734 42936 29790 42945
rect 29932 42906 29960 43930
rect 30024 43790 30052 44678
rect 30300 44402 30328 44814
rect 30288 44396 30340 44402
rect 30288 44338 30340 44344
rect 30380 44328 30432 44334
rect 30380 44270 30432 44276
rect 30012 43784 30064 43790
rect 30012 43726 30064 43732
rect 30196 43172 30248 43178
rect 30196 43114 30248 43120
rect 30012 43104 30064 43110
rect 30012 43046 30064 43052
rect 29734 42871 29790 42880
rect 29920 42900 29972 42906
rect 29920 42842 29972 42848
rect 30024 42702 30052 43046
rect 29736 42696 29788 42702
rect 30012 42696 30064 42702
rect 29736 42638 29788 42644
rect 29932 42656 30012 42684
rect 29644 42356 29696 42362
rect 29644 42298 29696 42304
rect 29748 41614 29776 42638
rect 29828 42560 29880 42566
rect 29828 42502 29880 42508
rect 29552 41608 29604 41614
rect 29736 41608 29788 41614
rect 29552 41550 29604 41556
rect 29656 41568 29736 41596
rect 29564 41414 29592 41550
rect 29472 41386 29592 41414
rect 29472 38758 29500 41386
rect 29550 39944 29606 39953
rect 29550 39879 29606 39888
rect 29564 39846 29592 39879
rect 29552 39840 29604 39846
rect 29552 39782 29604 39788
rect 29656 39409 29684 41568
rect 29736 41550 29788 41556
rect 29736 39976 29788 39982
rect 29736 39918 29788 39924
rect 29748 39438 29776 39918
rect 29840 39574 29868 42502
rect 29932 41614 29960 42656
rect 30012 42638 30064 42644
rect 30012 42288 30064 42294
rect 30012 42230 30064 42236
rect 29920 41608 29972 41614
rect 29920 41550 29972 41556
rect 29932 41206 29960 41550
rect 30024 41478 30052 42230
rect 30012 41472 30064 41478
rect 30012 41414 30064 41420
rect 29920 41200 29972 41206
rect 29920 41142 29972 41148
rect 29920 40996 29972 41002
rect 29920 40938 29972 40944
rect 29932 40526 29960 40938
rect 29920 40520 29972 40526
rect 29920 40462 29972 40468
rect 29828 39568 29880 39574
rect 29828 39510 29880 39516
rect 29840 39438 29868 39510
rect 29736 39432 29788 39438
rect 29642 39400 29698 39409
rect 29736 39374 29788 39380
rect 29828 39432 29880 39438
rect 29828 39374 29880 39380
rect 29642 39335 29698 39344
rect 29656 38962 29684 39335
rect 29748 39030 29776 39374
rect 29736 39024 29788 39030
rect 29736 38966 29788 38972
rect 29932 38962 29960 40462
rect 30024 39846 30052 41414
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 30116 39846 30144 41074
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 30104 39840 30156 39846
rect 30104 39782 30156 39788
rect 29644 38956 29696 38962
rect 29644 38898 29696 38904
rect 29920 38956 29972 38962
rect 29920 38898 29972 38904
rect 29828 38888 29880 38894
rect 29828 38830 29880 38836
rect 29736 38820 29788 38826
rect 29736 38762 29788 38768
rect 29460 38752 29512 38758
rect 29460 38694 29512 38700
rect 29644 38752 29696 38758
rect 29644 38694 29696 38700
rect 29472 38282 29500 38694
rect 29460 38276 29512 38282
rect 29460 38218 29512 38224
rect 29472 37806 29500 38218
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29656 36786 29684 38694
rect 29748 38214 29776 38762
rect 29840 38654 29868 38830
rect 30024 38758 30052 39782
rect 30116 39370 30144 39782
rect 30104 39364 30156 39370
rect 30104 39306 30156 39312
rect 30012 38752 30064 38758
rect 30012 38694 30064 38700
rect 29840 38626 30052 38654
rect 30024 38214 30052 38626
rect 29736 38208 29788 38214
rect 29736 38150 29788 38156
rect 30012 38208 30064 38214
rect 30012 38150 30064 38156
rect 29644 36780 29696 36786
rect 29644 36722 29696 36728
rect 29748 36718 29776 38150
rect 29828 37732 29880 37738
rect 29828 37674 29880 37680
rect 29736 36712 29788 36718
rect 29736 36654 29788 36660
rect 29644 36576 29696 36582
rect 29644 36518 29696 36524
rect 29552 35624 29604 35630
rect 29552 35566 29604 35572
rect 29368 35216 29420 35222
rect 29196 35142 29316 35170
rect 29368 35158 29420 35164
rect 29458 35184 29514 35193
rect 29184 35012 29236 35018
rect 29184 34954 29236 34960
rect 29092 33992 29144 33998
rect 29092 33934 29144 33940
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28724 33856 28776 33862
rect 28724 33798 28776 33804
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 26976 32224 27028 32230
rect 26976 32166 27028 32172
rect 26988 32026 27016 32166
rect 26976 32020 27028 32026
rect 26976 31962 27028 31968
rect 26884 31952 26936 31958
rect 26884 31894 26936 31900
rect 26896 30938 26924 31894
rect 27172 31890 27200 32846
rect 27356 32524 27568 32552
rect 27252 32496 27304 32502
rect 27250 32464 27252 32473
rect 27304 32464 27306 32473
rect 27250 32399 27306 32408
rect 27252 32224 27304 32230
rect 27252 32166 27304 32172
rect 27264 31958 27292 32166
rect 27252 31952 27304 31958
rect 27252 31894 27304 31900
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26988 31482 27016 31758
rect 27068 31748 27120 31754
rect 27068 31690 27120 31696
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 26884 30932 26936 30938
rect 26884 30874 26936 30880
rect 26988 30734 27016 31418
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 27080 30598 27108 31690
rect 27356 31396 27384 32524
rect 27540 32434 27568 32524
rect 28356 32496 28408 32502
rect 28356 32438 28408 32444
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27448 31498 27476 32370
rect 28368 32026 28396 32438
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27448 31470 27660 31498
rect 27632 31414 27660 31470
rect 27436 31408 27488 31414
rect 27356 31368 27436 31396
rect 27620 31408 27672 31414
rect 27488 31368 27568 31396
rect 27436 31350 27488 31356
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 26884 30592 26936 30598
rect 26884 30534 26936 30540
rect 27068 30592 27120 30598
rect 27068 30534 27120 30540
rect 26896 29646 26924 30534
rect 27080 30326 27108 30534
rect 27068 30320 27120 30326
rect 27068 30262 27120 30268
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26976 29096 27028 29102
rect 26976 29038 27028 29044
rect 26988 28422 27016 29038
rect 26976 28416 27028 28422
rect 26976 28358 27028 28364
rect 26976 27600 27028 27606
rect 26976 27542 27028 27548
rect 26988 27334 27016 27542
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 27172 27130 27200 31078
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27448 29170 27476 30534
rect 27540 30394 27568 31368
rect 27620 31350 27672 31356
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27540 29850 27568 30330
rect 27632 30190 27660 31350
rect 27816 30598 27844 31690
rect 28368 31142 28396 31962
rect 28356 31136 28408 31142
rect 28356 31078 28408 31084
rect 28460 30734 28488 33798
rect 28736 33658 28764 33798
rect 28724 33652 28776 33658
rect 28724 33594 28776 33600
rect 29196 33386 29224 34954
rect 29288 34610 29316 35142
rect 29458 35119 29460 35128
rect 29512 35119 29514 35128
rect 29460 35090 29512 35096
rect 29276 34604 29328 34610
rect 29276 34546 29328 34552
rect 29184 33380 29236 33386
rect 29184 33322 29236 33328
rect 29092 32972 29144 32978
rect 29092 32914 29144 32920
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 28828 32434 28856 32846
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 29104 32366 29132 32914
rect 29368 32428 29420 32434
rect 29368 32370 29420 32376
rect 29092 32360 29144 32366
rect 29092 32302 29144 32308
rect 28632 31680 28684 31686
rect 28632 31622 28684 31628
rect 28538 31376 28594 31385
rect 28644 31346 28672 31622
rect 28538 31311 28594 31320
rect 28632 31340 28684 31346
rect 28552 31278 28580 31311
rect 28632 31282 28684 31288
rect 28540 31272 28592 31278
rect 28540 31214 28592 31220
rect 28264 30728 28316 30734
rect 28264 30670 28316 30676
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 27804 30592 27856 30598
rect 27804 30534 27856 30540
rect 28276 30433 28304 30670
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28262 30424 28318 30433
rect 28262 30359 28318 30368
rect 28460 30258 28488 30534
rect 28644 30394 28672 31282
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28632 30388 28684 30394
rect 28632 30330 28684 30336
rect 28736 30258 28764 30670
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 27620 30184 27672 30190
rect 27620 30126 27672 30132
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 27528 29844 27580 29850
rect 27528 29786 27580 29792
rect 27632 29730 27660 30126
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 27540 29702 27660 29730
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27540 29102 27568 29702
rect 28920 29646 28948 29990
rect 29012 29714 29040 30126
rect 29104 29850 29132 32302
rect 29184 31748 29236 31754
rect 29184 31690 29236 31696
rect 29196 31346 29224 31690
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 29196 30938 29224 31282
rect 29184 30932 29236 30938
rect 29184 30874 29236 30880
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 29092 29844 29144 29850
rect 29092 29786 29144 29792
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29012 29306 29040 29650
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 27528 29096 27580 29102
rect 27528 29038 27580 29044
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 28172 29096 28224 29102
rect 28172 29038 28224 29044
rect 27540 28422 27568 29038
rect 27632 28558 27660 29038
rect 28184 28558 28212 29038
rect 28552 28558 28580 29106
rect 29104 28558 29132 29786
rect 29288 29714 29316 30534
rect 29380 30326 29408 32370
rect 29564 30598 29592 35566
rect 29656 31346 29684 36518
rect 29840 35766 29868 37674
rect 29920 36916 29972 36922
rect 29920 36858 29972 36864
rect 29828 35760 29880 35766
rect 29828 35702 29880 35708
rect 29840 35154 29868 35702
rect 29932 35698 29960 36858
rect 30024 36854 30052 38150
rect 30116 37210 30144 39306
rect 30208 39098 30236 43114
rect 30288 42900 30340 42906
rect 30288 42842 30340 42848
rect 30300 42226 30328 42842
rect 30288 42220 30340 42226
rect 30288 42162 30340 42168
rect 30392 40934 30420 44270
rect 30576 43994 30604 44882
rect 30668 44810 30696 45426
rect 30656 44804 30708 44810
rect 30656 44746 30708 44752
rect 30564 43988 30616 43994
rect 30564 43930 30616 43936
rect 30656 43784 30708 43790
rect 30656 43726 30708 43732
rect 30472 43716 30524 43722
rect 30472 43658 30524 43664
rect 30484 42226 30512 43658
rect 30668 42906 30696 43726
rect 30656 42900 30708 42906
rect 30656 42842 30708 42848
rect 30760 42294 30788 46038
rect 30944 45626 30972 46990
rect 31036 45626 31064 46990
rect 31312 46986 31340 47398
rect 31772 47122 31800 47670
rect 32600 47666 32628 48286
rect 32588 47660 32640 47666
rect 32588 47602 32640 47608
rect 32600 47258 32628 47602
rect 33232 47592 33284 47598
rect 33232 47534 33284 47540
rect 32588 47252 32640 47258
rect 32588 47194 32640 47200
rect 31760 47116 31812 47122
rect 31760 47058 31812 47064
rect 31300 46980 31352 46986
rect 31300 46922 31352 46928
rect 31312 46578 31340 46922
rect 31300 46572 31352 46578
rect 31300 46514 31352 46520
rect 31208 46164 31260 46170
rect 31208 46106 31260 46112
rect 31220 45626 31248 46106
rect 31300 45824 31352 45830
rect 31300 45766 31352 45772
rect 30932 45620 30984 45626
rect 30932 45562 30984 45568
rect 31024 45620 31076 45626
rect 31208 45620 31260 45626
rect 31076 45580 31156 45608
rect 31024 45562 31076 45568
rect 30840 45348 30892 45354
rect 30840 45290 30892 45296
rect 30748 42288 30800 42294
rect 30748 42230 30800 42236
rect 30472 42220 30524 42226
rect 30472 42162 30524 42168
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 30288 40928 30340 40934
rect 30288 40870 30340 40876
rect 30380 40928 30432 40934
rect 30380 40870 30432 40876
rect 30300 40746 30328 40870
rect 30300 40718 30420 40746
rect 30288 40384 30340 40390
rect 30288 40326 30340 40332
rect 30300 40186 30328 40326
rect 30288 40180 30340 40186
rect 30288 40122 30340 40128
rect 30288 39500 30340 39506
rect 30288 39442 30340 39448
rect 30196 39092 30248 39098
rect 30196 39034 30248 39040
rect 30300 38962 30328 39442
rect 30392 39438 30420 40718
rect 30380 39432 30432 39438
rect 30380 39374 30432 39380
rect 30484 39273 30512 42162
rect 30668 41818 30696 42162
rect 30748 42016 30800 42022
rect 30748 41958 30800 41964
rect 30656 41812 30708 41818
rect 30656 41754 30708 41760
rect 30760 41614 30788 41958
rect 30748 41608 30800 41614
rect 30748 41550 30800 41556
rect 30564 40656 30616 40662
rect 30564 40598 30616 40604
rect 30576 40390 30604 40598
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30576 39642 30604 40326
rect 30564 39636 30616 39642
rect 30564 39578 30616 39584
rect 30470 39264 30526 39273
rect 30470 39199 30526 39208
rect 30380 39092 30432 39098
rect 30380 39034 30432 39040
rect 30472 39092 30524 39098
rect 30472 39034 30524 39040
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 30288 38956 30340 38962
rect 30288 38898 30340 38904
rect 30208 38486 30236 38898
rect 30196 38480 30248 38486
rect 30196 38422 30248 38428
rect 30392 38350 30420 39034
rect 30380 38344 30432 38350
rect 30380 38286 30432 38292
rect 30484 37992 30512 39034
rect 30576 38554 30604 39578
rect 30656 38752 30708 38758
rect 30656 38694 30708 38700
rect 30564 38548 30616 38554
rect 30564 38490 30616 38496
rect 30484 37964 30604 37992
rect 30472 37868 30524 37874
rect 30472 37810 30524 37816
rect 30380 37664 30432 37670
rect 30380 37606 30432 37612
rect 30196 37460 30248 37466
rect 30196 37402 30248 37408
rect 30208 37330 30236 37402
rect 30288 37392 30340 37398
rect 30286 37360 30288 37369
rect 30340 37360 30342 37369
rect 30196 37324 30248 37330
rect 30286 37295 30342 37304
rect 30196 37266 30248 37272
rect 30116 37182 30236 37210
rect 30104 37120 30156 37126
rect 30104 37062 30156 37068
rect 30012 36848 30064 36854
rect 30012 36790 30064 36796
rect 30116 36718 30144 37062
rect 30104 36712 30156 36718
rect 30104 36654 30156 36660
rect 30104 36372 30156 36378
rect 30104 36314 30156 36320
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 30116 35154 30144 36314
rect 29828 35148 29880 35154
rect 29828 35090 29880 35096
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 29748 34610 29776 35022
rect 29840 34678 29868 35090
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29828 34672 29880 34678
rect 29828 34614 29880 34620
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29840 34066 29868 34614
rect 29932 34542 29960 35022
rect 30208 34610 30236 37182
rect 30288 37120 30340 37126
rect 30286 37088 30288 37097
rect 30340 37088 30342 37097
rect 30286 37023 30342 37032
rect 30392 36174 30420 37606
rect 30484 36786 30512 37810
rect 30576 37097 30604 37964
rect 30562 37088 30618 37097
rect 30562 37023 30618 37032
rect 30472 36780 30524 36786
rect 30472 36722 30524 36728
rect 30576 36174 30604 37023
rect 30668 36242 30696 38694
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30760 36786 30788 38286
rect 30852 37244 30880 45290
rect 30944 44878 30972 45562
rect 31024 45484 31076 45490
rect 31024 45426 31076 45432
rect 30932 44872 30984 44878
rect 30932 44814 30984 44820
rect 31036 44198 31064 45426
rect 31128 44402 31156 45580
rect 31208 45562 31260 45568
rect 31312 45490 31340 45766
rect 31300 45484 31352 45490
rect 31300 45426 31352 45432
rect 31312 45370 31340 45426
rect 31312 45342 31432 45370
rect 31300 45280 31352 45286
rect 31300 45222 31352 45228
rect 31312 44742 31340 45222
rect 31300 44736 31352 44742
rect 31300 44678 31352 44684
rect 31116 44396 31168 44402
rect 31116 44338 31168 44344
rect 31024 44192 31076 44198
rect 31024 44134 31076 44140
rect 31036 43790 31064 44134
rect 31128 43926 31156 44338
rect 31208 43988 31260 43994
rect 31208 43930 31260 43936
rect 31116 43920 31168 43926
rect 31116 43862 31168 43868
rect 31024 43784 31076 43790
rect 31024 43726 31076 43732
rect 31116 43784 31168 43790
rect 31116 43726 31168 43732
rect 30932 41608 30984 41614
rect 30932 41550 30984 41556
rect 30944 41002 30972 41550
rect 31036 41274 31064 43726
rect 31024 41268 31076 41274
rect 31024 41210 31076 41216
rect 30932 40996 30984 41002
rect 30932 40938 30984 40944
rect 31036 40594 31064 41210
rect 31024 40588 31076 40594
rect 31024 40530 31076 40536
rect 30932 39636 30984 39642
rect 30932 39578 30984 39584
rect 30944 39506 30972 39578
rect 30932 39500 30984 39506
rect 30932 39442 30984 39448
rect 31128 38842 31156 43726
rect 31220 41818 31248 43930
rect 31312 43790 31340 44678
rect 31404 44402 31432 45342
rect 31392 44396 31444 44402
rect 31392 44338 31444 44344
rect 31300 43784 31352 43790
rect 31300 43726 31352 43732
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31208 41812 31260 41818
rect 31208 41754 31260 41760
rect 31220 39438 31248 41754
rect 31312 41750 31340 43046
rect 31300 41744 31352 41750
rect 31300 41686 31352 41692
rect 31404 41614 31432 44338
rect 31484 43648 31536 43654
rect 31484 43590 31536 43596
rect 31496 42208 31524 43590
rect 31668 43240 31720 43246
rect 31668 43182 31720 43188
rect 31576 42220 31628 42226
rect 31496 42180 31576 42208
rect 31392 41608 31444 41614
rect 31392 41550 31444 41556
rect 31496 41460 31524 42180
rect 31576 42162 31628 42168
rect 31576 41608 31628 41614
rect 31576 41550 31628 41556
rect 31404 41432 31524 41460
rect 31300 40384 31352 40390
rect 31300 40326 31352 40332
rect 31208 39432 31260 39438
rect 31208 39374 31260 39380
rect 31312 38962 31340 40326
rect 31300 38956 31352 38962
rect 31300 38898 31352 38904
rect 31036 38814 31156 38842
rect 30932 37460 30984 37466
rect 30932 37402 30984 37408
rect 30944 37369 30972 37402
rect 30930 37360 30986 37369
rect 31036 37346 31064 38814
rect 31116 38752 31168 38758
rect 31114 38720 31116 38729
rect 31168 38720 31170 38729
rect 31114 38655 31170 38664
rect 31300 38344 31352 38350
rect 31300 38286 31352 38292
rect 31208 38208 31260 38214
rect 31208 38150 31260 38156
rect 31220 37670 31248 38150
rect 31208 37664 31260 37670
rect 31208 37606 31260 37612
rect 31036 37318 31156 37346
rect 30930 37295 30986 37304
rect 30932 37256 30984 37262
rect 30852 37216 30932 37244
rect 30748 36780 30800 36786
rect 30748 36722 30800 36728
rect 30852 36378 30880 37216
rect 30932 37198 30984 37204
rect 31024 37188 31076 37194
rect 31024 37130 31076 37136
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 30944 36582 30972 37062
rect 30932 36576 30984 36582
rect 30932 36518 30984 36524
rect 31036 36394 31064 37130
rect 31128 36786 31156 37318
rect 31208 37120 31260 37126
rect 31208 37062 31260 37068
rect 31116 36780 31168 36786
rect 31116 36722 31168 36728
rect 31116 36576 31168 36582
rect 31116 36518 31168 36524
rect 30840 36372 30892 36378
rect 30840 36314 30892 36320
rect 30944 36366 31064 36394
rect 30656 36236 30708 36242
rect 30656 36178 30708 36184
rect 30380 36168 30432 36174
rect 30380 36110 30432 36116
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30300 35698 30328 35974
rect 30470 35728 30526 35737
rect 30288 35692 30340 35698
rect 30470 35663 30526 35672
rect 30288 35634 30340 35640
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 29828 34060 29880 34066
rect 29828 34002 29880 34008
rect 30484 33590 30512 35663
rect 30576 35018 30604 36110
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30852 35290 30880 35430
rect 30840 35284 30892 35290
rect 30840 35226 30892 35232
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30564 35012 30616 35018
rect 30564 34954 30616 34960
rect 30656 34536 30708 34542
rect 30852 34524 30880 35022
rect 30944 35018 30972 36366
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 31036 35154 31064 36110
rect 31128 35698 31156 36518
rect 31116 35692 31168 35698
rect 31116 35634 31168 35640
rect 31024 35148 31076 35154
rect 31024 35090 31076 35096
rect 30932 35012 30984 35018
rect 30932 34954 30984 34960
rect 31036 34542 31064 35090
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 31128 34610 31156 34886
rect 31116 34604 31168 34610
rect 31116 34546 31168 34552
rect 30932 34536 30984 34542
rect 30852 34496 30932 34524
rect 30656 34478 30708 34484
rect 30932 34478 30984 34484
rect 31024 34536 31076 34542
rect 31024 34478 31076 34484
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30472 33584 30524 33590
rect 30472 33526 30524 33532
rect 30288 33516 30340 33522
rect 30288 33458 30340 33464
rect 30300 32570 30328 33458
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30392 32026 30420 32302
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30484 32026 30512 32234
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30576 31890 30604 33798
rect 30668 32502 30696 34478
rect 30944 34066 30972 34478
rect 31024 34128 31076 34134
rect 31024 34070 31076 34076
rect 31116 34128 31168 34134
rect 31116 34070 31168 34076
rect 30932 34060 30984 34066
rect 30932 34002 30984 34008
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30656 32496 30708 32502
rect 30656 32438 30708 32444
rect 30564 31884 30616 31890
rect 30564 31826 30616 31832
rect 29644 31340 29696 31346
rect 29644 31282 29696 31288
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 29552 30592 29604 30598
rect 29552 30534 29604 30540
rect 29368 30320 29420 30326
rect 29368 30262 29420 30268
rect 29276 29708 29328 29714
rect 29276 29650 29328 29656
rect 30116 29646 30144 31214
rect 30852 30802 30880 33254
rect 31036 31346 31064 34070
rect 31128 33998 31156 34070
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 31220 33522 31248 37062
rect 31312 36718 31340 38286
rect 31404 37874 31432 41432
rect 31484 41268 31536 41274
rect 31484 41210 31536 41216
rect 31496 40050 31524 41210
rect 31484 40044 31536 40050
rect 31484 39986 31536 39992
rect 31588 39846 31616 41550
rect 31576 39840 31628 39846
rect 31576 39782 31628 39788
rect 31588 38457 31616 39782
rect 31680 38865 31708 43182
rect 31772 42702 31800 47058
rect 32312 46912 32364 46918
rect 32312 46854 32364 46860
rect 32324 46646 32352 46854
rect 32312 46640 32364 46646
rect 32312 46582 32364 46588
rect 32496 46572 32548 46578
rect 32496 46514 32548 46520
rect 32312 46504 32364 46510
rect 32508 46458 32536 46514
rect 32600 46510 32628 47194
rect 33140 46640 33192 46646
rect 33140 46582 33192 46588
rect 32364 46452 32536 46458
rect 32312 46446 32536 46452
rect 32588 46504 32640 46510
rect 32588 46446 32640 46452
rect 32324 46430 32536 46446
rect 31852 46368 31904 46374
rect 31852 46310 31904 46316
rect 31864 46034 31892 46310
rect 31852 46028 31904 46034
rect 31852 45970 31904 45976
rect 32508 45966 32536 46430
rect 32496 45960 32548 45966
rect 32496 45902 32548 45908
rect 32312 45348 32364 45354
rect 32508 45336 32536 45902
rect 32588 45348 32640 45354
rect 32508 45308 32588 45336
rect 32312 45290 32364 45296
rect 32588 45290 32640 45296
rect 32128 45008 32180 45014
rect 32128 44950 32180 44956
rect 31852 44464 31904 44470
rect 31852 44406 31904 44412
rect 31864 43926 31892 44406
rect 31852 43920 31904 43926
rect 31852 43862 31904 43868
rect 31760 42696 31812 42702
rect 31760 42638 31812 42644
rect 31864 42634 31892 43862
rect 32140 43450 32168 44950
rect 32324 44538 32352 45290
rect 32496 44940 32548 44946
rect 32496 44882 32548 44888
rect 32312 44532 32364 44538
rect 32312 44474 32364 44480
rect 32128 43444 32180 43450
rect 32128 43386 32180 43392
rect 31944 42832 31996 42838
rect 31944 42774 31996 42780
rect 31852 42628 31904 42634
rect 31852 42570 31904 42576
rect 31956 42514 31984 42774
rect 31772 42486 31984 42514
rect 31772 41274 31800 42486
rect 31852 42356 31904 42362
rect 31852 42298 31904 42304
rect 31760 41268 31812 41274
rect 31760 41210 31812 41216
rect 31760 40044 31812 40050
rect 31760 39986 31812 39992
rect 31772 39953 31800 39986
rect 31758 39944 31814 39953
rect 31758 39879 31814 39888
rect 31666 38856 31722 38865
rect 31666 38791 31722 38800
rect 31574 38448 31630 38457
rect 31574 38383 31630 38392
rect 31484 38004 31536 38010
rect 31484 37946 31536 37952
rect 31392 37868 31444 37874
rect 31392 37810 31444 37816
rect 31496 37670 31524 37946
rect 31392 37664 31444 37670
rect 31392 37606 31444 37612
rect 31484 37664 31536 37670
rect 31484 37606 31536 37612
rect 31300 36712 31352 36718
rect 31300 36654 31352 36660
rect 31312 36378 31340 36654
rect 31300 36372 31352 36378
rect 31300 36314 31352 36320
rect 31404 35834 31432 37606
rect 31588 36802 31616 38383
rect 31668 37936 31720 37942
rect 31668 37878 31720 37884
rect 31680 37720 31708 37878
rect 31864 37720 31892 42298
rect 31944 42220 31996 42226
rect 31944 42162 31996 42168
rect 31956 41750 31984 42162
rect 32036 42016 32088 42022
rect 32036 41958 32088 41964
rect 31944 41744 31996 41750
rect 31944 41686 31996 41692
rect 31956 41449 31984 41686
rect 31942 41440 31998 41449
rect 31942 41375 31998 41384
rect 31944 40724 31996 40730
rect 31944 40666 31996 40672
rect 31956 40594 31984 40666
rect 31944 40588 31996 40594
rect 31944 40530 31996 40536
rect 32048 40526 32076 41958
rect 32140 41274 32168 43386
rect 32324 42650 32352 44474
rect 32404 44192 32456 44198
rect 32404 44134 32456 44140
rect 32416 43790 32444 44134
rect 32404 43784 32456 43790
rect 32404 43726 32456 43732
rect 32416 43382 32444 43726
rect 32404 43376 32456 43382
rect 32404 43318 32456 43324
rect 32416 42770 32444 43318
rect 32404 42764 32456 42770
rect 32404 42706 32456 42712
rect 32324 42622 32444 42650
rect 32312 42288 32364 42294
rect 32312 42230 32364 42236
rect 32128 41268 32180 41274
rect 32128 41210 32180 41216
rect 32220 41132 32272 41138
rect 32220 41074 32272 41080
rect 32128 40996 32180 41002
rect 32128 40938 32180 40944
rect 32036 40520 32088 40526
rect 32036 40462 32088 40468
rect 32140 40118 32168 40938
rect 32232 40186 32260 41074
rect 32324 40934 32352 42230
rect 32416 41414 32444 42622
rect 32508 41562 32536 44882
rect 32600 43722 32628 45290
rect 33152 44878 33180 46582
rect 33140 44872 33192 44878
rect 33140 44814 33192 44820
rect 33244 44810 33272 47534
rect 34428 47456 34480 47462
rect 34428 47398 34480 47404
rect 33600 46980 33652 46986
rect 33600 46922 33652 46928
rect 33324 46912 33376 46918
rect 33324 46854 33376 46860
rect 33336 46714 33364 46854
rect 33324 46708 33376 46714
rect 33324 46650 33376 46656
rect 33336 46034 33364 46650
rect 33324 46028 33376 46034
rect 33324 45970 33376 45976
rect 33336 45490 33364 45970
rect 33612 45966 33640 46922
rect 33968 46912 34020 46918
rect 33968 46854 34020 46860
rect 33784 46368 33836 46374
rect 33784 46310 33836 46316
rect 33796 45966 33824 46310
rect 33600 45960 33652 45966
rect 33600 45902 33652 45908
rect 33784 45960 33836 45966
rect 33784 45902 33836 45908
rect 33416 45620 33468 45626
rect 33416 45562 33468 45568
rect 33324 45484 33376 45490
rect 33324 45426 33376 45432
rect 33232 44804 33284 44810
rect 33232 44746 33284 44752
rect 33244 44334 33272 44746
rect 33336 44402 33364 45426
rect 33324 44396 33376 44402
rect 33324 44338 33376 44344
rect 33232 44328 33284 44334
rect 33232 44270 33284 44276
rect 32770 44160 32826 44169
rect 32770 44095 32826 44104
rect 32588 43716 32640 43722
rect 32588 43658 32640 43664
rect 32600 42770 32628 43658
rect 32680 43104 32732 43110
rect 32680 43046 32732 43052
rect 32588 42764 32640 42770
rect 32588 42706 32640 42712
rect 32586 42528 32642 42537
rect 32586 42463 32642 42472
rect 32600 42022 32628 42463
rect 32692 42226 32720 43046
rect 32680 42220 32732 42226
rect 32680 42162 32732 42168
rect 32588 42016 32640 42022
rect 32588 41958 32640 41964
rect 32600 41750 32628 41958
rect 32588 41744 32640 41750
rect 32588 41686 32640 41692
rect 32508 41534 32628 41562
rect 32416 41386 32536 41414
rect 32312 40928 32364 40934
rect 32312 40870 32364 40876
rect 32312 40724 32364 40730
rect 32312 40666 32364 40672
rect 32220 40180 32272 40186
rect 32220 40122 32272 40128
rect 32128 40112 32180 40118
rect 32128 40054 32180 40060
rect 32128 39976 32180 39982
rect 32128 39918 32180 39924
rect 32140 39642 32168 39918
rect 32220 39840 32272 39846
rect 32220 39782 32272 39788
rect 32128 39636 32180 39642
rect 32128 39578 32180 39584
rect 32128 39296 32180 39302
rect 32128 39238 32180 39244
rect 32140 38962 32168 39238
rect 32128 38956 32180 38962
rect 32128 38898 32180 38904
rect 32034 38856 32090 38865
rect 31944 38820 31996 38826
rect 32034 38791 32090 38800
rect 31944 38762 31996 38768
rect 31956 38457 31984 38762
rect 31942 38448 31998 38457
rect 31942 38383 31998 38392
rect 31944 38344 31996 38350
rect 31944 38286 31996 38292
rect 31956 38010 31984 38286
rect 31944 38004 31996 38010
rect 31944 37946 31996 37952
rect 31680 37692 31892 37720
rect 31668 37392 31720 37398
rect 31668 37334 31720 37340
rect 31680 36922 31708 37334
rect 31772 37262 31800 37692
rect 32048 37670 32076 38791
rect 32140 37738 32168 38898
rect 32128 37732 32180 37738
rect 32128 37674 32180 37680
rect 32036 37664 32088 37670
rect 32036 37606 32088 37612
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 31484 36780 31536 36786
rect 31588 36774 31708 36802
rect 31484 36722 31536 36728
rect 31496 36582 31524 36722
rect 31484 36576 31536 36582
rect 31484 36518 31536 36524
rect 31496 36174 31524 36518
rect 31484 36168 31536 36174
rect 31484 36110 31536 36116
rect 31392 35828 31444 35834
rect 31392 35770 31444 35776
rect 31484 35148 31536 35154
rect 31484 35090 31536 35096
rect 31392 34536 31444 34542
rect 31392 34478 31444 34484
rect 31404 33930 31432 34478
rect 31496 33998 31524 35090
rect 31576 34944 31628 34950
rect 31576 34886 31628 34892
rect 31484 33992 31536 33998
rect 31484 33934 31536 33940
rect 31392 33924 31444 33930
rect 31392 33866 31444 33872
rect 31300 33856 31352 33862
rect 31300 33798 31352 33804
rect 31312 33590 31340 33798
rect 31300 33584 31352 33590
rect 31300 33526 31352 33532
rect 31404 33522 31432 33866
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 31312 32774 31340 33050
rect 31116 32768 31168 32774
rect 31116 32710 31168 32716
rect 31300 32768 31352 32774
rect 31300 32710 31352 32716
rect 31128 32230 31156 32710
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31116 32224 31168 32230
rect 31116 32166 31168 32172
rect 31128 31822 31156 32166
rect 31220 31890 31248 32370
rect 31208 31884 31260 31890
rect 31208 31826 31260 31832
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 31392 31408 31444 31414
rect 31392 31350 31444 31356
rect 31024 31340 31076 31346
rect 31024 31282 31076 31288
rect 31036 30802 31064 31282
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 31024 30796 31076 30802
rect 31024 30738 31076 30744
rect 31404 30734 31432 31350
rect 31484 31340 31536 31346
rect 31484 31282 31536 31288
rect 31496 30938 31524 31282
rect 31484 30932 31536 30938
rect 31484 30874 31536 30880
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 30932 30592 30984 30598
rect 30932 30534 30984 30540
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 29656 29170 29684 29582
rect 30116 29170 30144 29582
rect 30840 29572 30892 29578
rect 30840 29514 30892 29520
rect 30852 29238 30880 29514
rect 30944 29238 30972 30534
rect 31588 30258 31616 34886
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31312 29510 31340 29786
rect 31680 29594 31708 36774
rect 32128 36100 32180 36106
rect 32128 36042 32180 36048
rect 31944 36032 31996 36038
rect 31944 35974 31996 35980
rect 31852 35148 31904 35154
rect 31852 35090 31904 35096
rect 31864 35018 31892 35090
rect 31956 35086 31984 35974
rect 32140 35086 32168 36042
rect 32232 35737 32260 39782
rect 32324 38418 32352 40666
rect 32508 40526 32536 41386
rect 32600 41070 32628 41534
rect 32692 41206 32720 42162
rect 32784 41585 32812 44095
rect 33336 43722 33364 44338
rect 33428 43994 33456 45562
rect 33612 45490 33640 45902
rect 33600 45484 33652 45490
rect 33600 45426 33652 45432
rect 33612 44878 33640 45426
rect 33508 44872 33560 44878
rect 33508 44814 33560 44820
rect 33600 44872 33652 44878
rect 33600 44814 33652 44820
rect 33520 44402 33548 44814
rect 33508 44396 33560 44402
rect 33508 44338 33560 44344
rect 33612 44282 33640 44814
rect 33520 44254 33640 44282
rect 33416 43988 33468 43994
rect 33416 43930 33468 43936
rect 33324 43716 33376 43722
rect 33324 43658 33376 43664
rect 33520 43246 33548 44254
rect 33690 43344 33746 43353
rect 33690 43279 33692 43288
rect 33744 43279 33746 43288
rect 33692 43250 33744 43256
rect 33508 43240 33560 43246
rect 33508 43182 33560 43188
rect 32956 42832 33008 42838
rect 32956 42774 33008 42780
rect 32770 41576 32826 41585
rect 32770 41511 32826 41520
rect 32784 41478 32812 41511
rect 32772 41472 32824 41478
rect 32772 41414 32824 41420
rect 32680 41200 32732 41206
rect 32732 41160 32904 41188
rect 32680 41142 32732 41148
rect 32588 41064 32640 41070
rect 32640 41012 32812 41018
rect 32588 41006 32812 41012
rect 32600 40990 32812 41006
rect 32600 40941 32628 40990
rect 32680 40928 32732 40934
rect 32680 40870 32732 40876
rect 32404 40520 32456 40526
rect 32404 40462 32456 40468
rect 32496 40520 32548 40526
rect 32496 40462 32548 40468
rect 32416 39030 32444 40462
rect 32496 40384 32548 40390
rect 32496 40326 32548 40332
rect 32508 40186 32536 40326
rect 32496 40180 32548 40186
rect 32496 40122 32548 40128
rect 32508 39574 32536 40122
rect 32496 39568 32548 39574
rect 32496 39510 32548 39516
rect 32496 39432 32548 39438
rect 32496 39374 32548 39380
rect 32508 39302 32536 39374
rect 32496 39296 32548 39302
rect 32496 39238 32548 39244
rect 32404 39024 32456 39030
rect 32404 38966 32456 38972
rect 32312 38412 32364 38418
rect 32312 38354 32364 38360
rect 32416 35766 32444 38966
rect 32588 38956 32640 38962
rect 32588 38898 32640 38904
rect 32600 38554 32628 38898
rect 32588 38548 32640 38554
rect 32588 38490 32640 38496
rect 32588 38412 32640 38418
rect 32588 38354 32640 38360
rect 32496 38344 32548 38350
rect 32496 38286 32548 38292
rect 32508 37874 32536 38286
rect 32496 37868 32548 37874
rect 32496 37810 32548 37816
rect 32600 37466 32628 38354
rect 32588 37460 32640 37466
rect 32588 37402 32640 37408
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 32496 36780 32548 36786
rect 32600 36768 32628 37198
rect 32692 36786 32720 40870
rect 32784 39506 32812 40990
rect 32772 39500 32824 39506
rect 32772 39442 32824 39448
rect 32876 39370 32904 41160
rect 32968 39574 32996 42774
rect 33520 42634 33548 43182
rect 33796 42702 33824 45902
rect 33980 45830 34008 46854
rect 34152 46368 34204 46374
rect 34152 46310 34204 46316
rect 33876 45824 33928 45830
rect 33874 45792 33876 45801
rect 33968 45824 34020 45830
rect 33928 45792 33930 45801
rect 33968 45766 34020 45772
rect 33874 45727 33930 45736
rect 33980 45490 34008 45766
rect 33968 45484 34020 45490
rect 33968 45426 34020 45432
rect 34164 45082 34192 46310
rect 34440 45490 34468 47398
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34704 46368 34756 46374
rect 34704 46310 34756 46316
rect 34716 45830 34744 46310
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34704 45824 34756 45830
rect 34704 45766 34756 45772
rect 34520 45552 34572 45558
rect 34520 45494 34572 45500
rect 34428 45484 34480 45490
rect 34428 45426 34480 45432
rect 34440 45286 34468 45426
rect 34428 45280 34480 45286
rect 34428 45222 34480 45228
rect 34152 45076 34204 45082
rect 34152 45018 34204 45024
rect 34164 44538 34192 45018
rect 34152 44532 34204 44538
rect 34152 44474 34204 44480
rect 34428 44464 34480 44470
rect 34428 44406 34480 44412
rect 34440 44334 34468 44406
rect 34428 44328 34480 44334
rect 34428 44270 34480 44276
rect 33876 44260 33928 44266
rect 33876 44202 33928 44208
rect 33888 44169 33916 44202
rect 33874 44160 33930 44169
rect 33874 44095 33930 44104
rect 33876 43988 33928 43994
rect 33876 43930 33928 43936
rect 33784 42696 33836 42702
rect 33784 42638 33836 42644
rect 33048 42628 33100 42634
rect 33048 42570 33100 42576
rect 33508 42628 33560 42634
rect 33508 42570 33560 42576
rect 33060 42226 33088 42570
rect 33416 42560 33468 42566
rect 33416 42502 33468 42508
rect 33140 42356 33192 42362
rect 33140 42298 33192 42304
rect 33048 42220 33100 42226
rect 33048 42162 33100 42168
rect 33060 41682 33088 42162
rect 33048 41676 33100 41682
rect 33048 41618 33100 41624
rect 33060 41002 33088 41618
rect 33152 41138 33180 42298
rect 33140 41132 33192 41138
rect 33140 41074 33192 41080
rect 33048 40996 33100 41002
rect 33048 40938 33100 40944
rect 32956 39568 33008 39574
rect 32956 39510 33008 39516
rect 32864 39364 32916 39370
rect 32864 39306 32916 39312
rect 32876 38486 32904 39306
rect 32968 39098 32996 39510
rect 32956 39092 33008 39098
rect 32956 39034 33008 39040
rect 32864 38480 32916 38486
rect 32864 38422 32916 38428
rect 33060 37874 33088 40938
rect 33152 38962 33180 41074
rect 33232 40928 33284 40934
rect 33232 40870 33284 40876
rect 33140 38956 33192 38962
rect 33140 38898 33192 38904
rect 33048 37868 33100 37874
rect 33048 37810 33100 37816
rect 33152 37262 33180 38898
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32548 36740 32628 36768
rect 32680 36780 32732 36786
rect 32496 36722 32548 36728
rect 32732 36740 32812 36768
rect 32680 36722 32732 36728
rect 32404 35760 32456 35766
rect 32218 35728 32274 35737
rect 32404 35702 32456 35708
rect 32218 35663 32274 35672
rect 32508 35494 32536 36722
rect 32680 36236 32732 36242
rect 32680 36178 32732 36184
rect 32692 35834 32720 36178
rect 32784 36174 32812 36740
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 33152 36174 33180 36314
rect 32772 36168 32824 36174
rect 32772 36110 32824 36116
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 32680 35828 32732 35834
rect 32680 35770 32732 35776
rect 32956 35624 33008 35630
rect 33008 35572 33180 35578
rect 32956 35566 33180 35572
rect 32968 35550 33180 35566
rect 32496 35488 32548 35494
rect 32496 35430 32548 35436
rect 32508 35086 32536 35430
rect 33048 35216 33100 35222
rect 33048 35158 33100 35164
rect 33060 35086 33088 35158
rect 31944 35080 31996 35086
rect 31944 35022 31996 35028
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 32496 35080 32548 35086
rect 32496 35022 32548 35028
rect 33048 35080 33100 35086
rect 33048 35022 33100 35028
rect 31852 35012 31904 35018
rect 31852 34954 31904 34960
rect 31760 34060 31812 34066
rect 31760 34002 31812 34008
rect 31772 33658 31800 34002
rect 31864 33862 31892 34954
rect 33152 34950 33180 35550
rect 32680 34944 32732 34950
rect 32680 34886 32732 34892
rect 33140 34944 33192 34950
rect 33140 34886 33192 34892
rect 31944 34536 31996 34542
rect 31944 34478 31996 34484
rect 31852 33856 31904 33862
rect 31852 33798 31904 33804
rect 31760 33652 31812 33658
rect 31760 33594 31812 33600
rect 31956 33114 31984 34478
rect 32128 34128 32180 34134
rect 32128 34070 32180 34076
rect 31944 33108 31996 33114
rect 31944 33050 31996 33056
rect 32140 32910 32168 34070
rect 32692 33998 32720 34886
rect 33140 34672 33192 34678
rect 33140 34614 33192 34620
rect 33048 34468 33100 34474
rect 33048 34410 33100 34416
rect 32680 33992 32732 33998
rect 32680 33934 32732 33940
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 32220 33448 32272 33454
rect 32220 33390 32272 33396
rect 32232 32978 32260 33390
rect 32508 33114 32536 33458
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 32220 32972 32272 32978
rect 32220 32914 32272 32920
rect 32692 32910 32720 33934
rect 32772 33856 32824 33862
rect 32772 33798 32824 33804
rect 32784 33522 32812 33798
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32784 32978 32812 33458
rect 32956 33312 33008 33318
rect 32956 33254 33008 33260
rect 32772 32972 32824 32978
rect 32772 32914 32824 32920
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32680 32904 32732 32910
rect 32680 32846 32732 32852
rect 31772 32774 31800 32846
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 32140 32366 32168 32846
rect 32692 32434 32720 32846
rect 32784 32774 32812 32914
rect 32772 32768 32824 32774
rect 32772 32710 32824 32716
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 32140 30870 32168 32302
rect 32968 31890 32996 33254
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32588 31680 32640 31686
rect 32588 31622 32640 31628
rect 32128 30864 32180 30870
rect 32128 30806 32180 30812
rect 32496 30864 32548 30870
rect 32496 30806 32548 30812
rect 32140 30190 32168 30806
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32508 30054 32536 30806
rect 32600 30734 32628 31622
rect 32692 31482 32720 31758
rect 32680 31476 32732 31482
rect 32680 31418 32732 31424
rect 32968 31414 32996 31826
rect 32956 31408 33008 31414
rect 32956 31350 33008 31356
rect 32956 31136 33008 31142
rect 32956 31078 33008 31084
rect 32968 30734 32996 31078
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32772 30252 32824 30258
rect 32772 30194 32824 30200
rect 32496 30048 32548 30054
rect 32496 29990 32548 29996
rect 31588 29578 31708 29594
rect 31576 29572 31708 29578
rect 31628 29566 31708 29572
rect 31576 29514 31628 29520
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 30840 29232 30892 29238
rect 30840 29174 30892 29180
rect 30932 29232 30984 29238
rect 30984 29180 31064 29186
rect 30932 29174 31064 29180
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30852 29050 30880 29174
rect 30944 29158 31064 29174
rect 31312 29170 31340 29446
rect 31484 29232 31536 29238
rect 31484 29174 31536 29180
rect 29828 29028 29880 29034
rect 30852 29022 30972 29050
rect 29828 28970 29880 28976
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 28082 27568 28358
rect 27632 28150 27660 28494
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27252 28008 27304 28014
rect 27252 27950 27304 27956
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 26332 26444 26384 26450
rect 26332 26386 26384 26392
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 24216 26308 24268 26314
rect 24216 26250 24268 26256
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 26344 25838 26372 26386
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 27080 25702 27108 26318
rect 27172 26042 27200 26862
rect 27160 26036 27212 26042
rect 27160 25978 27212 25984
rect 27264 25838 27292 27950
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 27448 27062 27476 27270
rect 27540 27062 27568 28018
rect 28184 27674 28212 28494
rect 28552 28218 28580 28494
rect 29104 28234 29132 28494
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 29012 28206 29132 28234
rect 29012 28150 29040 28206
rect 29196 28150 29224 28426
rect 29000 28144 29052 28150
rect 29000 28086 29052 28092
rect 29184 28144 29236 28150
rect 29184 28086 29236 28092
rect 29840 27878 29868 28970
rect 30104 28960 30156 28966
rect 30104 28902 30156 28908
rect 30380 28960 30432 28966
rect 30380 28902 30432 28908
rect 30116 28490 30144 28902
rect 30104 28484 30156 28490
rect 30104 28426 30156 28432
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 28184 27334 28212 27610
rect 30392 27606 30420 28902
rect 30944 28558 30972 29022
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30932 28552 30984 28558
rect 30932 28494 30984 28500
rect 30760 27606 30788 28494
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30748 27600 30800 27606
rect 30748 27542 30800 27548
rect 31036 27470 31064 29158
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31496 28694 31524 29174
rect 32312 29096 32364 29102
rect 32310 29064 32312 29073
rect 32364 29064 32366 29073
rect 32310 28999 32366 29008
rect 31484 28688 31536 28694
rect 31484 28630 31536 28636
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31128 28150 31156 28358
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 32416 28014 32444 29446
rect 32508 28558 32536 29990
rect 32680 29028 32732 29034
rect 32600 28976 32680 28994
rect 32600 28970 32732 28976
rect 32600 28966 32720 28970
rect 32588 28960 32640 28966
rect 32588 28902 32640 28908
rect 32784 28558 32812 30194
rect 33060 29646 33088 34410
rect 33152 33998 33180 34614
rect 33140 33992 33192 33998
rect 33140 33934 33192 33940
rect 33152 33590 33180 33934
rect 33140 33584 33192 33590
rect 33140 33526 33192 33532
rect 33244 33114 33272 40870
rect 33428 40526 33456 42502
rect 33416 40520 33468 40526
rect 33416 40462 33468 40468
rect 33324 40384 33376 40390
rect 33324 40326 33376 40332
rect 33336 40118 33364 40326
rect 33324 40112 33376 40118
rect 33324 40054 33376 40060
rect 33520 39914 33548 42570
rect 33692 42560 33744 42566
rect 33692 42502 33744 42508
rect 33704 42294 33732 42502
rect 33692 42288 33744 42294
rect 33692 42230 33744 42236
rect 33600 41812 33652 41818
rect 33600 41754 33652 41760
rect 33612 41614 33640 41754
rect 33600 41608 33652 41614
rect 33600 41550 33652 41556
rect 33704 41478 33732 42230
rect 33784 41540 33836 41546
rect 33784 41482 33836 41488
rect 33692 41472 33744 41478
rect 33692 41414 33744 41420
rect 33796 41274 33824 41482
rect 33784 41268 33836 41274
rect 33784 41210 33836 41216
rect 33600 41200 33652 41206
rect 33600 41142 33652 41148
rect 33690 41168 33746 41177
rect 33508 39908 33560 39914
rect 33508 39850 33560 39856
rect 33612 39522 33640 41142
rect 33690 41103 33692 41112
rect 33744 41103 33746 41112
rect 33692 41074 33744 41080
rect 33704 40662 33732 41074
rect 33784 40996 33836 41002
rect 33784 40938 33836 40944
rect 33692 40656 33744 40662
rect 33692 40598 33744 40604
rect 33796 40474 33824 40938
rect 33336 39494 33640 39522
rect 33704 40446 33824 40474
rect 33336 38418 33364 39494
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33520 38418 33548 39374
rect 33704 39302 33732 40446
rect 33888 40066 33916 43930
rect 33968 42016 34020 42022
rect 33968 41958 34020 41964
rect 33980 41449 34008 41958
rect 33966 41440 34022 41449
rect 33966 41375 34022 41384
rect 33980 41138 34008 41375
rect 33968 41132 34020 41138
rect 33968 41074 34020 41080
rect 33796 40038 33916 40066
rect 33692 39296 33744 39302
rect 33692 39238 33744 39244
rect 33600 38888 33652 38894
rect 33600 38830 33652 38836
rect 33324 38412 33376 38418
rect 33324 38354 33376 38360
rect 33508 38412 33560 38418
rect 33508 38354 33560 38360
rect 33336 37330 33364 38354
rect 33324 37324 33376 37330
rect 33324 37266 33376 37272
rect 33520 37194 33548 38354
rect 33612 37670 33640 38830
rect 33600 37664 33652 37670
rect 33600 37606 33652 37612
rect 33612 37398 33640 37606
rect 33600 37392 33652 37398
rect 33600 37334 33652 37340
rect 33508 37188 33560 37194
rect 33508 37130 33560 37136
rect 33416 36304 33468 36310
rect 33416 36246 33468 36252
rect 33324 35080 33376 35086
rect 33428 35068 33456 36246
rect 33520 36174 33548 37130
rect 33612 37126 33640 37334
rect 33600 37120 33652 37126
rect 33600 37062 33652 37068
rect 33612 36786 33640 37062
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33520 35834 33548 36110
rect 33508 35828 33560 35834
rect 33508 35770 33560 35776
rect 33520 35154 33548 35770
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 33376 35040 33456 35068
rect 33600 35080 33652 35086
rect 33324 35022 33376 35028
rect 33600 35022 33652 35028
rect 33324 34944 33376 34950
rect 33324 34886 33376 34892
rect 33416 34944 33468 34950
rect 33416 34886 33468 34892
rect 33336 34610 33364 34886
rect 33324 34604 33376 34610
rect 33324 34546 33376 34552
rect 33428 34134 33456 34886
rect 33416 34128 33468 34134
rect 33416 34070 33468 34076
rect 33612 33590 33640 35022
rect 33704 34610 33732 39238
rect 33796 37806 33824 40038
rect 33876 39976 33928 39982
rect 33876 39918 33928 39924
rect 33888 39098 33916 39918
rect 34060 39432 34112 39438
rect 34060 39374 34112 39380
rect 33876 39092 33928 39098
rect 33876 39034 33928 39040
rect 34072 38894 34100 39374
rect 34532 39370 34560 45494
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35348 44192 35400 44198
rect 35348 44134 35400 44140
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34978 43888 35034 43897
rect 34978 43823 34980 43832
rect 35032 43823 35034 43832
rect 34980 43794 35032 43800
rect 35360 43790 35388 44134
rect 35348 43784 35400 43790
rect 35348 43726 35400 43732
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34796 42220 34848 42226
rect 34796 42162 34848 42168
rect 34704 42152 34756 42158
rect 34704 42094 34756 42100
rect 34716 41818 34744 42094
rect 34704 41812 34756 41818
rect 34704 41754 34756 41760
rect 34808 41614 34836 42162
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41750 35388 43726
rect 35440 43308 35492 43314
rect 35440 43250 35492 43256
rect 35348 41744 35400 41750
rect 35348 41686 35400 41692
rect 34796 41608 34848 41614
rect 34610 41576 34666 41585
rect 34796 41550 34848 41556
rect 34610 41511 34666 41520
rect 34520 39364 34572 39370
rect 34520 39306 34572 39312
rect 34244 39296 34296 39302
rect 34244 39238 34296 39244
rect 34256 38894 34284 39238
rect 34532 39098 34560 39306
rect 34520 39092 34572 39098
rect 34520 39034 34572 39040
rect 34532 38962 34560 39034
rect 34520 38956 34572 38962
rect 34520 38898 34572 38904
rect 34624 38894 34652 41511
rect 35164 41472 35216 41478
rect 35164 41414 35216 41420
rect 35176 41070 35204 41414
rect 35164 41064 35216 41070
rect 35164 41006 35216 41012
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40526 35388 41686
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34796 38956 34848 38962
rect 34796 38898 34848 38904
rect 34060 38888 34112 38894
rect 34060 38830 34112 38836
rect 34244 38888 34296 38894
rect 34244 38830 34296 38836
rect 34336 38888 34388 38894
rect 34336 38830 34388 38836
rect 34612 38888 34664 38894
rect 34612 38830 34664 38836
rect 34152 38208 34204 38214
rect 34152 38150 34204 38156
rect 33784 37800 33836 37806
rect 33784 37742 33836 37748
rect 33876 37460 33928 37466
rect 33876 37402 33928 37408
rect 33888 36922 33916 37402
rect 33968 37256 34020 37262
rect 33968 37198 34020 37204
rect 34060 37256 34112 37262
rect 34060 37198 34112 37204
rect 33876 36916 33928 36922
rect 33876 36858 33928 36864
rect 33784 36780 33836 36786
rect 33784 36722 33836 36728
rect 33876 36780 33928 36786
rect 33980 36768 34008 37198
rect 33928 36740 34008 36768
rect 33876 36722 33928 36728
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33600 33584 33652 33590
rect 33600 33526 33652 33532
rect 33796 33402 33824 36722
rect 33888 36310 33916 36722
rect 34072 36650 34100 37198
rect 34060 36644 34112 36650
rect 34060 36586 34112 36592
rect 33876 36304 33928 36310
rect 33876 36246 33928 36252
rect 33968 36032 34020 36038
rect 33968 35974 34020 35980
rect 33876 34604 33928 34610
rect 33876 34546 33928 34552
rect 33888 33658 33916 34546
rect 33980 34542 34008 35974
rect 34058 35184 34114 35193
rect 34058 35119 34114 35128
rect 34072 35086 34100 35119
rect 34060 35080 34112 35086
rect 34060 35022 34112 35028
rect 34060 34672 34112 34678
rect 34060 34614 34112 34620
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 33428 33374 33824 33402
rect 33232 33108 33284 33114
rect 33232 33050 33284 33056
rect 33244 32434 33272 33050
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 33428 29714 33456 33374
rect 34072 33114 34100 34614
rect 34164 33590 34192 38150
rect 34348 38010 34376 38830
rect 34428 38820 34480 38826
rect 34428 38762 34480 38768
rect 34336 38004 34388 38010
rect 34336 37946 34388 37952
rect 34440 37466 34468 38762
rect 34520 38752 34572 38758
rect 34520 38694 34572 38700
rect 34428 37460 34480 37466
rect 34428 37402 34480 37408
rect 34336 37188 34388 37194
rect 34336 37130 34388 37136
rect 34348 36174 34376 37130
rect 34336 36168 34388 36174
rect 34336 36110 34388 36116
rect 34348 35986 34376 36110
rect 34256 35958 34376 35986
rect 34256 35766 34284 35958
rect 34244 35760 34296 35766
rect 34244 35702 34296 35708
rect 34532 35630 34560 38694
rect 34624 38554 34652 38830
rect 34704 38752 34756 38758
rect 34704 38694 34756 38700
rect 34612 38548 34664 38554
rect 34612 38490 34664 38496
rect 34716 38010 34744 38694
rect 34704 38004 34756 38010
rect 34704 37946 34756 37952
rect 34704 37868 34756 37874
rect 34808 37856 34836 38898
rect 35360 38894 35388 40462
rect 35452 40186 35480 43250
rect 35440 40180 35492 40186
rect 35440 40122 35492 40128
rect 35440 39500 35492 39506
rect 35440 39442 35492 39448
rect 35072 38888 35124 38894
rect 35072 38830 35124 38836
rect 35348 38888 35400 38894
rect 35348 38830 35400 38836
rect 35084 38758 35112 38830
rect 35072 38752 35124 38758
rect 35072 38694 35124 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35452 38418 35480 39442
rect 35440 38412 35492 38418
rect 35440 38354 35492 38360
rect 35348 38276 35400 38282
rect 35348 38218 35400 38224
rect 35360 38010 35388 38218
rect 35348 38004 35400 38010
rect 35348 37946 35400 37952
rect 34756 37828 34836 37856
rect 34704 37810 34756 37816
rect 34716 36242 34744 37810
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34980 37120 35032 37126
rect 34980 37062 35032 37068
rect 34992 36786 35020 37062
rect 34980 36780 35032 36786
rect 34980 36722 35032 36728
rect 35452 36718 35480 38354
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 35440 36712 35492 36718
rect 35440 36654 35492 36660
rect 34704 36236 34756 36242
rect 34704 36178 34756 36184
rect 34520 35624 34572 35630
rect 34520 35566 34572 35572
rect 34428 33992 34480 33998
rect 34428 33934 34480 33940
rect 34152 33584 34204 33590
rect 34152 33526 34204 33532
rect 34440 33386 34468 33934
rect 34428 33380 34480 33386
rect 34428 33322 34480 33328
rect 34060 33108 34112 33114
rect 34060 33050 34112 33056
rect 33600 32768 33652 32774
rect 33600 32710 33652 32716
rect 33612 32434 33640 32710
rect 34072 32434 34100 33050
rect 34440 33046 34468 33322
rect 34428 33040 34480 33046
rect 34428 32982 34480 32988
rect 33600 32428 33652 32434
rect 33600 32370 33652 32376
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 34060 32428 34112 32434
rect 34060 32370 34112 32376
rect 33508 32360 33560 32366
rect 33508 32302 33560 32308
rect 33520 31822 33548 32302
rect 33612 32230 33640 32370
rect 33692 32292 33744 32298
rect 33692 32234 33744 32240
rect 33600 32224 33652 32230
rect 33600 32166 33652 32172
rect 33508 31816 33560 31822
rect 33508 31758 33560 31764
rect 33600 30660 33652 30666
rect 33600 30602 33652 30608
rect 33612 30054 33640 30602
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33704 29850 33732 32234
rect 33796 31890 33824 32370
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 33888 31890 33916 32166
rect 34072 31890 34100 32370
rect 34428 32360 34480 32366
rect 34428 32302 34480 32308
rect 33784 31884 33836 31890
rect 33784 31826 33836 31832
rect 33876 31884 33928 31890
rect 33876 31826 33928 31832
rect 34060 31884 34112 31890
rect 34060 31826 34112 31832
rect 34440 31754 34468 32302
rect 34348 31726 34468 31754
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 31482 34100 31622
rect 34060 31476 34112 31482
rect 34060 31418 34112 31424
rect 33968 31272 34020 31278
rect 33968 31214 34020 31220
rect 33980 30734 34008 31214
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 33980 30326 34008 30670
rect 33968 30320 34020 30326
rect 33968 30262 34020 30268
rect 34072 30258 34100 31418
rect 34244 31408 34296 31414
rect 34244 31350 34296 31356
rect 34152 30932 34204 30938
rect 34152 30874 34204 30880
rect 34164 30326 34192 30874
rect 34256 30802 34284 31350
rect 34348 31142 34376 31726
rect 34336 31136 34388 31142
rect 34336 31078 34388 31084
rect 34244 30796 34296 30802
rect 34244 30738 34296 30744
rect 34152 30320 34204 30326
rect 34152 30262 34204 30268
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 34348 30190 34376 31078
rect 34336 30184 34388 30190
rect 34336 30126 34388 30132
rect 33692 29844 33744 29850
rect 33692 29786 33744 29792
rect 34060 29776 34112 29782
rect 34060 29718 34112 29724
rect 33416 29708 33468 29714
rect 33416 29650 33468 29656
rect 33048 29640 33100 29646
rect 33048 29582 33100 29588
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 33152 28082 33180 29242
rect 33140 28076 33192 28082
rect 33140 28018 33192 28024
rect 31760 28008 31812 28014
rect 31760 27950 31812 27956
rect 32404 28008 32456 28014
rect 32404 27950 32456 27956
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 27436 27056 27488 27062
rect 27436 26998 27488 27004
rect 27528 27056 27580 27062
rect 27528 26998 27580 27004
rect 31208 27056 31260 27062
rect 31208 26998 31260 27004
rect 27448 26518 27476 26998
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27540 26330 27568 26998
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 27356 26314 27568 26330
rect 27344 26308 27568 26314
rect 27396 26302 27568 26308
rect 27344 26250 27396 26256
rect 29472 25974 29500 26726
rect 30470 26480 30526 26489
rect 30470 26415 30472 26424
rect 30524 26415 30526 26424
rect 30472 26386 30524 26392
rect 30484 26042 30512 26386
rect 31220 26314 31248 26998
rect 31312 26586 31340 27406
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31496 27062 31524 27270
rect 31484 27056 31536 27062
rect 31484 26998 31536 27004
rect 31772 26994 31800 27950
rect 33232 27600 33284 27606
rect 33232 27542 33284 27548
rect 33244 27334 33272 27542
rect 31944 27328 31996 27334
rect 31944 27270 31996 27276
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 31760 26988 31812 26994
rect 31760 26930 31812 26936
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 30656 26240 30708 26246
rect 30656 26182 30708 26188
rect 30472 26036 30524 26042
rect 30472 25978 30524 25984
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27252 25832 27304 25838
rect 27252 25774 27304 25780
rect 27540 25702 27568 25842
rect 27068 25696 27120 25702
rect 27068 25638 27120 25644
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27080 25226 27108 25638
rect 27540 25498 27568 25638
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 30484 25294 30512 25978
rect 30668 25702 30696 26182
rect 31220 25974 31248 26250
rect 31208 25968 31260 25974
rect 31208 25910 31260 25916
rect 30656 25696 30708 25702
rect 30656 25638 30708 25644
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30472 25288 30524 25294
rect 30472 25230 30524 25236
rect 27068 25220 27120 25226
rect 27068 25162 27120 25168
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24964 23866 24992 24754
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25056 23798 25084 24686
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23322 24900 23462
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 24596 22778 24624 22986
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24780 22642 24808 22918
rect 24964 22778 24992 23666
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 25056 22642 25084 23734
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25148 22982 25176 23598
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25240 23118 25268 23462
rect 25424 23322 25452 23734
rect 25976 23730 26004 24142
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25424 23118 25452 23258
rect 25608 23118 25636 23598
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24872 22234 24900 22578
rect 25148 22574 25176 22918
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 25044 21412 25096 21418
rect 25044 21354 25096 21360
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24964 19854 24992 20742
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24228 18630 24256 19314
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24320 18766 24348 19110
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24412 18290 24440 19314
rect 25056 18766 25084 21354
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24308 18148 24360 18154
rect 24308 18090 24360 18096
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24228 14890 24256 17138
rect 24320 15502 24348 18090
rect 24412 17882 24440 18226
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24596 17678 24624 18702
rect 25056 17678 25084 18702
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24596 16726 24624 17614
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 24584 16720 24636 16726
rect 24584 16662 24636 16668
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 24964 16046 24992 16526
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 25056 15978 25084 17138
rect 25148 16794 25176 22510
rect 25608 22030 25636 23054
rect 25976 22166 26004 23666
rect 26148 23588 26200 23594
rect 26148 23530 26200 23536
rect 26160 23118 26188 23530
rect 26436 23186 26464 24142
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 26160 22710 26188 23054
rect 26148 22704 26200 22710
rect 26148 22646 26200 22652
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 25964 22160 26016 22166
rect 25964 22102 26016 22108
rect 26988 22098 27016 22510
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 21690 25636 21966
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25700 21554 25728 22034
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25700 21010 25728 21490
rect 25792 21146 25820 21966
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 25976 20942 26004 21286
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 25608 20466 25636 20810
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20466 25728 20742
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25412 19984 25464 19990
rect 25412 19926 25464 19932
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25332 19378 25360 19722
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25424 19310 25452 19926
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25608 18630 25636 20402
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25412 17808 25464 17814
rect 25412 17750 25464 17756
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25424 16590 25452 17750
rect 25516 17678 25544 18022
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25332 16250 25360 16390
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25424 16182 25452 16390
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25516 16114 25544 17614
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 25700 15638 25728 19314
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18766 25820 19110
rect 25976 18970 26004 20878
rect 26068 20874 26096 21422
rect 26056 20868 26108 20874
rect 26056 20810 26108 20816
rect 26068 20058 26096 20810
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25792 18290 25820 18702
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25976 18154 26004 18702
rect 25964 18148 26016 18154
rect 25964 18090 26016 18096
rect 26528 17678 26556 21898
rect 26988 20602 27016 22034
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 26620 19514 26648 19790
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 25884 16726 25912 17614
rect 25976 16998 26004 17614
rect 26056 17536 26108 17542
rect 26056 17478 26108 17484
rect 26068 17202 26096 17478
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25872 16720 25924 16726
rect 25872 16662 25924 16668
rect 25884 16114 25912 16662
rect 25976 16182 26004 16934
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 26528 15910 26556 17614
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 25688 15632 25740 15638
rect 25688 15574 25740 15580
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 24320 15026 24348 15438
rect 25608 15162 25636 15438
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24216 14884 24268 14890
rect 24216 14826 24268 14832
rect 24228 14414 24256 14826
rect 25608 14414 25636 15098
rect 26160 14958 26188 15370
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 26160 14618 26188 14894
rect 26436 14890 26464 15438
rect 26896 15434 26924 15506
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25424 14006 25452 14214
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23860 12850 23888 13670
rect 24320 12850 24348 13806
rect 24412 13326 24440 13874
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24688 13190 24716 13942
rect 25504 13932 25556 13938
rect 25780 13932 25832 13938
rect 25556 13892 25780 13920
rect 25504 13874 25556 13880
rect 25780 13874 25832 13880
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 24768 13796 24820 13802
rect 24768 13738 24820 13744
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24780 12434 24808 13738
rect 25148 13394 25176 13806
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 26252 13326 26280 13670
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26332 13320 26384 13326
rect 26436 13274 26464 14826
rect 26896 14618 26924 15370
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26988 15026 27016 15302
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26804 13462 26832 13806
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26384 13268 26464 13274
rect 26332 13262 26464 13268
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24780 12406 24900 12434
rect 24872 12306 24900 12406
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11354 24900 12242
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22296 2446 22324 7142
rect 24964 6934 24992 12582
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25240 11694 25268 12174
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 25424 2446 25452 13126
rect 25884 12986 25912 13262
rect 26252 13002 26280 13262
rect 26160 12986 26280 13002
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 26148 12980 26280 12986
rect 26200 12974 26280 12980
rect 26344 13246 26464 13262
rect 26148 12922 26200 12928
rect 26344 12646 26372 13246
rect 26896 13190 26924 14554
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 26436 12918 26464 13126
rect 26424 12912 26476 12918
rect 26424 12854 26476 12860
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25516 11762 25544 12038
rect 25700 11898 25728 12174
rect 26160 11898 26188 12174
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26252 11286 26280 11630
rect 26240 11280 26292 11286
rect 26240 11222 26292 11228
rect 26436 10470 26464 12854
rect 27080 10674 27108 25162
rect 28356 25152 28408 25158
rect 28356 25094 28408 25100
rect 28264 24200 28316 24206
rect 27434 24168 27490 24177
rect 28264 24142 28316 24148
rect 27434 24103 27436 24112
rect 27488 24103 27490 24112
rect 27436 24074 27488 24080
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 27252 23588 27304 23594
rect 27252 23530 27304 23536
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27172 22642 27200 23122
rect 27264 22778 27292 23530
rect 27816 23118 27844 24006
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27908 23186 27936 23734
rect 28000 23730 28028 24006
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 28276 23662 28304 24142
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27908 22778 27936 23122
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 27172 22030 27200 22578
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 28184 21690 28212 22578
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 28172 21684 28224 21690
rect 28172 21626 28224 21632
rect 27908 21350 27936 21626
rect 28368 21554 28396 25094
rect 30484 24954 30512 25230
rect 30472 24948 30524 24954
rect 30472 24890 30524 24896
rect 28448 24608 28500 24614
rect 28448 24550 28500 24556
rect 28460 24138 28488 24550
rect 29000 24268 29052 24274
rect 29000 24210 29052 24216
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 28460 23798 28488 24074
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28920 23186 28948 23666
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 29012 23118 29040 24210
rect 29092 24200 29144 24206
rect 29092 24142 29144 24148
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 29104 23866 29132 24142
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 30116 23798 30144 24142
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30300 23118 30328 23666
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30576 23186 30604 23462
rect 30564 23180 30616 23186
rect 30564 23122 30616 23128
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 29012 22710 29040 23054
rect 29000 22704 29052 22710
rect 29000 22646 29052 22652
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29276 22500 29328 22506
rect 29276 22442 29328 22448
rect 29288 22098 29316 22442
rect 29276 22092 29328 22098
rect 29276 22034 29328 22040
rect 29840 21622 29868 22510
rect 30668 22030 30696 25638
rect 30944 25430 30972 25638
rect 30932 25424 30984 25430
rect 30932 25366 30984 25372
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31404 25129 31432 25162
rect 31390 25120 31446 25129
rect 31390 25055 31446 25064
rect 30748 24268 30800 24274
rect 30748 24210 30800 24216
rect 30760 23594 30788 24210
rect 31668 24200 31720 24206
rect 31668 24142 31720 24148
rect 30748 23588 30800 23594
rect 30748 23530 30800 23536
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27264 20058 27292 20402
rect 27540 20330 27568 20742
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27632 19446 27660 19722
rect 27620 19440 27672 19446
rect 27620 19382 27672 19388
rect 27632 18970 27660 19382
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27264 17066 27292 18022
rect 27540 17882 27568 18226
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27264 16658 27292 17002
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27448 16454 27476 16594
rect 27632 16590 27660 17070
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27448 16114 27476 16390
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27264 15094 27292 15438
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27172 13326 27200 14894
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27264 13394 27292 13874
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27264 12918 27292 13194
rect 27540 13190 27568 14554
rect 27632 14550 27660 16526
rect 27724 14618 27752 21014
rect 27908 20874 27936 21286
rect 28368 21078 28396 21490
rect 30484 21486 30512 21830
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28356 21072 28408 21078
rect 28356 21014 28408 21020
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27908 20466 27936 20810
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27908 19922 27936 20402
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27908 19378 27936 19858
rect 28276 19854 28304 19994
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27816 18222 27844 18838
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27804 17604 27856 17610
rect 27908 17592 27936 19314
rect 28080 18692 28132 18698
rect 28080 18634 28132 18640
rect 28092 17814 28120 18634
rect 28080 17808 28132 17814
rect 28080 17750 28132 17756
rect 27856 17564 27936 17592
rect 27804 17546 27856 17552
rect 27816 15858 27844 17546
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27908 15978 27936 16526
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27816 15830 27936 15858
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 27816 14074 27844 14894
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27908 13954 27936 15830
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28000 14618 28028 14962
rect 28276 14929 28304 19790
rect 28736 19310 28764 20334
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28460 18834 28488 19110
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28736 18222 28764 19246
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28736 17610 28764 18158
rect 28724 17604 28776 17610
rect 28724 17546 28776 17552
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28368 16522 28396 16730
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28368 16250 28396 16458
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 28262 14920 28318 14929
rect 28172 14884 28224 14890
rect 28262 14855 28318 14864
rect 28172 14826 28224 14832
rect 27988 14612 28040 14618
rect 27988 14554 28040 14560
rect 27724 13926 27936 13954
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27540 12918 27568 13126
rect 27252 12912 27304 12918
rect 27252 12854 27304 12860
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27264 12306 27292 12854
rect 27540 12434 27568 12854
rect 27448 12406 27568 12434
rect 27252 12300 27304 12306
rect 27252 12242 27304 12248
rect 27448 12170 27476 12406
rect 27724 12238 27752 13926
rect 28000 13870 28028 14554
rect 28184 14482 28212 14826
rect 28172 14476 28224 14482
rect 28172 14418 28224 14424
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27908 12646 27936 13330
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 27896 12640 27948 12646
rect 27896 12582 27948 12588
rect 27908 12306 27936 12582
rect 27896 12300 27948 12306
rect 27896 12242 27948 12248
rect 28368 12238 28396 12786
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 27436 12164 27488 12170
rect 27436 12106 27488 12112
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27356 11898 27384 12038
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27448 11354 27476 12106
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27540 11762 27568 12038
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27724 10742 27752 12174
rect 28460 11558 28488 17478
rect 28540 16584 28592 16590
rect 28540 16526 28592 16532
rect 28552 16250 28580 16526
rect 28540 16244 28592 16250
rect 28540 16186 28592 16192
rect 28552 15706 28580 16186
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28644 15910 28672 16118
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28828 15502 28856 15982
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28540 13932 28592 13938
rect 28540 13874 28592 13880
rect 28552 13530 28580 13874
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28540 13184 28592 13190
rect 28540 13126 28592 13132
rect 28552 12782 28580 13126
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28552 12442 28580 12718
rect 28540 12436 28592 12442
rect 28540 12378 28592 12384
rect 28828 11898 28856 15438
rect 28920 15026 28948 21286
rect 29104 19922 29132 21422
rect 30196 20868 30248 20874
rect 30196 20810 30248 20816
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29748 20398 29776 20742
rect 30208 20466 30236 20810
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 29748 19854 29776 20198
rect 29736 19848 29788 19854
rect 29656 19796 29736 19802
rect 29656 19790 29788 19796
rect 29656 19774 29776 19790
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29196 16794 29224 17138
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29472 16114 29500 17546
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29104 15502 29132 16050
rect 29368 15972 29420 15978
rect 29368 15914 29420 15920
rect 29184 15904 29236 15910
rect 29236 15864 29316 15892
rect 29184 15846 29236 15852
rect 29288 15706 29316 15864
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29012 15094 29040 15302
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 28920 14414 28948 14962
rect 29012 14482 29040 15030
rect 29196 14618 29224 15098
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 28908 14408 28960 14414
rect 28908 14350 28960 14356
rect 29196 14346 29224 14554
rect 29184 14340 29236 14346
rect 29184 14282 29236 14288
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 29012 12442 29040 12786
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 29012 12238 29040 12378
rect 29104 12306 29132 12854
rect 29196 12850 29224 13942
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 29104 11830 29132 12242
rect 29092 11824 29144 11830
rect 29092 11766 29144 11772
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 29012 11286 29040 11698
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 29196 11218 29224 11630
rect 29288 11354 29316 15642
rect 29380 15570 29408 15914
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29472 13326 29500 16050
rect 29656 15434 29684 19774
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29748 17882 29776 19654
rect 29932 19378 29960 20402
rect 30208 19514 30236 20402
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30300 19854 30328 20198
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30392 19718 30420 20402
rect 30668 19938 30696 21966
rect 30760 20058 30788 23530
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 30840 22500 30892 22506
rect 30840 22442 30892 22448
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30484 19910 30696 19938
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29932 18290 29960 19314
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29932 17678 29960 18226
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29932 16114 29960 17614
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29644 15428 29696 15434
rect 29644 15370 29696 15376
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29656 14074 29684 14758
rect 30024 14618 30052 18022
rect 30208 17814 30236 18022
rect 30196 17808 30248 17814
rect 30196 17750 30248 17756
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30116 16182 30144 17138
rect 30104 16176 30156 16182
rect 30104 16118 30156 16124
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29460 13320 29512 13326
rect 29460 13262 29512 13268
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29932 11150 29960 12582
rect 30024 12442 30052 12650
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28736 10742 28764 10950
rect 27712 10736 27764 10742
rect 27712 10678 27764 10684
rect 28724 10736 28776 10742
rect 28724 10678 28776 10684
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26436 8974 26464 10406
rect 27080 10266 27108 10610
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27080 9586 27108 10202
rect 28736 9926 28764 10678
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29104 10266 29132 10542
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29748 10062 29776 11086
rect 29932 10198 29960 11086
rect 30024 10742 30052 11766
rect 30012 10736 30064 10742
rect 30012 10678 30064 10684
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 28724 9920 28776 9926
rect 28724 9862 28776 9868
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 27080 8634 27108 9522
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27448 9178 27476 9454
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27908 8974 27936 9862
rect 28736 9654 28764 9862
rect 28920 9722 28948 9998
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 28736 9178 28764 9590
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 27172 8430 27200 8910
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27356 8362 27384 8842
rect 27344 8356 27396 8362
rect 27344 8298 27396 8304
rect 27356 2582 27384 8298
rect 28184 8090 28212 9114
rect 30024 8974 30052 9318
rect 30012 8968 30064 8974
rect 30012 8910 30064 8916
rect 30116 8430 30144 16118
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30208 12782 30236 13262
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30208 12442 30236 12718
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 30300 10266 30328 15098
rect 30392 13802 30420 16050
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 30484 13530 30512 19910
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30576 19174 30604 19790
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30576 18358 30604 19110
rect 30564 18352 30616 18358
rect 30564 18294 30616 18300
rect 30576 15094 30604 18294
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 30668 15434 30696 15506
rect 30656 15428 30708 15434
rect 30656 15370 30708 15376
rect 30564 15088 30616 15094
rect 30564 15030 30616 15036
rect 30576 14414 30604 15030
rect 30668 15026 30696 15370
rect 30656 15020 30708 15026
rect 30656 14962 30708 14968
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30576 13938 30604 14350
rect 30852 14074 30880 22442
rect 31404 22438 31432 23054
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31392 22432 31444 22438
rect 31392 22374 31444 22380
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21690 31064 21966
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31220 21554 31248 22374
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31220 21146 31248 21490
rect 31208 21140 31260 21146
rect 31208 21082 31260 21088
rect 31404 19242 31432 22374
rect 31484 22024 31536 22030
rect 31484 21966 31536 21972
rect 31496 21554 31524 21966
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31680 20913 31708 24142
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31772 23118 31800 23598
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31666 20904 31722 20913
rect 31666 20839 31722 20848
rect 31392 19236 31444 19242
rect 31392 19178 31444 19184
rect 31404 18766 31432 19178
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 31392 18760 31444 18766
rect 31392 18702 31444 18708
rect 31036 15366 31064 18702
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 31128 18358 31156 18566
rect 31116 18352 31168 18358
rect 31116 18294 31168 18300
rect 31404 18170 31432 18702
rect 31312 18142 31432 18170
rect 31116 17536 31168 17542
rect 31116 17478 31168 17484
rect 31128 16114 31156 17478
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31312 15162 31340 18142
rect 31392 18080 31444 18086
rect 31392 18022 31444 18028
rect 31404 17678 31432 18022
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31404 17270 31432 17478
rect 31392 17264 31444 17270
rect 31392 17206 31444 17212
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31404 14618 31432 16050
rect 31588 15706 31616 16526
rect 31576 15700 31628 15706
rect 31576 15642 31628 15648
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31208 14476 31260 14482
rect 31208 14418 31260 14424
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30392 12170 30420 13262
rect 30484 13138 30512 13466
rect 30576 13258 30604 13874
rect 30656 13796 30708 13802
rect 30656 13738 30708 13744
rect 30564 13252 30616 13258
rect 30564 13194 30616 13200
rect 30484 13110 30604 13138
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30392 11898 30420 12106
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30484 11762 30512 12922
rect 30576 12918 30604 13110
rect 30668 12918 30696 13738
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 30564 12912 30616 12918
rect 30564 12854 30616 12860
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30576 11354 30604 12854
rect 30760 12850 30788 13262
rect 30852 13190 30880 14010
rect 31036 13530 31064 14214
rect 31220 14113 31248 14418
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31206 14104 31262 14113
rect 31206 14039 31208 14048
rect 31260 14039 31262 14048
rect 31208 14010 31260 14016
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31300 13932 31352 13938
rect 31300 13874 31352 13880
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 31024 13388 31076 13394
rect 31024 13330 31076 13336
rect 30932 13252 30984 13258
rect 30932 13194 30984 13200
rect 30840 13184 30892 13190
rect 30840 13126 30892 13132
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30852 12782 30880 13126
rect 30840 12776 30892 12782
rect 30840 12718 30892 12724
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30668 11626 30696 12174
rect 30944 12102 30972 13194
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 30656 11620 30708 11626
rect 30656 11562 30708 11568
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30392 8634 30420 9590
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30576 9178 30604 9454
rect 30564 9172 30616 9178
rect 30564 9114 30616 9120
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30484 8498 30512 8774
rect 30576 8566 30604 9114
rect 30668 9110 30696 11562
rect 31036 10742 31064 13330
rect 31128 12918 31156 13874
rect 31312 13326 31340 13874
rect 31300 13320 31352 13326
rect 31300 13262 31352 13268
rect 31312 12918 31340 13262
rect 31116 12912 31168 12918
rect 31116 12854 31168 12860
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31128 11762 31156 12854
rect 31588 12850 31616 14350
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31392 12776 31444 12782
rect 31392 12718 31444 12724
rect 31300 12640 31352 12646
rect 31300 12582 31352 12588
rect 31312 12238 31340 12582
rect 31300 12232 31352 12238
rect 31208 12210 31260 12216
rect 31300 12174 31352 12180
rect 31404 12220 31432 12718
rect 31484 12232 31536 12238
rect 31404 12192 31484 12220
rect 31208 12152 31260 12158
rect 31220 11898 31248 12152
rect 31404 11898 31432 12192
rect 31484 12174 31536 12180
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31392 11892 31444 11898
rect 31392 11834 31444 11840
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 31024 10736 31076 10742
rect 30944 10696 31024 10724
rect 30944 9518 30972 10696
rect 31024 10678 31076 10684
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 31036 9586 31064 10066
rect 31312 10062 31340 10678
rect 31300 10056 31352 10062
rect 31300 9998 31352 10004
rect 31312 9654 31340 9998
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 30932 9512 30984 9518
rect 30932 9454 30984 9460
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30564 8560 30616 8566
rect 30564 8502 30616 8508
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 30668 8362 30696 9046
rect 31036 9042 31064 9522
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31128 9178 31156 9318
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 31024 9036 31076 9042
rect 31024 8978 31076 8984
rect 31220 8974 31248 9454
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 31404 8634 31432 9318
rect 31496 8906 31524 12038
rect 31588 11762 31616 12786
rect 31576 11756 31628 11762
rect 31576 11698 31628 11704
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30668 8090 30696 8298
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 31036 7954 31064 8434
rect 31024 7948 31076 7954
rect 31024 7890 31076 7896
rect 31220 7886 31248 8434
rect 31404 8022 31432 8570
rect 31496 8498 31524 8842
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 31392 8016 31444 8022
rect 31392 7958 31444 7964
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31220 7342 31248 7822
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7410 31432 7686
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 27712 6928 27764 6934
rect 27712 6870 27764 6876
rect 27344 2576 27396 2582
rect 27344 2518 27396 2524
rect 27724 2446 27752 6870
rect 31680 2650 31708 20839
rect 31772 18834 31800 23054
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31864 22030 31892 22578
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 31864 21418 31892 21966
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31956 20890 31984 27270
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33244 26382 33272 26726
rect 33428 26586 33456 29650
rect 34072 29238 34100 29718
rect 34060 29232 34112 29238
rect 34060 29174 34112 29180
rect 33784 29096 33836 29102
rect 33598 29064 33654 29073
rect 33784 29038 33836 29044
rect 33598 28999 33654 29008
rect 33612 28490 33640 28999
rect 33796 28558 33824 29038
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 33600 28484 33652 28490
rect 33600 28426 33652 28432
rect 33612 28082 33640 28426
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33796 26994 33824 27270
rect 33980 26994 34008 28494
rect 34716 28150 34744 36178
rect 34808 35698 34836 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34888 36168 34940 36174
rect 34888 36110 34940 36116
rect 35256 36168 35308 36174
rect 35256 36110 35308 36116
rect 34900 35834 34928 36110
rect 35164 36032 35216 36038
rect 35164 35974 35216 35980
rect 34888 35828 34940 35834
rect 34888 35770 34940 35776
rect 35176 35698 35204 35974
rect 35268 35698 35296 36110
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 35164 35692 35216 35698
rect 35164 35634 35216 35640
rect 35256 35692 35308 35698
rect 35256 35634 35308 35640
rect 34808 35154 34836 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 35148 34848 35154
rect 34796 35090 34848 35096
rect 35636 34932 35664 56646
rect 35900 45280 35952 45286
rect 35900 45222 35952 45228
rect 35808 43648 35860 43654
rect 35808 43590 35860 43596
rect 35820 42770 35848 43590
rect 35808 42764 35860 42770
rect 35808 42706 35860 42712
rect 35820 42566 35848 42706
rect 35808 42560 35860 42566
rect 35808 42502 35860 42508
rect 35912 41614 35940 45222
rect 35992 43172 36044 43178
rect 35992 43114 36044 43120
rect 35900 41608 35952 41614
rect 35900 41550 35952 41556
rect 35716 41472 35768 41478
rect 35716 41414 35768 41420
rect 35728 40118 35756 41414
rect 35808 40384 35860 40390
rect 35808 40326 35860 40332
rect 35900 40384 35952 40390
rect 35900 40326 35952 40332
rect 35716 40112 35768 40118
rect 35716 40054 35768 40060
rect 35820 40050 35848 40326
rect 35808 40044 35860 40050
rect 35808 39986 35860 39992
rect 35716 39840 35768 39846
rect 35716 39782 35768 39788
rect 35728 39506 35756 39782
rect 35716 39500 35768 39506
rect 35716 39442 35768 39448
rect 35820 39302 35848 39986
rect 35912 39982 35940 40326
rect 35900 39976 35952 39982
rect 35900 39918 35952 39924
rect 35912 39506 35940 39918
rect 35900 39500 35952 39506
rect 35900 39442 35952 39448
rect 35808 39296 35860 39302
rect 35808 39238 35860 39244
rect 36004 37670 36032 43114
rect 37096 42560 37148 42566
rect 37096 42502 37148 42508
rect 36084 39840 36136 39846
rect 36084 39782 36136 39788
rect 36096 39506 36124 39782
rect 36084 39500 36136 39506
rect 36084 39442 36136 39448
rect 36176 39296 36228 39302
rect 36176 39238 36228 39244
rect 36188 38758 36216 39238
rect 36360 39024 36412 39030
rect 36360 38966 36412 38972
rect 36176 38752 36228 38758
rect 36176 38694 36228 38700
rect 36188 38282 36216 38694
rect 36176 38276 36228 38282
rect 36176 38218 36228 38224
rect 35992 37664 36044 37670
rect 35992 37606 36044 37612
rect 36004 35630 36032 37606
rect 36188 37126 36216 38218
rect 36176 37120 36228 37126
rect 36176 37062 36228 37068
rect 36188 36854 36216 37062
rect 36176 36848 36228 36854
rect 36176 36790 36228 36796
rect 36188 36038 36216 36790
rect 36372 36718 36400 38966
rect 37108 38282 37136 42502
rect 37464 41472 37516 41478
rect 37464 41414 37516 41420
rect 37476 39506 37504 41414
rect 37464 39500 37516 39506
rect 37464 39442 37516 39448
rect 37096 38276 37148 38282
rect 37096 38218 37148 38224
rect 36360 36712 36412 36718
rect 36360 36654 36412 36660
rect 36176 36032 36228 36038
rect 36176 35974 36228 35980
rect 36188 35766 36216 35974
rect 36176 35760 36228 35766
rect 36176 35702 36228 35708
rect 35992 35624 36044 35630
rect 35992 35566 36044 35572
rect 35452 34904 35664 34932
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34980 34060 35032 34066
rect 34980 34002 35032 34008
rect 34992 33658 35020 34002
rect 34980 33652 35032 33658
rect 34980 33594 35032 33600
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35452 32026 35480 34904
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35716 34604 35768 34610
rect 35716 34546 35768 34552
rect 35544 34202 35572 34546
rect 35624 34400 35676 34406
rect 35624 34342 35676 34348
rect 35532 34196 35584 34202
rect 35532 34138 35584 34144
rect 35636 33522 35664 34342
rect 35728 33998 35756 34546
rect 35716 33992 35768 33998
rect 35716 33934 35768 33940
rect 35808 33856 35860 33862
rect 35808 33798 35860 33804
rect 35820 33522 35848 33798
rect 35624 33516 35676 33522
rect 35624 33458 35676 33464
rect 35808 33516 35860 33522
rect 35808 33458 35860 33464
rect 35532 33448 35584 33454
rect 35532 33390 35584 33396
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35348 31340 35400 31346
rect 35348 31282 35400 31288
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 34808 30394 34836 31214
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30938 35388 31282
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 35452 30326 35480 31758
rect 35440 30320 35492 30326
rect 35440 30262 35492 30268
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35544 29102 35572 33390
rect 35716 33312 35768 33318
rect 35716 33254 35768 33260
rect 35624 32768 35676 32774
rect 35624 32710 35676 32716
rect 35636 31822 35664 32710
rect 35728 32434 35756 33254
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 35820 32230 35848 32846
rect 36004 32570 36032 32846
rect 35992 32564 36044 32570
rect 35992 32506 36044 32512
rect 35808 32224 35860 32230
rect 35808 32166 35860 32172
rect 35624 31816 35676 31822
rect 35676 31776 35756 31804
rect 35624 31758 35676 31764
rect 35728 30734 35756 31776
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35716 30728 35768 30734
rect 35716 30670 35768 30676
rect 35912 30598 35940 31282
rect 35992 31136 36044 31142
rect 35992 31078 36044 31084
rect 36004 30734 36032 31078
rect 36084 30796 36136 30802
rect 36084 30738 36136 30744
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 35900 30592 35952 30598
rect 35900 30534 35952 30540
rect 35912 30258 35940 30534
rect 36004 30326 36032 30670
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 36096 30258 36124 30738
rect 35900 30252 35952 30258
rect 35900 30194 35952 30200
rect 36084 30252 36136 30258
rect 36084 30194 36136 30200
rect 36096 30122 36124 30194
rect 36084 30116 36136 30122
rect 36084 30058 36136 30064
rect 36096 29170 36124 30058
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 35532 29096 35584 29102
rect 35532 29038 35584 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35532 28484 35584 28490
rect 35532 28426 35584 28432
rect 34152 28144 34204 28150
rect 34152 28086 34204 28092
rect 34704 28144 34756 28150
rect 34704 28086 34756 28092
rect 33784 26988 33836 26994
rect 33784 26930 33836 26936
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 33796 26858 33824 26930
rect 33784 26852 33836 26858
rect 33784 26794 33836 26800
rect 33416 26580 33468 26586
rect 33416 26522 33468 26528
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 32588 26308 32640 26314
rect 32640 26268 32720 26296
rect 32588 26250 32640 26256
rect 32692 25226 32720 26268
rect 33428 26042 33456 26522
rect 33980 26450 34008 26930
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 33876 26240 33928 26246
rect 33876 26182 33928 26188
rect 33888 26042 33916 26182
rect 33416 26036 33468 26042
rect 33416 25978 33468 25984
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 33428 25838 33456 25978
rect 33600 25900 33652 25906
rect 33600 25842 33652 25848
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25362 33180 25638
rect 33428 25378 33456 25774
rect 33612 25498 33640 25842
rect 33600 25492 33652 25498
rect 33600 25434 33652 25440
rect 33876 25492 33928 25498
rect 33876 25434 33928 25440
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 33336 25350 33456 25378
rect 32680 25220 32732 25226
rect 32680 25162 32732 25168
rect 32588 24132 32640 24138
rect 32692 24120 32720 25162
rect 33336 24818 33364 25350
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 33428 24206 33456 25230
rect 33888 24834 33916 25434
rect 33980 25430 34008 26386
rect 33968 25424 34020 25430
rect 33968 25366 34020 25372
rect 34072 25226 34100 26794
rect 34060 25220 34112 25226
rect 34060 25162 34112 25168
rect 34072 24954 34100 25162
rect 34060 24948 34112 24954
rect 33980 24886 34008 24917
rect 34060 24890 34112 24896
rect 33968 24880 34020 24886
rect 33888 24828 33968 24834
rect 33888 24822 34020 24828
rect 33888 24806 34008 24822
rect 33876 24744 33928 24750
rect 33876 24686 33928 24692
rect 33600 24608 33652 24614
rect 33600 24550 33652 24556
rect 33416 24200 33468 24206
rect 33416 24142 33468 24148
rect 32640 24092 32720 24120
rect 32588 24074 32640 24080
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 32232 22642 32260 24006
rect 32956 23724 33008 23730
rect 32956 23666 33008 23672
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 32404 23180 32456 23186
rect 32404 23122 32456 23128
rect 32416 22778 32444 23122
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 32784 22778 32812 22918
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32772 22772 32824 22778
rect 32772 22714 32824 22720
rect 32312 22704 32364 22710
rect 32312 22646 32364 22652
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32232 20942 32260 21490
rect 32324 21418 32352 22646
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 32600 22234 32628 22578
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32600 21962 32628 22170
rect 32588 21956 32640 21962
rect 32588 21898 32640 21904
rect 32586 21720 32642 21729
rect 32586 21655 32642 21664
rect 32600 21622 32628 21655
rect 32588 21616 32640 21622
rect 32588 21558 32640 21564
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32312 21412 32364 21418
rect 32312 21354 32364 21360
rect 32416 21146 32444 21490
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 32784 21146 32812 21422
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32772 21140 32824 21146
rect 32772 21082 32824 21088
rect 31864 20862 31984 20890
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 31864 20806 31892 20862
rect 31852 20800 31904 20806
rect 31852 20742 31904 20748
rect 32404 20800 32456 20806
rect 32404 20742 32456 20748
rect 31864 20330 31892 20742
rect 31852 20324 31904 20330
rect 31852 20266 31904 20272
rect 31864 19718 31892 20266
rect 31852 19712 31904 19718
rect 31852 19654 31904 19660
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31864 17610 31892 19314
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 32048 18290 32076 18634
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31944 18148 31996 18154
rect 31944 18090 31996 18096
rect 31956 17746 31984 18090
rect 32140 17785 32168 18362
rect 32232 18222 32260 18702
rect 32220 18216 32272 18222
rect 32220 18158 32272 18164
rect 32126 17776 32182 17785
rect 31944 17740 31996 17746
rect 32126 17711 32182 17720
rect 31944 17682 31996 17688
rect 31852 17604 31904 17610
rect 31852 17546 31904 17552
rect 31864 14006 31892 17546
rect 31956 17338 31984 17682
rect 32140 17678 32168 17711
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 32416 16590 32444 20742
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 32508 20058 32536 20470
rect 32784 20466 32812 21082
rect 32968 20874 32996 23666
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 32956 20868 33008 20874
rect 32956 20810 33008 20816
rect 33060 20466 33088 22170
rect 33244 22098 33272 23054
rect 33416 22976 33468 22982
rect 33416 22918 33468 22924
rect 33428 22166 33456 22918
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 33232 22092 33284 22098
rect 33232 22034 33284 22040
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 32772 20460 32824 20466
rect 33048 20460 33100 20466
rect 32772 20402 32824 20408
rect 32968 20420 33048 20448
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 32864 19984 32916 19990
rect 32864 19926 32916 19932
rect 32876 19242 32904 19926
rect 32864 19236 32916 19242
rect 32864 19178 32916 19184
rect 32876 18873 32904 19178
rect 32862 18864 32918 18873
rect 32862 18799 32918 18808
rect 32680 18624 32732 18630
rect 32680 18566 32732 18572
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 31944 15904 31996 15910
rect 31944 15846 31996 15852
rect 31956 15502 31984 15846
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 32232 14958 32260 16526
rect 32508 16114 32536 18226
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32600 17202 32628 18022
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32508 15570 32536 16050
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32496 15564 32548 15570
rect 32496 15506 32548 15512
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 31852 14000 31904 14006
rect 31852 13942 31904 13948
rect 32508 13462 32536 15506
rect 32600 15502 32628 15846
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32600 15162 32628 15438
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32692 15026 32720 18566
rect 32968 18272 32996 20420
rect 33048 20402 33100 20408
rect 33152 20058 33180 21966
rect 33244 21894 33272 22034
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 33244 21010 33272 21830
rect 33336 21690 33364 21966
rect 33520 21729 33548 23666
rect 33612 23662 33640 24550
rect 33888 24274 33916 24686
rect 33980 24274 34008 24806
rect 33876 24268 33928 24274
rect 33876 24210 33928 24216
rect 33968 24268 34020 24274
rect 33968 24210 34020 24216
rect 33692 24200 33744 24206
rect 33692 24142 33744 24148
rect 33704 23730 33732 24142
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33612 22438 33640 23598
rect 33600 22432 33652 22438
rect 33600 22374 33652 22380
rect 33506 21720 33562 21729
rect 33324 21684 33376 21690
rect 33506 21655 33562 21664
rect 33324 21626 33376 21632
rect 33232 21004 33284 21010
rect 33232 20946 33284 20952
rect 33416 20256 33468 20262
rect 33416 20198 33468 20204
rect 33140 20052 33192 20058
rect 33140 19994 33192 20000
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33060 18970 33088 19790
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 33232 19440 33284 19446
rect 33232 19382 33284 19388
rect 33048 18964 33100 18970
rect 33048 18906 33100 18912
rect 33060 18766 33088 18906
rect 33048 18760 33100 18766
rect 33048 18702 33100 18708
rect 33244 18426 33272 19382
rect 33336 19378 33364 19654
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33336 19174 33364 19314
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33336 18698 33364 19110
rect 33324 18692 33376 18698
rect 33324 18634 33376 18640
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 33336 18290 33364 18634
rect 33324 18284 33376 18290
rect 32968 18244 33088 18272
rect 32956 18148 33008 18154
rect 32956 18090 33008 18096
rect 32968 17882 32996 18090
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 33060 17626 33088 18244
rect 33324 18226 33376 18232
rect 33428 17882 33456 20198
rect 33520 19854 33548 21655
rect 33600 20800 33652 20806
rect 33600 20742 33652 20748
rect 33508 19848 33560 19854
rect 33508 19790 33560 19796
rect 33612 18766 33640 20742
rect 33704 20346 33732 23666
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33796 23322 33824 23462
rect 33784 23316 33836 23322
rect 33784 23258 33836 23264
rect 34060 22772 34112 22778
rect 34060 22714 34112 22720
rect 33876 22432 33928 22438
rect 33876 22374 33928 22380
rect 33888 22137 33916 22374
rect 33874 22128 33930 22137
rect 33874 22063 33930 22072
rect 33876 21888 33928 21894
rect 33876 21830 33928 21836
rect 33888 20466 33916 21830
rect 34072 21690 34100 22714
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 33968 21548 34020 21554
rect 33968 21490 34020 21496
rect 33980 20942 34008 21490
rect 33968 20936 34020 20942
rect 33968 20878 34020 20884
rect 34060 20868 34112 20874
rect 34060 20810 34112 20816
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33704 20318 33916 20346
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33416 17876 33468 17882
rect 33416 17818 33468 17824
rect 33416 17672 33468 17678
rect 33230 17640 33286 17649
rect 33060 17598 33230 17626
rect 33416 17614 33468 17620
rect 33230 17575 33286 17584
rect 33244 17270 33272 17575
rect 33428 17338 33456 17614
rect 33416 17332 33468 17338
rect 33416 17274 33468 17280
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 32772 15088 32824 15094
rect 32772 15030 32824 15036
rect 32680 15020 32732 15026
rect 32680 14962 32732 14968
rect 32784 14890 32812 15030
rect 32968 14890 32996 17138
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 33336 16726 33364 16934
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 33336 16590 33364 16662
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 33324 16584 33376 16590
rect 33324 16526 33376 16532
rect 33060 15366 33088 16526
rect 33140 16108 33192 16114
rect 33140 16050 33192 16056
rect 33152 15570 33180 16050
rect 33232 15700 33284 15706
rect 33232 15642 33284 15648
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 33060 15162 33088 15302
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32772 14884 32824 14890
rect 32956 14884 33008 14890
rect 32824 14844 32904 14872
rect 32772 14826 32824 14832
rect 32772 14340 32824 14346
rect 32772 14282 32824 14288
rect 32784 13530 32812 14282
rect 32876 13870 32904 14844
rect 32956 14826 33008 14832
rect 32956 14340 33008 14346
rect 32956 14282 33008 14288
rect 32968 14074 32996 14282
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 33060 13938 33088 14962
rect 33140 14952 33192 14958
rect 33140 14894 33192 14900
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32496 13456 32548 13462
rect 32496 13398 32548 13404
rect 32876 13258 32904 13806
rect 33060 13530 33088 13874
rect 33152 13870 33180 14894
rect 33244 13938 33272 15642
rect 33336 15502 33364 16526
rect 33612 16250 33640 18702
rect 33600 16244 33652 16250
rect 33600 16186 33652 16192
rect 33704 16114 33732 20198
rect 33782 19952 33838 19961
rect 33782 19887 33838 19896
rect 33796 19854 33824 19887
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33888 19281 33916 20318
rect 34072 20262 34100 20810
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 34072 20058 34100 20198
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 33968 19780 34020 19786
rect 33968 19722 34020 19728
rect 34060 19780 34112 19786
rect 34060 19722 34112 19728
rect 33874 19272 33930 19281
rect 33874 19207 33930 19216
rect 33876 18080 33928 18086
rect 33876 18022 33928 18028
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33796 16794 33824 17478
rect 33784 16788 33836 16794
rect 33784 16730 33836 16736
rect 33692 16108 33744 16114
rect 33692 16050 33744 16056
rect 33888 15910 33916 18022
rect 33980 17218 34008 19722
rect 34072 18358 34100 19722
rect 34060 18352 34112 18358
rect 34060 18294 34112 18300
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 34072 17338 34100 17478
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 33980 17190 34100 17218
rect 33968 17128 34020 17134
rect 33968 17070 34020 17076
rect 33980 16998 34008 17070
rect 33968 16992 34020 16998
rect 33968 16934 34020 16940
rect 33980 16590 34008 16934
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 33876 15904 33928 15910
rect 33876 15846 33928 15852
rect 34072 15638 34100 17190
rect 34060 15632 34112 15638
rect 34060 15574 34112 15580
rect 33692 15564 33744 15570
rect 33692 15506 33744 15512
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33704 15162 33732 15506
rect 33968 15496 34020 15502
rect 33968 15438 34020 15444
rect 33692 15156 33744 15162
rect 33692 15098 33744 15104
rect 33980 14618 34008 15438
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33876 14272 33928 14278
rect 33876 14214 33928 14220
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33048 13524 33100 13530
rect 33048 13466 33100 13472
rect 32956 13456 33008 13462
rect 32956 13398 33008 13404
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32968 12850 32996 13398
rect 33060 13326 33088 13466
rect 33048 13320 33100 13326
rect 33048 13262 33100 13268
rect 33152 13190 33180 13806
rect 33232 13388 33284 13394
rect 33232 13330 33284 13336
rect 33140 13184 33192 13190
rect 33140 13126 33192 13132
rect 33152 12986 33180 13126
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 32588 12776 32640 12782
rect 32588 12718 32640 12724
rect 32600 12442 32628 12718
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 32036 12300 32088 12306
rect 32036 12242 32088 12248
rect 32048 12102 32076 12242
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 32692 11694 32720 12310
rect 32784 12238 32812 12378
rect 32772 12232 32824 12238
rect 32772 12174 32824 12180
rect 32784 11762 32812 12174
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32680 11688 32732 11694
rect 32680 11630 32732 11636
rect 32312 11212 32364 11218
rect 32312 11154 32364 11160
rect 32324 10810 32352 11154
rect 32968 11098 32996 12786
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 33060 11830 33088 12174
rect 33152 11898 33180 12310
rect 33140 11892 33192 11898
rect 33140 11834 33192 11840
rect 33048 11824 33100 11830
rect 33048 11766 33100 11772
rect 33244 11354 33272 13330
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33520 12306 33548 12922
rect 33796 12434 33824 13874
rect 33888 13734 33916 14214
rect 34072 13870 34100 14350
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33876 13728 33928 13734
rect 33876 13670 33928 13676
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33612 12406 33824 12434
rect 33508 12300 33560 12306
rect 33508 12242 33560 12248
rect 33612 12238 33640 12406
rect 33600 12232 33652 12238
rect 33600 12174 33652 12180
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33520 11898 33548 12106
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33888 11354 33916 12174
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 33876 11348 33928 11354
rect 33876 11290 33928 11296
rect 33244 11218 33272 11290
rect 33980 11218 34008 13330
rect 33232 11212 33284 11218
rect 33232 11154 33284 11160
rect 33968 11212 34020 11218
rect 33968 11154 34020 11160
rect 32968 11082 33088 11098
rect 32968 11076 33100 11082
rect 32968 11070 33048 11076
rect 33048 11018 33100 11024
rect 32496 11008 32548 11014
rect 32496 10950 32548 10956
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32508 10470 32536 10950
rect 33060 10674 33088 11018
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32508 9654 32536 10202
rect 33060 10062 33088 10610
rect 33244 10470 33272 11154
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33692 11144 33744 11150
rect 33692 11086 33744 11092
rect 33520 10674 33548 11086
rect 33704 10810 33732 11086
rect 33876 11076 33928 11082
rect 33876 11018 33928 11024
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 33244 10266 33272 10406
rect 33704 10266 33732 10746
rect 33232 10260 33284 10266
rect 33232 10202 33284 10208
rect 33692 10260 33744 10266
rect 33692 10202 33744 10208
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 33048 9648 33100 9654
rect 33048 9590 33100 9596
rect 32956 9444 33008 9450
rect 32956 9386 33008 9392
rect 32968 9194 32996 9386
rect 32876 9178 32996 9194
rect 32876 9172 33008 9178
rect 32876 9166 32956 9172
rect 32876 9058 32904 9166
rect 32956 9114 33008 9120
rect 32784 9042 32904 9058
rect 32772 9036 32904 9042
rect 32824 9030 32904 9036
rect 32772 8978 32824 8984
rect 32876 8566 32904 9030
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32864 8560 32916 8566
rect 32864 8502 32916 8508
rect 32968 8498 32996 8978
rect 33060 8906 33088 9590
rect 33704 9586 33732 9862
rect 33888 9586 33916 11018
rect 33980 10538 34008 11154
rect 33968 10532 34020 10538
rect 33968 10474 34020 10480
rect 33980 10062 34008 10474
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33704 9042 33732 9522
rect 33692 9036 33744 9042
rect 33692 8978 33744 8984
rect 33888 8974 33916 9522
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33048 8900 33100 8906
rect 33048 8842 33100 8848
rect 33876 8832 33928 8838
rect 33876 8774 33928 8780
rect 33888 8498 33916 8774
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 32956 8492 33008 8498
rect 32956 8434 33008 8440
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33232 8288 33284 8294
rect 33232 8230 33284 8236
rect 33244 7886 33272 8230
rect 33888 8090 33916 8434
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33140 7812 33192 7818
rect 33140 7754 33192 7760
rect 32956 7200 33008 7206
rect 32956 7142 33008 7148
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32968 2446 32996 7142
rect 33152 6798 33180 7754
rect 33244 6934 33272 7822
rect 33692 7404 33744 7410
rect 33692 7346 33744 7352
rect 33704 7002 33732 7346
rect 33796 7342 33824 7822
rect 33980 7818 34008 8366
rect 34072 7818 34100 8570
rect 33968 7812 34020 7818
rect 33968 7754 34020 7760
rect 34060 7812 34112 7818
rect 34060 7754 34112 7760
rect 33784 7336 33836 7342
rect 33784 7278 33836 7284
rect 33692 6996 33744 7002
rect 33692 6938 33744 6944
rect 33232 6928 33284 6934
rect 33232 6870 33284 6876
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 34164 2774 34192 28086
rect 34716 27418 34744 28086
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34624 27390 34744 27418
rect 34244 27328 34296 27334
rect 34244 27270 34296 27276
rect 34256 27062 34284 27270
rect 34624 27130 34652 27390
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34612 27124 34664 27130
rect 34612 27066 34664 27072
rect 34244 27056 34296 27062
rect 34244 26998 34296 27004
rect 34716 26994 34744 27270
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34808 26586 34836 28018
rect 35348 28008 35400 28014
rect 35348 27950 35400 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27402 35388 27950
rect 35440 27872 35492 27878
rect 35440 27814 35492 27820
rect 35452 27674 35480 27814
rect 35440 27668 35492 27674
rect 35440 27610 35492 27616
rect 35348 27396 35400 27402
rect 35348 27338 35400 27344
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26586 35388 27338
rect 35544 27130 35572 28426
rect 35624 28076 35676 28082
rect 35624 28018 35676 28024
rect 35532 27124 35584 27130
rect 35532 27066 35584 27072
rect 35636 27010 35664 28018
rect 35900 27464 35952 27470
rect 35900 27406 35952 27412
rect 35452 26994 35664 27010
rect 35440 26988 35664 26994
rect 35492 26982 35664 26988
rect 35440 26930 35492 26936
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 34336 26376 34388 26382
rect 34336 26318 34388 26324
rect 34244 25764 34296 25770
rect 34244 25706 34296 25712
rect 34256 25226 34284 25706
rect 34244 25220 34296 25226
rect 34244 25162 34296 25168
rect 34256 24614 34284 25162
rect 34348 24818 34376 26318
rect 34796 26308 34848 26314
rect 34796 26250 34848 26256
rect 34808 24818 34836 26250
rect 35452 26042 35480 26930
rect 35532 26920 35584 26926
rect 35532 26862 35584 26868
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 35544 25906 35572 26862
rect 35912 26790 35940 27406
rect 35900 26784 35952 26790
rect 35900 26726 35952 26732
rect 35912 26246 35940 26726
rect 36188 26586 36216 35702
rect 36912 34944 36964 34950
rect 36912 34886 36964 34892
rect 36728 34536 36780 34542
rect 36728 34478 36780 34484
rect 36636 33992 36688 33998
rect 36636 33934 36688 33940
rect 36648 33522 36676 33934
rect 36636 33516 36688 33522
rect 36636 33458 36688 33464
rect 36648 33046 36676 33458
rect 36740 33454 36768 34478
rect 36728 33448 36780 33454
rect 36728 33390 36780 33396
rect 36636 33040 36688 33046
rect 36636 32982 36688 32988
rect 36740 32842 36768 33390
rect 36820 33312 36872 33318
rect 36820 33254 36872 33260
rect 36832 32910 36860 33254
rect 36820 32904 36872 32910
rect 36820 32846 36872 32852
rect 36728 32836 36780 32842
rect 36728 32778 36780 32784
rect 36452 32292 36504 32298
rect 36452 32234 36504 32240
rect 36464 31890 36492 32234
rect 36452 31884 36504 31890
rect 36452 31826 36504 31832
rect 36464 30938 36492 31826
rect 36452 30932 36504 30938
rect 36452 30874 36504 30880
rect 36636 30252 36688 30258
rect 36636 30194 36688 30200
rect 36648 30122 36676 30194
rect 36636 30116 36688 30122
rect 36636 30058 36688 30064
rect 36544 28416 36596 28422
rect 36544 28358 36596 28364
rect 36452 27872 36504 27878
rect 36452 27814 36504 27820
rect 36464 27334 36492 27814
rect 36452 27328 36504 27334
rect 36452 27270 36504 27276
rect 36176 26580 36228 26586
rect 36176 26522 36228 26528
rect 36084 26308 36136 26314
rect 36084 26250 36136 26256
rect 35900 26240 35952 26246
rect 35900 26182 35952 26188
rect 35440 25900 35492 25906
rect 35440 25842 35492 25848
rect 35532 25900 35584 25906
rect 35532 25842 35584 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35452 25362 35480 25842
rect 35544 25430 35572 25842
rect 35808 25492 35860 25498
rect 35808 25434 35860 25440
rect 35532 25424 35584 25430
rect 35532 25366 35584 25372
rect 35440 25356 35492 25362
rect 35440 25298 35492 25304
rect 35256 25288 35308 25294
rect 35256 25230 35308 25236
rect 35268 24954 35296 25230
rect 35256 24948 35308 24954
rect 35256 24890 35308 24896
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34796 24812 34848 24818
rect 34796 24754 34848 24760
rect 34244 24608 34296 24614
rect 34244 24550 34296 24556
rect 34348 24410 34376 24754
rect 34336 24404 34388 24410
rect 34336 24346 34388 24352
rect 34532 24342 34560 24754
rect 34520 24336 34572 24342
rect 34572 24296 34652 24324
rect 34520 24278 34572 24284
rect 34336 23860 34388 23866
rect 34336 23802 34388 23808
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34256 23186 34284 23258
rect 34244 23180 34296 23186
rect 34244 23122 34296 23128
rect 34244 22772 34296 22778
rect 34244 22714 34296 22720
rect 34256 19854 34284 22714
rect 34348 20330 34376 23802
rect 34428 23520 34480 23526
rect 34428 23462 34480 23468
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34440 22642 34468 23462
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34532 22506 34560 23462
rect 34624 23118 34652 24296
rect 34704 23520 34756 23526
rect 34704 23462 34756 23468
rect 34612 23112 34664 23118
rect 34612 23054 34664 23060
rect 34624 22778 34652 23054
rect 34612 22772 34664 22778
rect 34612 22714 34664 22720
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34520 22500 34572 22506
rect 34520 22442 34572 22448
rect 34532 21962 34560 22442
rect 34624 22166 34652 22578
rect 34612 22160 34664 22166
rect 34612 22102 34664 22108
rect 34520 21956 34572 21962
rect 34520 21898 34572 21904
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 34336 20324 34388 20330
rect 34336 20266 34388 20272
rect 34244 19848 34296 19854
rect 34244 19790 34296 19796
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34336 19168 34388 19174
rect 34336 19110 34388 19116
rect 34348 18766 34376 19110
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34440 18290 34468 19314
rect 34532 19310 34560 21490
rect 34624 19344 34652 22102
rect 34716 22094 34744 23462
rect 34808 23202 34836 24754
rect 35348 24744 35400 24750
rect 35348 24686 35400 24692
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24426 35388 24686
rect 35268 24398 35388 24426
rect 35452 24426 35480 25298
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 35532 25152 35584 25158
rect 35532 25094 35584 25100
rect 35544 24750 35572 25094
rect 35532 24744 35584 24750
rect 35728 24698 35756 25162
rect 35532 24686 35584 24692
rect 35636 24682 35756 24698
rect 35624 24676 35756 24682
rect 35676 24670 35756 24676
rect 35624 24618 35676 24624
rect 35452 24398 35664 24426
rect 35268 23662 35296 24398
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 35256 23656 35308 23662
rect 35256 23598 35308 23604
rect 35268 23526 35296 23598
rect 35256 23520 35308 23526
rect 35256 23462 35308 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35256 23248 35308 23254
rect 34808 23174 34928 23202
rect 35256 23190 35308 23196
rect 34900 22522 34928 23174
rect 35268 22642 35296 23190
rect 35360 23118 35388 24006
rect 35452 23322 35480 24142
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 35440 23180 35492 23186
rect 35440 23122 35492 23128
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35256 22636 35308 22642
rect 35256 22578 35308 22584
rect 34900 22494 35388 22522
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34716 22066 34836 22094
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34716 21690 34744 21966
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34716 21554 34744 21626
rect 34704 21548 34756 21554
rect 34704 21490 34756 21496
rect 34612 19338 34664 19344
rect 34520 19304 34572 19310
rect 34612 19280 34664 19286
rect 34520 19246 34572 19252
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34244 17332 34296 17338
rect 34244 17274 34296 17280
rect 34256 16561 34284 17274
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34348 16794 34376 17138
rect 34336 16788 34388 16794
rect 34336 16730 34388 16736
rect 34242 16552 34298 16561
rect 34242 16487 34298 16496
rect 34440 16046 34468 17614
rect 34532 17202 34560 19246
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34428 16040 34480 16046
rect 34428 15982 34480 15988
rect 34336 15904 34388 15910
rect 34336 15846 34388 15852
rect 34348 14822 34376 15846
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14414 34376 14758
rect 34336 14408 34388 14414
rect 34336 14350 34388 14356
rect 34426 14240 34482 14249
rect 34426 14175 34482 14184
rect 34440 14074 34468 14175
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34242 13832 34298 13841
rect 34242 13767 34298 13776
rect 34256 13394 34284 13767
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34440 13326 34468 14010
rect 34428 13320 34480 13326
rect 34428 13262 34480 13268
rect 34532 13258 34560 16390
rect 34624 16250 34652 18702
rect 34716 18426 34744 21490
rect 34808 20398 34836 22066
rect 35072 22024 35124 22030
rect 35072 21966 35124 21972
rect 35084 21622 35112 21966
rect 35360 21944 35388 22494
rect 35452 22098 35480 23122
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35360 21916 35480 21944
rect 35346 21856 35402 21865
rect 35346 21791 35402 21800
rect 35072 21616 35124 21622
rect 35072 21558 35124 21564
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34888 20936 34940 20942
rect 34888 20878 34940 20884
rect 34900 20466 34928 20878
rect 35360 20482 35388 21791
rect 35452 21690 35480 21916
rect 35544 21894 35572 23666
rect 35636 23610 35664 24398
rect 35820 24070 35848 25434
rect 35912 25294 35940 26182
rect 36096 26042 36124 26250
rect 36084 26036 36136 26042
rect 36084 25978 36136 25984
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35900 24812 35952 24818
rect 35900 24754 35952 24760
rect 35912 24206 35940 24754
rect 35900 24200 35952 24206
rect 35900 24142 35952 24148
rect 35808 24064 35860 24070
rect 35808 24006 35860 24012
rect 35820 23730 35848 24006
rect 35808 23724 35860 23730
rect 35808 23666 35860 23672
rect 35636 23582 35848 23610
rect 35716 23248 35768 23254
rect 35716 23190 35768 23196
rect 35728 23050 35756 23190
rect 35624 23044 35676 23050
rect 35624 22986 35676 22992
rect 35716 23044 35768 23050
rect 35716 22986 35768 22992
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 35636 21706 35664 22986
rect 35716 22432 35768 22438
rect 35716 22374 35768 22380
rect 35728 22098 35756 22374
rect 35716 22092 35768 22098
rect 35716 22034 35768 22040
rect 35820 21978 35848 23582
rect 36004 23526 36032 24890
rect 36556 24818 36584 28358
rect 36924 27130 36952 34886
rect 36912 27124 36964 27130
rect 36912 27066 36964 27072
rect 36820 26784 36872 26790
rect 36818 26752 36820 26761
rect 36872 26752 36874 26761
rect 36818 26687 36874 26696
rect 36544 24812 36596 24818
rect 36820 24812 36872 24818
rect 36596 24772 36676 24800
rect 36544 24754 36596 24760
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 36556 23526 36584 24142
rect 35992 23520 36044 23526
rect 35992 23462 36044 23468
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36360 23044 36412 23050
rect 36360 22986 36412 22992
rect 36084 22976 36136 22982
rect 36004 22936 36084 22964
rect 36004 22658 36032 22936
rect 36084 22918 36136 22924
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 35912 22642 36032 22658
rect 35900 22636 36032 22642
rect 35952 22630 36032 22636
rect 35900 22578 35952 22584
rect 35992 22568 36044 22574
rect 35992 22510 36044 22516
rect 36004 22234 36032 22510
rect 36176 22500 36228 22506
rect 36176 22442 36228 22448
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 36188 22166 36216 22442
rect 36176 22160 36228 22166
rect 36176 22102 36228 22108
rect 35728 21950 35848 21978
rect 35728 21865 35756 21950
rect 35808 21888 35860 21894
rect 35714 21856 35770 21865
rect 35808 21830 35860 21836
rect 35714 21791 35770 21800
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 35544 21678 35756 21706
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35452 20777 35480 21490
rect 35544 20942 35572 21678
rect 35728 21554 35756 21678
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35636 21146 35664 21490
rect 35716 21344 35768 21350
rect 35714 21312 35716 21321
rect 35768 21312 35770 21321
rect 35714 21247 35770 21256
rect 35624 21140 35676 21146
rect 35624 21082 35676 21088
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 35532 20800 35584 20806
rect 35438 20768 35494 20777
rect 35532 20742 35584 20748
rect 35438 20703 35494 20712
rect 35544 20602 35572 20742
rect 35636 20641 35664 21082
rect 35820 21026 35848 21830
rect 36188 21690 36216 22102
rect 36280 21962 36308 22714
rect 36268 21956 36320 21962
rect 36268 21898 36320 21904
rect 36176 21684 36228 21690
rect 36176 21626 36228 21632
rect 36084 21616 36136 21622
rect 36136 21564 36308 21570
rect 36084 21558 36308 21564
rect 36096 21542 36308 21558
rect 35992 21412 36044 21418
rect 35992 21354 36044 21360
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35728 20998 35848 21026
rect 35622 20632 35678 20641
rect 35532 20596 35584 20602
rect 35622 20567 35678 20576
rect 35532 20538 35584 20544
rect 35728 20482 35756 20998
rect 35808 20868 35860 20874
rect 35808 20810 35860 20816
rect 34888 20460 34940 20466
rect 35360 20454 35572 20482
rect 34888 20402 34940 20408
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34704 18420 34756 18426
rect 34704 18362 34756 18368
rect 34716 17746 34744 18362
rect 34704 17740 34756 17746
rect 34704 17682 34756 17688
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34808 15994 34836 20334
rect 35440 20256 35492 20262
rect 35440 20198 35492 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35452 19854 35480 20198
rect 35544 19922 35572 20454
rect 35636 20454 35756 20482
rect 35636 20058 35664 20454
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35624 20052 35676 20058
rect 35624 19994 35676 20000
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 35360 19378 35388 19790
rect 35544 19718 35572 19858
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 35532 19712 35584 19718
rect 35532 19654 35584 19660
rect 35452 19378 35480 19654
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 35440 19372 35492 19378
rect 35492 19320 35572 19334
rect 35440 19314 35572 19320
rect 35360 19258 35388 19314
rect 35452 19306 35572 19314
rect 35360 19230 35480 19258
rect 35256 19168 35308 19174
rect 35308 19128 35388 19156
rect 35256 19110 35308 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18630 35388 19128
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35452 18290 35480 19230
rect 35544 18902 35572 19306
rect 35532 18896 35584 18902
rect 35532 18838 35584 18844
rect 35532 18760 35584 18766
rect 35530 18728 35532 18737
rect 35584 18728 35586 18737
rect 35530 18663 35586 18672
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 35624 18148 35676 18154
rect 35624 18090 35676 18096
rect 35440 18080 35492 18086
rect 35440 18022 35492 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35452 17746 35480 18022
rect 35440 17740 35492 17746
rect 35440 17682 35492 17688
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35256 16516 35308 16522
rect 35256 16458 35308 16464
rect 34716 15966 34836 15994
rect 34716 15434 34744 15966
rect 34796 15904 34848 15910
rect 34796 15846 34848 15852
rect 35268 15858 35296 16458
rect 35360 16250 35388 17206
rect 35532 16720 35584 16726
rect 35532 16662 35584 16668
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 35440 16108 35492 16114
rect 35440 16050 35492 16056
rect 34808 15706 34836 15846
rect 35268 15830 35388 15858
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15706 35388 15830
rect 34796 15700 34848 15706
rect 35348 15700 35400 15706
rect 34796 15642 34848 15648
rect 35268 15660 35348 15688
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 34716 15026 34744 15370
rect 35268 15162 35296 15660
rect 35348 15642 35400 15648
rect 35346 15192 35402 15201
rect 35256 15156 35308 15162
rect 35346 15127 35402 15136
rect 35256 15098 35308 15104
rect 35268 15026 35296 15098
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 35360 14958 35388 15127
rect 35452 15026 35480 16050
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35348 14952 35400 14958
rect 35348 14894 35400 14900
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34980 14544 35032 14550
rect 34980 14486 35032 14492
rect 34992 13938 35020 14486
rect 35360 14328 35388 14758
rect 35268 14300 35388 14328
rect 35268 13938 35296 14300
rect 34980 13932 35032 13938
rect 34980 13874 35032 13880
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 35348 13932 35400 13938
rect 35348 13874 35400 13880
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34428 12844 34480 12850
rect 34532 12832 34560 13194
rect 34808 12918 34836 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 12986 35388 13874
rect 35544 13530 35572 16662
rect 35636 16017 35664 18090
rect 35622 16008 35678 16017
rect 35622 15943 35678 15952
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 35636 15570 35664 15846
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 35636 15026 35664 15506
rect 35624 15020 35676 15026
rect 35624 14962 35676 14968
rect 35532 13524 35584 13530
rect 35532 13466 35584 13472
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 35544 12850 35572 13466
rect 35636 13462 35664 14962
rect 35728 14482 35756 20334
rect 35820 20058 35848 20810
rect 35912 20466 35940 21286
rect 36004 20942 36032 21354
rect 36176 21140 36228 21146
rect 36176 21082 36228 21088
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 36084 20868 36136 20874
rect 36084 20810 36136 20816
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 36004 20534 36032 20742
rect 36096 20534 36124 20810
rect 35992 20528 36044 20534
rect 35992 20470 36044 20476
rect 36084 20528 36136 20534
rect 36084 20470 36136 20476
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35900 19984 35952 19990
rect 35900 19926 35952 19932
rect 35992 19984 36044 19990
rect 35992 19926 36044 19932
rect 35808 19780 35860 19786
rect 35808 19722 35860 19728
rect 35820 19378 35848 19722
rect 35808 19372 35860 19378
rect 35808 19314 35860 19320
rect 35912 18873 35940 19926
rect 36004 19446 36032 19926
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36096 19446 36124 19790
rect 35992 19440 36044 19446
rect 35992 19382 36044 19388
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 35898 18864 35954 18873
rect 35898 18799 35954 18808
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 35820 16130 35848 18226
rect 35900 18080 35952 18086
rect 35900 18022 35952 18028
rect 35912 17542 35940 18022
rect 35900 17536 35952 17542
rect 35900 17478 35952 17484
rect 35820 16102 35940 16130
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35728 14006 35756 14418
rect 35716 14000 35768 14006
rect 35716 13942 35768 13948
rect 35624 13456 35676 13462
rect 35624 13398 35676 13404
rect 35532 12844 35584 12850
rect 34480 12804 34652 12832
rect 34428 12786 34480 12792
rect 34520 12708 34572 12714
rect 34520 12650 34572 12656
rect 34532 12434 34560 12650
rect 34348 12406 34560 12434
rect 34348 12238 34376 12406
rect 34624 12322 34652 12804
rect 35532 12786 35584 12792
rect 35820 12714 35848 15982
rect 35912 15434 35940 16102
rect 36004 15586 36032 19246
rect 36096 18970 36124 19382
rect 36084 18964 36136 18970
rect 36084 18906 36136 18912
rect 36188 18290 36216 21082
rect 36280 20346 36308 21542
rect 36372 21010 36400 22986
rect 36464 22642 36492 23462
rect 36452 22636 36504 22642
rect 36452 22578 36504 22584
rect 36452 22092 36504 22098
rect 36452 22034 36504 22040
rect 36464 21894 36492 22034
rect 36452 21888 36504 21894
rect 36452 21830 36504 21836
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 36372 20466 36400 20946
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36360 20460 36412 20466
rect 36360 20402 36412 20408
rect 36464 20346 36492 20878
rect 36280 20318 36492 20346
rect 36360 20256 36412 20262
rect 36360 20198 36412 20204
rect 36372 19854 36400 20198
rect 36464 19990 36492 20318
rect 36452 19984 36504 19990
rect 36452 19926 36504 19932
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 36372 19378 36400 19790
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36360 19372 36412 19378
rect 36280 19320 36360 19334
rect 36280 19314 36412 19320
rect 36280 19306 36400 19314
rect 36176 18284 36228 18290
rect 36176 18226 36228 18232
rect 36188 17882 36216 18226
rect 36176 17876 36228 17882
rect 36176 17818 36228 17824
rect 36280 17746 36308 19306
rect 36464 19174 36492 19654
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 36360 18896 36412 18902
rect 36360 18838 36412 18844
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 36096 16590 36124 17478
rect 36268 16992 36320 16998
rect 36268 16934 36320 16940
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 36176 15972 36228 15978
rect 36176 15914 36228 15920
rect 36004 15558 36124 15586
rect 35992 15496 36044 15502
rect 35992 15438 36044 15444
rect 35900 15428 35952 15434
rect 35900 15370 35952 15376
rect 35900 15020 35952 15026
rect 35900 14962 35952 14968
rect 35912 12918 35940 14962
rect 36004 14550 36032 15438
rect 36096 15026 36124 15558
rect 36188 15366 36216 15914
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 36084 15020 36136 15026
rect 36084 14962 36136 14968
rect 36084 14884 36136 14890
rect 36084 14826 36136 14832
rect 35992 14544 36044 14550
rect 35992 14486 36044 14492
rect 36096 14414 36124 14826
rect 36188 14521 36216 15098
rect 36280 15026 36308 16934
rect 36372 15502 36400 18838
rect 36464 18698 36492 19110
rect 36452 18692 36504 18698
rect 36452 18634 36504 18640
rect 36464 18086 36492 18634
rect 36556 18290 36584 23462
rect 36648 22642 36676 24772
rect 36820 24754 36872 24760
rect 36832 24682 36860 24754
rect 36820 24676 36872 24682
rect 36820 24618 36872 24624
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 36740 23118 36768 23666
rect 36832 23526 36860 24142
rect 37004 23656 37056 23662
rect 37002 23624 37004 23633
rect 37056 23624 37058 23633
rect 37002 23559 37058 23568
rect 36820 23520 36872 23526
rect 36820 23462 36872 23468
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36636 22636 36688 22642
rect 36636 22578 36688 22584
rect 36832 22094 36860 23462
rect 36912 23044 36964 23050
rect 36912 22986 36964 22992
rect 36740 22066 36860 22094
rect 36740 21962 36768 22066
rect 36820 22024 36872 22030
rect 36820 21966 36872 21972
rect 36728 21956 36780 21962
rect 36728 21898 36780 21904
rect 36636 21616 36688 21622
rect 36636 21558 36688 21564
rect 36648 20942 36676 21558
rect 36740 21146 36768 21898
rect 36832 21690 36860 21966
rect 36820 21684 36872 21690
rect 36820 21626 36872 21632
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36820 21140 36872 21146
rect 36820 21082 36872 21088
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36648 20466 36676 20878
rect 36832 20806 36860 21082
rect 36820 20800 36872 20806
rect 36820 20742 36872 20748
rect 36636 20460 36688 20466
rect 36636 20402 36688 20408
rect 36648 20262 36676 20402
rect 36636 20256 36688 20262
rect 36636 20198 36688 20204
rect 36634 19408 36690 19417
rect 36634 19343 36636 19352
rect 36688 19343 36690 19352
rect 36636 19314 36688 19320
rect 36636 19236 36688 19242
rect 36636 19178 36688 19184
rect 36648 18902 36676 19178
rect 36636 18896 36688 18902
rect 36636 18838 36688 18844
rect 36648 18698 36676 18838
rect 36636 18692 36688 18698
rect 36636 18634 36688 18640
rect 36924 18358 36952 22986
rect 37004 22092 37056 22098
rect 37004 22034 37056 22040
rect 37016 21622 37044 22034
rect 37004 21616 37056 21622
rect 37004 21558 37056 21564
rect 37004 19984 37056 19990
rect 37004 19926 37056 19932
rect 36912 18352 36964 18358
rect 36912 18294 36964 18300
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 36556 17338 36584 18226
rect 36820 17808 36872 17814
rect 37016 17762 37044 19926
rect 36820 17750 36872 17756
rect 36728 17672 36780 17678
rect 36726 17640 36728 17649
rect 36780 17640 36782 17649
rect 36726 17575 36782 17584
rect 36832 17338 36860 17750
rect 36924 17734 37044 17762
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36820 17332 36872 17338
rect 36820 17274 36872 17280
rect 36556 17218 36584 17274
rect 36556 17202 36676 17218
rect 36556 17196 36688 17202
rect 36556 17190 36636 17196
rect 36636 17138 36688 17144
rect 36636 17060 36688 17066
rect 36636 17002 36688 17008
rect 36544 16992 36596 16998
rect 36544 16934 36596 16940
rect 36452 16584 36504 16590
rect 36452 16526 36504 16532
rect 36464 16028 36492 16526
rect 36556 16182 36584 16934
rect 36648 16658 36676 17002
rect 36728 16992 36780 16998
rect 36728 16934 36780 16940
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36544 16176 36596 16182
rect 36648 16153 36676 16594
rect 36544 16118 36596 16124
rect 36634 16144 36690 16153
rect 36634 16079 36690 16088
rect 36544 16040 36596 16046
rect 36464 16000 36544 16028
rect 36544 15982 36596 15988
rect 36452 15632 36504 15638
rect 36452 15574 36504 15580
rect 36360 15496 36412 15502
rect 36360 15438 36412 15444
rect 36360 15360 36412 15366
rect 36360 15302 36412 15308
rect 36372 15162 36400 15302
rect 36464 15162 36492 15574
rect 36360 15156 36412 15162
rect 36360 15098 36412 15104
rect 36452 15156 36504 15162
rect 36452 15098 36504 15104
rect 36268 15020 36320 15026
rect 36320 14980 36400 15008
rect 36268 14962 36320 14968
rect 36174 14512 36230 14521
rect 36174 14447 36230 14456
rect 36268 14476 36320 14482
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 35900 12912 35952 12918
rect 35900 12854 35952 12860
rect 36188 12850 36216 14447
rect 36268 14418 36320 14424
rect 36280 13462 36308 14418
rect 36372 14346 36400 14980
rect 36360 14340 36412 14346
rect 36360 14282 36412 14288
rect 36464 14226 36492 15098
rect 36556 14618 36584 15982
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 36464 14198 36584 14226
rect 36556 14074 36584 14198
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 36360 13728 36412 13734
rect 36360 13670 36412 13676
rect 36268 13456 36320 13462
rect 36268 13398 36320 13404
rect 36176 12844 36228 12850
rect 36176 12786 36228 12792
rect 35808 12708 35860 12714
rect 35808 12650 35860 12656
rect 34704 12640 34756 12646
rect 34704 12582 34756 12588
rect 34440 12306 34652 12322
rect 34428 12300 34652 12306
rect 34480 12294 34652 12300
rect 34428 12242 34480 12248
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34244 12096 34296 12102
rect 34244 12038 34296 12044
rect 34428 12096 34480 12102
rect 34428 12038 34480 12044
rect 34256 11898 34284 12038
rect 34244 11892 34296 11898
rect 34244 11834 34296 11840
rect 34440 11830 34468 12038
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34440 10742 34468 11086
rect 34428 10736 34480 10742
rect 34428 10678 34480 10684
rect 34624 10674 34652 12174
rect 34716 11830 34744 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36372 12434 36400 13670
rect 36464 13530 36492 14010
rect 36648 13938 36676 16079
rect 36740 15910 36768 16934
rect 36728 15904 36780 15910
rect 36728 15846 36780 15852
rect 36636 13932 36688 13938
rect 36636 13874 36688 13880
rect 36452 13524 36504 13530
rect 36452 13466 36504 13472
rect 36636 13456 36688 13462
rect 36636 13398 36688 13404
rect 36726 13424 36782 13433
rect 36648 12986 36676 13398
rect 36726 13359 36728 13368
rect 36780 13359 36782 13368
rect 36728 13330 36780 13336
rect 36636 12980 36688 12986
rect 36636 12922 36688 12928
rect 36728 12844 36780 12850
rect 36728 12786 36780 12792
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 36372 12406 36492 12434
rect 35348 12368 35400 12374
rect 35532 12368 35584 12374
rect 35400 12316 35532 12322
rect 35348 12310 35584 12316
rect 34796 12300 34848 12306
rect 35360 12294 35572 12310
rect 34796 12242 34848 12248
rect 34704 11824 34756 11830
rect 34704 11766 34756 11772
rect 34808 11642 34836 12242
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 35820 11830 35848 12038
rect 35532 11824 35584 11830
rect 35532 11766 35584 11772
rect 35808 11824 35860 11830
rect 35808 11766 35860 11772
rect 34716 11614 34836 11642
rect 34716 10742 34744 11614
rect 34796 11552 34848 11558
rect 34796 11494 34848 11500
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 34716 10606 34744 10678
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34532 9586 34560 10134
rect 34808 9586 34836 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35544 11354 35572 11766
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 35900 11552 35952 11558
rect 35900 11494 35952 11500
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35728 10742 35756 11086
rect 35716 10736 35768 10742
rect 35716 10678 35768 10684
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35716 9920 35768 9926
rect 35716 9862 35768 9868
rect 35728 9586 35756 9862
rect 34520 9580 34572 9586
rect 34520 9522 34572 9528
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35716 9580 35768 9586
rect 35716 9522 35768 9528
rect 34532 8974 34560 9522
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34808 8498 34836 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35544 8974 35572 9522
rect 35624 9376 35676 9382
rect 35624 9318 35676 9324
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35636 8634 35664 9318
rect 35728 9042 35756 9522
rect 35716 9036 35768 9042
rect 35716 8978 35768 8984
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35912 8498 35940 11494
rect 36280 10742 36308 11698
rect 36360 11552 36412 11558
rect 36360 11494 36412 11500
rect 36372 11286 36400 11494
rect 36360 11280 36412 11286
rect 36360 11222 36412 11228
rect 36464 11150 36492 12406
rect 36648 12306 36676 12582
rect 36740 12442 36768 12786
rect 36832 12782 36860 17274
rect 36924 17066 36952 17734
rect 37002 17640 37058 17649
rect 37002 17575 37058 17584
rect 36912 17060 36964 17066
rect 36912 17002 36964 17008
rect 37016 16114 37044 17575
rect 37004 16108 37056 16114
rect 37004 16050 37056 16056
rect 36912 15904 36964 15910
rect 36912 15846 36964 15852
rect 36924 15638 36952 15846
rect 36912 15632 36964 15638
rect 36912 15574 36964 15580
rect 36912 15496 36964 15502
rect 36912 15438 36964 15444
rect 36924 15094 36952 15438
rect 36912 15088 36964 15094
rect 36912 15030 36964 15036
rect 36924 14414 36952 15030
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 36924 12850 36952 14350
rect 36912 12844 36964 12850
rect 36912 12786 36964 12792
rect 36820 12776 36872 12782
rect 36820 12718 36872 12724
rect 36728 12436 36780 12442
rect 36728 12378 36780 12384
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 36556 11626 36584 12038
rect 36728 11756 36780 11762
rect 36728 11698 36780 11704
rect 36912 11756 36964 11762
rect 36912 11698 36964 11704
rect 36544 11620 36596 11626
rect 36544 11562 36596 11568
rect 36740 11354 36768 11698
rect 36728 11348 36780 11354
rect 36728 11290 36780 11296
rect 36924 11150 36952 11698
rect 37004 11348 37056 11354
rect 37004 11290 37056 11296
rect 37016 11218 37044 11290
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36912 11144 36964 11150
rect 36912 11086 36964 11092
rect 36464 10742 36492 11086
rect 36268 10736 36320 10742
rect 36268 10678 36320 10684
rect 36452 10736 36504 10742
rect 36452 10678 36504 10684
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 36096 10130 36124 10406
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 36924 9722 36952 11086
rect 36912 9716 36964 9722
rect 36912 9658 36964 9664
rect 36084 8832 36136 8838
rect 36084 8774 36136 8780
rect 36096 8498 36124 8774
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34164 2746 34468 2774
rect 34440 2582 34468 2746
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 37108 2650 37136 38218
rect 37464 34604 37516 34610
rect 37464 34546 37516 34552
rect 37476 33658 37504 34546
rect 38936 34468 38988 34474
rect 38936 34410 38988 34416
rect 38948 33998 38976 34410
rect 40224 34128 40276 34134
rect 40224 34070 40276 34076
rect 38936 33992 38988 33998
rect 38936 33934 38988 33940
rect 38844 33924 38896 33930
rect 38844 33866 38896 33872
rect 38752 33856 38804 33862
rect 38752 33798 38804 33804
rect 38764 33658 38792 33798
rect 37464 33652 37516 33658
rect 38752 33652 38804 33658
rect 37464 33594 37516 33600
rect 38672 33612 38752 33640
rect 37476 33522 37504 33594
rect 37464 33516 37516 33522
rect 37464 33458 37516 33464
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 37292 31822 37320 32914
rect 37556 32904 37608 32910
rect 37556 32846 37608 32852
rect 37464 32224 37516 32230
rect 37464 32166 37516 32172
rect 37476 32065 37504 32166
rect 37462 32056 37518 32065
rect 37462 31991 37518 32000
rect 37568 31958 37596 32846
rect 38672 32842 38700 33612
rect 38752 33594 38804 33600
rect 38856 33590 38884 33866
rect 38844 33584 38896 33590
rect 38844 33526 38896 33532
rect 38752 33312 38804 33318
rect 38752 33254 38804 33260
rect 38660 32836 38712 32842
rect 38660 32778 38712 32784
rect 37924 32768 37976 32774
rect 37924 32710 37976 32716
rect 37936 32434 37964 32710
rect 38764 32502 38792 33254
rect 38856 33114 38884 33526
rect 38948 33522 38976 33934
rect 38936 33516 38988 33522
rect 38936 33458 38988 33464
rect 39672 33516 39724 33522
rect 39672 33458 39724 33464
rect 40040 33516 40092 33522
rect 40040 33458 40092 33464
rect 38844 33108 38896 33114
rect 38844 33050 38896 33056
rect 38948 32842 38976 33458
rect 38936 32836 38988 32842
rect 38936 32778 38988 32784
rect 39028 32768 39080 32774
rect 39028 32710 39080 32716
rect 38752 32496 38804 32502
rect 38752 32438 38804 32444
rect 39040 32434 39068 32710
rect 39684 32570 39712 33458
rect 40052 33114 40080 33458
rect 40040 33108 40092 33114
rect 40040 33050 40092 33056
rect 40236 32910 40264 34070
rect 40224 32904 40276 32910
rect 40224 32846 40276 32852
rect 39672 32564 39724 32570
rect 39672 32506 39724 32512
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 37924 32428 37976 32434
rect 37924 32370 37976 32376
rect 39028 32428 39080 32434
rect 39028 32370 39080 32376
rect 37660 32026 37688 32370
rect 37648 32020 37700 32026
rect 37648 31962 37700 31968
rect 37556 31952 37608 31958
rect 37556 31894 37608 31900
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 37188 31136 37240 31142
rect 37188 31078 37240 31084
rect 37200 30734 37228 31078
rect 41340 30802 41368 57394
rect 37280 30796 37332 30802
rect 37280 30738 37332 30744
rect 41328 30796 41380 30802
rect 41328 30738 41380 30744
rect 37188 30728 37240 30734
rect 37188 30670 37240 30676
rect 37292 30326 37320 30738
rect 37280 30320 37332 30326
rect 37280 30262 37332 30268
rect 37188 29232 37240 29238
rect 37188 29174 37240 29180
rect 37200 28490 37228 29174
rect 37188 28484 37240 28490
rect 37188 28426 37240 28432
rect 39488 28484 39540 28490
rect 39488 28426 39540 28432
rect 37200 27402 37228 28426
rect 38382 27432 38438 27441
rect 37188 27396 37240 27402
rect 37924 27396 37976 27402
rect 37240 27356 37320 27384
rect 37188 27338 37240 27344
rect 37188 27124 37240 27130
rect 37188 27066 37240 27072
rect 37200 26586 37228 27066
rect 37188 26580 37240 26586
rect 37188 26522 37240 26528
rect 37292 26450 37320 27356
rect 38382 27367 38384 27376
rect 37924 27338 37976 27344
rect 38436 27367 38438 27376
rect 38384 27338 38436 27344
rect 37280 26444 37332 26450
rect 37280 26386 37332 26392
rect 37292 25294 37320 26386
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 37648 25152 37700 25158
rect 37648 25094 37700 25100
rect 37660 24886 37688 25094
rect 37648 24880 37700 24886
rect 37648 24822 37700 24828
rect 37936 24818 37964 27338
rect 38396 26994 38424 27338
rect 39500 27130 39528 28426
rect 39488 27124 39540 27130
rect 39488 27066 39540 27072
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38396 26450 38424 26930
rect 38844 26920 38896 26926
rect 38844 26862 38896 26868
rect 38752 26784 38804 26790
rect 38752 26726 38804 26732
rect 38384 26444 38436 26450
rect 38384 26386 38436 26392
rect 38016 26308 38068 26314
rect 38016 26250 38068 26256
rect 38028 25838 38056 26250
rect 38016 25832 38068 25838
rect 38016 25774 38068 25780
rect 38028 25430 38056 25774
rect 38396 25770 38424 26386
rect 38764 26314 38792 26726
rect 38752 26308 38804 26314
rect 38752 26250 38804 26256
rect 38384 25764 38436 25770
rect 38384 25706 38436 25712
rect 38016 25424 38068 25430
rect 38016 25366 38068 25372
rect 38028 24818 38056 25366
rect 38108 25152 38160 25158
rect 38108 25094 38160 25100
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37292 24206 37320 24550
rect 37830 24440 37886 24449
rect 37936 24410 37964 24754
rect 37830 24375 37832 24384
rect 37884 24375 37886 24384
rect 37924 24404 37976 24410
rect 37832 24346 37884 24352
rect 37924 24346 37976 24352
rect 37280 24200 37332 24206
rect 37280 24142 37332 24148
rect 37188 24132 37240 24138
rect 37188 24074 37240 24080
rect 37200 23254 37228 24074
rect 37188 23248 37240 23254
rect 37188 23190 37240 23196
rect 37292 23118 37320 24142
rect 38028 23730 38056 24754
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37200 22710 37228 22918
rect 37188 22704 37240 22710
rect 37188 22646 37240 22652
rect 37200 21554 37228 22646
rect 37384 21894 37412 23666
rect 37924 23656 37976 23662
rect 37476 23604 37924 23610
rect 37476 23598 37976 23604
rect 37476 23582 37964 23598
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37188 21412 37240 21418
rect 37188 21354 37240 21360
rect 37200 21010 37228 21354
rect 37188 21004 37240 21010
rect 37188 20946 37240 20952
rect 37292 20942 37320 21422
rect 37280 20936 37332 20942
rect 37476 20913 37504 23582
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 37556 22568 37608 22574
rect 37556 22510 37608 22516
rect 37568 21690 37596 22510
rect 38028 22234 38056 22578
rect 37740 22228 37792 22234
rect 37740 22170 37792 22176
rect 38016 22228 38068 22234
rect 38016 22170 38068 22176
rect 37752 21962 37780 22170
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 37740 21956 37792 21962
rect 37740 21898 37792 21904
rect 37752 21865 37780 21898
rect 37738 21856 37794 21865
rect 37738 21791 37794 21800
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 37648 21548 37700 21554
rect 37700 21508 37780 21536
rect 37648 21490 37700 21496
rect 37752 21146 37780 21508
rect 37648 21140 37700 21146
rect 37648 21082 37700 21088
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 37660 21010 37688 21082
rect 37648 21004 37700 21010
rect 37648 20946 37700 20952
rect 37740 20936 37792 20942
rect 37280 20878 37332 20884
rect 37462 20904 37518 20913
rect 37740 20878 37792 20884
rect 37462 20839 37464 20848
rect 37516 20839 37518 20848
rect 37464 20810 37516 20816
rect 37280 20800 37332 20806
rect 37280 20742 37332 20748
rect 37556 20800 37608 20806
rect 37556 20742 37608 20748
rect 37188 17604 37240 17610
rect 37188 17546 37240 17552
rect 37200 17066 37228 17546
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 37292 16794 37320 20742
rect 37462 20632 37518 20641
rect 37568 20602 37596 20742
rect 37462 20567 37518 20576
rect 37556 20596 37608 20602
rect 37476 20466 37504 20567
rect 37556 20538 37608 20544
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37752 20330 37780 20878
rect 37740 20324 37792 20330
rect 37740 20266 37792 20272
rect 37844 20233 37872 21626
rect 38028 21593 38056 21966
rect 38014 21584 38070 21593
rect 38014 21519 38070 21528
rect 37924 21480 37976 21486
rect 37924 21422 37976 21428
rect 37830 20224 37886 20233
rect 37830 20159 37886 20168
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37476 19718 37504 19790
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37464 19712 37516 19718
rect 37844 19689 37872 19790
rect 37464 19654 37516 19660
rect 37830 19680 37886 19689
rect 37384 19446 37412 19654
rect 37372 19440 37424 19446
rect 37372 19382 37424 19388
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37384 18763 37412 19246
rect 37476 18902 37504 19654
rect 37830 19615 37886 19624
rect 37740 19508 37792 19514
rect 37740 19450 37792 19456
rect 37752 19378 37780 19450
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 37556 19168 37608 19174
rect 37556 19110 37608 19116
rect 37464 18896 37516 18902
rect 37464 18838 37516 18844
rect 37381 18757 37433 18763
rect 37381 18699 37433 18705
rect 37384 18646 37421 18699
rect 37384 18290 37412 18646
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37384 16794 37412 17818
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 37372 16788 37424 16794
rect 37372 16730 37424 16736
rect 37292 16590 37320 16730
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37372 15904 37424 15910
rect 37372 15846 37424 15852
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 37292 13938 37320 15438
rect 37384 14890 37412 15846
rect 37372 14884 37424 14890
rect 37372 14826 37424 14832
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 37476 13394 37504 18838
rect 37568 17746 37596 19110
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 37740 18760 37792 18766
rect 37740 18702 37792 18708
rect 37556 17740 37608 17746
rect 37556 17682 37608 17688
rect 37554 17640 37610 17649
rect 37660 17610 37688 18702
rect 37752 18222 37780 18702
rect 37844 18426 37872 19615
rect 37936 19378 37964 21422
rect 37924 19372 37976 19378
rect 37924 19314 37976 19320
rect 37936 19174 37964 19314
rect 37924 19168 37976 19174
rect 37924 19110 37976 19116
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37936 18737 37964 18770
rect 37922 18728 37978 18737
rect 37922 18663 37978 18672
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37554 17575 37610 17584
rect 37648 17604 37700 17610
rect 37568 17338 37596 17575
rect 37648 17546 37700 17552
rect 37556 17332 37608 17338
rect 37556 17274 37608 17280
rect 37752 17202 37780 17682
rect 37844 17377 37872 18226
rect 38028 18193 38056 21519
rect 38120 21321 38148 25094
rect 38764 24886 38792 26250
rect 38856 25226 38884 26862
rect 39500 26858 39528 27066
rect 43996 26920 44048 26926
rect 43996 26862 44048 26868
rect 39488 26852 39540 26858
rect 39488 26794 39540 26800
rect 39212 26376 39264 26382
rect 39212 26318 39264 26324
rect 39224 26042 39252 26318
rect 39212 26036 39264 26042
rect 39212 25978 39264 25984
rect 39500 25906 39528 26794
rect 41880 26784 41932 26790
rect 41880 26726 41932 26732
rect 40224 26512 40276 26518
rect 40224 26454 40276 26460
rect 40040 26376 40092 26382
rect 40040 26318 40092 26324
rect 39488 25900 39540 25906
rect 39488 25842 39540 25848
rect 39212 25492 39264 25498
rect 39212 25434 39264 25440
rect 38844 25220 38896 25226
rect 38844 25162 38896 25168
rect 38752 24880 38804 24886
rect 38752 24822 38804 24828
rect 38856 24818 38884 25162
rect 39224 25158 39252 25434
rect 39304 25356 39356 25362
rect 39304 25298 39356 25304
rect 39212 25152 39264 25158
rect 39212 25094 39264 25100
rect 38568 24812 38620 24818
rect 38568 24754 38620 24760
rect 38844 24812 38896 24818
rect 38844 24754 38896 24760
rect 38580 24682 38608 24754
rect 38752 24744 38804 24750
rect 38752 24686 38804 24692
rect 38568 24676 38620 24682
rect 38568 24618 38620 24624
rect 38580 23662 38608 24618
rect 38764 24342 38792 24686
rect 39212 24608 39264 24614
rect 39316 24596 39344 25298
rect 39264 24568 39344 24596
rect 39212 24550 39264 24556
rect 38752 24336 38804 24342
rect 38752 24278 38804 24284
rect 38568 23656 38620 23662
rect 38568 23598 38620 23604
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38476 23180 38528 23186
rect 38476 23122 38528 23128
rect 38292 22432 38344 22438
rect 38292 22374 38344 22380
rect 38200 22024 38252 22030
rect 38200 21966 38252 21972
rect 38212 21690 38240 21966
rect 38200 21684 38252 21690
rect 38200 21626 38252 21632
rect 38200 21548 38252 21554
rect 38200 21490 38252 21496
rect 38106 21312 38162 21321
rect 38106 21247 38162 21256
rect 38120 19514 38148 21247
rect 38212 19854 38240 21490
rect 38200 19848 38252 19854
rect 38200 19790 38252 19796
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 38200 19304 38252 19310
rect 38200 19246 38252 19252
rect 38212 18902 38240 19246
rect 38200 18896 38252 18902
rect 38200 18838 38252 18844
rect 38200 18624 38252 18630
rect 38200 18566 38252 18572
rect 38014 18184 38070 18193
rect 38014 18119 38070 18128
rect 37830 17368 37886 17377
rect 37830 17303 37886 17312
rect 37924 17332 37976 17338
rect 37556 17196 37608 17202
rect 37740 17196 37792 17202
rect 37556 17138 37608 17144
rect 37660 17156 37740 17184
rect 37568 16946 37596 17138
rect 37660 17066 37688 17156
rect 37740 17138 37792 17144
rect 37648 17060 37700 17066
rect 37648 17002 37700 17008
rect 37740 16992 37792 16998
rect 37568 16940 37740 16946
rect 37568 16934 37792 16940
rect 37568 16918 37780 16934
rect 37568 16114 37596 16918
rect 37844 16810 37872 17303
rect 37924 17274 37976 17280
rect 37936 17066 37964 17274
rect 37924 17060 37976 17066
rect 37924 17002 37976 17008
rect 37752 16782 37872 16810
rect 37648 16652 37700 16658
rect 37648 16594 37700 16600
rect 37660 16454 37688 16594
rect 37648 16448 37700 16454
rect 37648 16390 37700 16396
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37568 14414 37596 16050
rect 37752 15026 37780 16782
rect 37832 16516 37884 16522
rect 37832 16458 37884 16464
rect 37844 16250 37872 16458
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37936 16114 37964 17002
rect 38028 16998 38056 18119
rect 38212 18086 38240 18566
rect 38200 18080 38252 18086
rect 38200 18022 38252 18028
rect 38212 17882 38240 18022
rect 38200 17876 38252 17882
rect 38200 17818 38252 17824
rect 38106 17776 38162 17785
rect 38106 17711 38108 17720
rect 38160 17711 38162 17720
rect 38108 17682 38160 17688
rect 38106 17368 38162 17377
rect 38106 17303 38108 17312
rect 38160 17303 38162 17312
rect 38108 17274 38160 17280
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 38108 16992 38160 16998
rect 38212 16980 38240 17818
rect 38160 16952 38240 16980
rect 38108 16934 38160 16940
rect 38016 16788 38068 16794
rect 38016 16730 38068 16736
rect 37924 16108 37976 16114
rect 37924 16050 37976 16056
rect 37924 15904 37976 15910
rect 37924 15846 37976 15852
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37648 14272 37700 14278
rect 37648 14214 37700 14220
rect 37660 13870 37688 14214
rect 37844 14006 37872 14350
rect 37832 14000 37884 14006
rect 37936 13977 37964 15846
rect 38028 14346 38056 16730
rect 38120 15910 38148 16934
rect 38200 16720 38252 16726
rect 38200 16662 38252 16668
rect 38108 15904 38160 15910
rect 38108 15846 38160 15852
rect 38108 15428 38160 15434
rect 38108 15370 38160 15376
rect 38016 14340 38068 14346
rect 38016 14282 38068 14288
rect 37832 13942 37884 13948
rect 37922 13968 37978 13977
rect 37922 13903 37924 13912
rect 37976 13903 37978 13912
rect 38028 13920 38056 14282
rect 38120 14056 38148 15370
rect 38212 14346 38240 16662
rect 38304 15502 38332 22374
rect 38488 22250 38516 23122
rect 38672 22982 38700 23258
rect 38660 22976 38712 22982
rect 38660 22918 38712 22924
rect 38672 22642 38700 22918
rect 38660 22636 38712 22642
rect 38660 22578 38712 22584
rect 38488 22234 38654 22250
rect 38488 22228 38666 22234
rect 38488 22222 38614 22228
rect 38614 22170 38666 22176
rect 38384 22160 38436 22166
rect 38384 22102 38436 22108
rect 38396 21146 38424 22102
rect 38660 22092 38712 22098
rect 38488 22052 38660 22080
rect 38488 21729 38516 22052
rect 38660 22034 38712 22040
rect 38474 21720 38530 21729
rect 38474 21655 38530 21664
rect 38568 21548 38620 21554
rect 38568 21490 38620 21496
rect 38476 21480 38528 21486
rect 38476 21422 38528 21428
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38488 20602 38516 21422
rect 38580 20874 38608 21490
rect 38568 20868 38620 20874
rect 38568 20810 38620 20816
rect 38476 20596 38528 20602
rect 38476 20538 38528 20544
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38384 19168 38436 19174
rect 38384 19110 38436 19116
rect 38396 18698 38424 19110
rect 38384 18692 38436 18698
rect 38384 18634 38436 18640
rect 38396 18426 38424 18634
rect 38384 18420 38436 18426
rect 38384 18362 38436 18368
rect 38382 18320 38438 18329
rect 38382 18255 38384 18264
rect 38436 18255 38438 18264
rect 38384 18226 38436 18232
rect 38488 18086 38516 19790
rect 38660 19508 38712 19514
rect 38660 19450 38712 19456
rect 38566 18864 38622 18873
rect 38566 18799 38622 18808
rect 38580 18630 38608 18799
rect 38568 18624 38620 18630
rect 38568 18566 38620 18572
rect 38672 18290 38700 19450
rect 38660 18284 38712 18290
rect 38580 18244 38660 18272
rect 38476 18080 38528 18086
rect 38476 18022 38528 18028
rect 38384 17876 38436 17882
rect 38384 17818 38436 17824
rect 38396 17134 38424 17818
rect 38476 17604 38528 17610
rect 38476 17546 38528 17552
rect 38384 17128 38436 17134
rect 38384 17070 38436 17076
rect 38396 16726 38424 17070
rect 38384 16720 38436 16726
rect 38384 16662 38436 16668
rect 38292 15496 38344 15502
rect 38292 15438 38344 15444
rect 38488 15026 38516 17546
rect 38580 17066 38608 18244
rect 38660 18226 38712 18232
rect 38660 18148 38712 18154
rect 38660 18090 38712 18096
rect 38672 18057 38700 18090
rect 38658 18048 38714 18057
rect 38658 17983 38714 17992
rect 38660 17196 38712 17202
rect 38660 17138 38712 17144
rect 38568 17060 38620 17066
rect 38568 17002 38620 17008
rect 38568 15088 38620 15094
rect 38672 15076 38700 17138
rect 38620 15048 38700 15076
rect 38568 15030 38620 15036
rect 38476 15020 38528 15026
rect 38476 14962 38528 14968
rect 38566 14920 38622 14929
rect 38566 14855 38568 14864
rect 38620 14855 38622 14864
rect 38568 14826 38620 14832
rect 38292 14544 38344 14550
rect 38292 14486 38344 14492
rect 38476 14544 38528 14550
rect 38476 14486 38528 14492
rect 38566 14512 38622 14521
rect 38200 14340 38252 14346
rect 38200 14282 38252 14288
rect 38304 14278 38332 14486
rect 38384 14476 38436 14482
rect 38384 14418 38436 14424
rect 38292 14272 38344 14278
rect 38292 14214 38344 14220
rect 38120 14028 38240 14056
rect 38108 13932 38160 13938
rect 37924 13874 37976 13880
rect 38028 13892 38108 13920
rect 37648 13864 37700 13870
rect 37648 13806 37700 13812
rect 37740 13728 37792 13734
rect 37740 13670 37792 13676
rect 37752 13462 37780 13670
rect 37740 13456 37792 13462
rect 37740 13398 37792 13404
rect 37464 13388 37516 13394
rect 38028 13376 38056 13892
rect 38108 13874 38160 13880
rect 37464 13330 37516 13336
rect 37844 13348 38056 13376
rect 37740 13320 37792 13326
rect 37844 13308 37872 13348
rect 37792 13280 37872 13308
rect 37740 13262 37792 13268
rect 37752 13190 37780 13262
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37832 13184 37884 13190
rect 37832 13126 37884 13132
rect 37844 12850 37872 13126
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 37200 11234 37228 12038
rect 38212 11762 38240 14028
rect 38396 14006 38424 14418
rect 38384 14000 38436 14006
rect 38290 13968 38346 13977
rect 38384 13942 38436 13948
rect 38290 13903 38346 13912
rect 38304 12986 38332 13903
rect 38488 13841 38516 14486
rect 38566 14447 38622 14456
rect 38580 14346 38608 14447
rect 38658 14376 38714 14385
rect 38568 14340 38620 14346
rect 38658 14311 38714 14320
rect 38568 14282 38620 14288
rect 38672 14278 38700 14311
rect 38660 14272 38712 14278
rect 38660 14214 38712 14220
rect 38474 13832 38530 13841
rect 38474 13767 38530 13776
rect 38764 13394 38792 24278
rect 38844 24132 38896 24138
rect 38844 24074 38896 24080
rect 38856 23322 38884 24074
rect 39224 23526 39252 24550
rect 39304 24200 39356 24206
rect 39304 24142 39356 24148
rect 39316 23866 39344 24142
rect 39304 23860 39356 23866
rect 39304 23802 39356 23808
rect 39212 23520 39264 23526
rect 39212 23462 39264 23468
rect 38844 23316 38896 23322
rect 38844 23258 38896 23264
rect 38856 21554 38884 23258
rect 39120 23248 39172 23254
rect 39120 23190 39172 23196
rect 39132 22817 39160 23190
rect 39316 23118 39344 23802
rect 39394 23760 39450 23769
rect 39500 23730 39528 25842
rect 39948 25696 40000 25702
rect 39948 25638 40000 25644
rect 39672 24812 39724 24818
rect 39724 24772 39804 24800
rect 39672 24754 39724 24760
rect 39776 23730 39804 24772
rect 39394 23695 39450 23704
rect 39488 23724 39540 23730
rect 39304 23112 39356 23118
rect 39304 23054 39356 23060
rect 39118 22808 39174 22817
rect 39118 22743 39174 22752
rect 39132 22574 39160 22743
rect 39304 22704 39356 22710
rect 39302 22672 39304 22681
rect 39356 22672 39358 22681
rect 39302 22607 39358 22616
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 39120 22568 39172 22574
rect 39120 22510 39172 22516
rect 39040 21894 39068 22510
rect 39120 22432 39172 22438
rect 39120 22374 39172 22380
rect 39028 21888 39080 21894
rect 39028 21830 39080 21836
rect 38844 21548 38896 21554
rect 38844 21490 38896 21496
rect 38856 20942 38884 21490
rect 39132 20942 39160 22374
rect 39304 22094 39356 22098
rect 39408 22094 39436 23695
rect 39488 23666 39540 23672
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39764 23724 39816 23730
rect 39764 23666 39816 23672
rect 39488 23316 39540 23322
rect 39488 23258 39540 23264
rect 39500 23118 39528 23258
rect 39488 23112 39540 23118
rect 39488 23054 39540 23060
rect 39488 22772 39540 22778
rect 39488 22714 39540 22720
rect 39500 22506 39528 22714
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39488 22500 39540 22506
rect 39488 22442 39540 22448
rect 39500 22234 39528 22442
rect 39488 22228 39540 22234
rect 39488 22170 39540 22176
rect 39304 22092 39436 22094
rect 39356 22066 39436 22092
rect 39304 22034 39356 22040
rect 39304 21684 39356 21690
rect 39304 21626 39356 21632
rect 39212 21548 39264 21554
rect 39212 21490 39264 21496
rect 39224 21078 39252 21490
rect 39212 21072 39264 21078
rect 39212 21014 39264 21020
rect 38844 20936 38896 20942
rect 38844 20878 38896 20884
rect 39120 20936 39172 20942
rect 39120 20878 39172 20884
rect 39212 20868 39264 20874
rect 39212 20810 39264 20816
rect 39120 20800 39172 20806
rect 39120 20742 39172 20748
rect 39028 20596 39080 20602
rect 39028 20538 39080 20544
rect 39040 19786 39068 20538
rect 39028 19780 39080 19786
rect 39028 19722 39080 19728
rect 39132 19666 39160 20742
rect 39040 19638 39160 19666
rect 38936 19372 38988 19378
rect 38936 19314 38988 19320
rect 38844 19168 38896 19174
rect 38844 19110 38896 19116
rect 38856 18834 38884 19110
rect 38948 18902 38976 19314
rect 39040 18970 39068 19638
rect 39028 18964 39080 18970
rect 39028 18906 39080 18912
rect 38936 18896 38988 18902
rect 38936 18838 38988 18844
rect 38844 18828 38896 18834
rect 38844 18770 38896 18776
rect 38948 18714 38976 18838
rect 38856 18686 38976 18714
rect 38856 18222 38884 18686
rect 39040 18630 39068 18906
rect 39224 18698 39252 20810
rect 39316 20602 39344 21626
rect 39488 21480 39540 21486
rect 39488 21422 39540 21428
rect 39396 21344 39448 21350
rect 39396 21286 39448 21292
rect 39408 21010 39436 21286
rect 39396 21004 39448 21010
rect 39396 20946 39448 20952
rect 39500 20602 39528 21422
rect 39304 20596 39356 20602
rect 39304 20538 39356 20544
rect 39488 20596 39540 20602
rect 39488 20538 39540 20544
rect 39304 20460 39356 20466
rect 39304 20402 39356 20408
rect 39316 20262 39344 20402
rect 39304 20256 39356 20262
rect 39304 20198 39356 20204
rect 39500 19854 39528 20538
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 39488 19712 39540 19718
rect 39488 19654 39540 19660
rect 39500 19378 39528 19654
rect 39304 19372 39356 19378
rect 39304 19314 39356 19320
rect 39488 19372 39540 19378
rect 39488 19314 39540 19320
rect 39316 18970 39344 19314
rect 39592 19145 39620 22578
rect 39684 21593 39712 23666
rect 39776 23594 39804 23666
rect 39856 23656 39908 23662
rect 39856 23598 39908 23604
rect 39764 23588 39816 23594
rect 39764 23530 39816 23536
rect 39764 22704 39816 22710
rect 39764 22646 39816 22652
rect 39776 22030 39804 22646
rect 39868 22094 39896 23598
rect 39960 23118 39988 25638
rect 40052 25294 40080 26318
rect 40132 26240 40184 26246
rect 40132 26182 40184 26188
rect 40144 25906 40172 26182
rect 40132 25900 40184 25906
rect 40132 25842 40184 25848
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40052 24342 40080 25230
rect 40144 25226 40172 25842
rect 40236 25294 40264 26454
rect 41892 26382 41920 26726
rect 41880 26376 41932 26382
rect 41880 26318 41932 26324
rect 41052 26308 41104 26314
rect 41052 26250 41104 26256
rect 41064 26042 41092 26250
rect 41052 26036 41104 26042
rect 41052 25978 41104 25984
rect 41144 25764 41196 25770
rect 41144 25706 41196 25712
rect 41052 25696 41104 25702
rect 41052 25638 41104 25644
rect 41064 25498 41092 25638
rect 41052 25492 41104 25498
rect 41052 25434 41104 25440
rect 40224 25288 40276 25294
rect 40224 25230 40276 25236
rect 40776 25288 40828 25294
rect 40776 25230 40828 25236
rect 40132 25220 40184 25226
rect 40132 25162 40184 25168
rect 40144 24410 40172 25162
rect 40316 25152 40368 25158
rect 40316 25094 40368 25100
rect 40224 24608 40276 24614
rect 40224 24550 40276 24556
rect 40132 24404 40184 24410
rect 40132 24346 40184 24352
rect 40040 24336 40092 24342
rect 40040 24278 40092 24284
rect 40132 24064 40184 24070
rect 40132 24006 40184 24012
rect 40144 23526 40172 24006
rect 40236 23712 40264 24550
rect 40328 24070 40356 25094
rect 40500 24948 40552 24954
rect 40500 24890 40552 24896
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 40316 24064 40368 24070
rect 40316 24006 40368 24012
rect 40236 23684 40356 23712
rect 40132 23520 40184 23526
rect 40132 23462 40184 23468
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 39960 22710 39988 23054
rect 40040 22976 40092 22982
rect 40040 22918 40092 22924
rect 39948 22704 40000 22710
rect 39948 22646 40000 22652
rect 39948 22568 40000 22574
rect 40052 22545 40080 22918
rect 40130 22808 40186 22817
rect 40130 22743 40186 22752
rect 40144 22574 40172 22743
rect 40132 22568 40184 22574
rect 39948 22510 40000 22516
rect 40038 22536 40094 22545
rect 39960 22420 39988 22510
rect 40132 22510 40184 22516
rect 40224 22568 40276 22574
rect 40224 22510 40276 22516
rect 40038 22471 40094 22480
rect 39960 22392 40080 22420
rect 40052 22137 40080 22392
rect 40038 22128 40094 22137
rect 39948 22094 40000 22098
rect 39868 22092 40000 22094
rect 39868 22066 39948 22092
rect 40038 22063 40094 22072
rect 39948 22034 40000 22040
rect 40052 22030 40080 22063
rect 40236 22030 40264 22510
rect 39764 22024 39816 22030
rect 39764 21966 39816 21972
rect 40040 22024 40092 22030
rect 40224 22024 40276 22030
rect 40040 21966 40092 21972
rect 40222 21992 40224 22001
rect 40276 21992 40278 22001
rect 39856 21888 39908 21894
rect 40052 21876 40080 21966
rect 40328 21962 40356 23684
rect 40222 21927 40278 21936
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 40132 21888 40184 21894
rect 40052 21848 40132 21876
rect 39856 21830 39908 21836
rect 40132 21830 40184 21836
rect 39764 21616 39816 21622
rect 39670 21584 39726 21593
rect 39764 21558 39816 21564
rect 39670 21519 39726 21528
rect 39776 19514 39804 21558
rect 39868 21554 39896 21830
rect 40420 21554 40448 24142
rect 39856 21548 39908 21554
rect 39856 21490 39908 21496
rect 40408 21548 40460 21554
rect 40408 21490 40460 21496
rect 40512 21486 40540 24890
rect 40592 24880 40644 24886
rect 40592 24822 40644 24828
rect 40604 23254 40632 24822
rect 40684 24608 40736 24614
rect 40684 24550 40736 24556
rect 40696 24410 40724 24550
rect 40684 24404 40736 24410
rect 40684 24346 40736 24352
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40592 23248 40644 23254
rect 40592 23190 40644 23196
rect 40592 23112 40644 23118
rect 40592 23054 40644 23060
rect 40604 22506 40632 23054
rect 40592 22500 40644 22506
rect 40592 22442 40644 22448
rect 40696 21570 40724 23598
rect 40604 21542 40724 21570
rect 40500 21480 40552 21486
rect 40500 21422 40552 21428
rect 39948 21412 40000 21418
rect 39948 21354 40000 21360
rect 39856 21344 39908 21350
rect 39856 21286 39908 21292
rect 39960 21298 39988 21354
rect 40132 21344 40184 21350
rect 39960 21292 40132 21298
rect 39960 21286 40184 21292
rect 39868 21078 39896 21286
rect 39960 21270 40172 21286
rect 39856 21072 39908 21078
rect 39856 21014 39908 21020
rect 39764 19508 39816 19514
rect 39764 19450 39816 19456
rect 39578 19136 39634 19145
rect 39578 19071 39634 19080
rect 39304 18964 39356 18970
rect 39304 18906 39356 18912
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 39028 18624 39080 18630
rect 39028 18566 39080 18572
rect 39224 18329 39252 18634
rect 39316 18426 39344 18906
rect 39488 18828 39540 18834
rect 39488 18770 39540 18776
rect 39304 18420 39356 18426
rect 39304 18362 39356 18368
rect 39210 18320 39266 18329
rect 39500 18290 39528 18770
rect 39592 18290 39620 19071
rect 39764 18420 39816 18426
rect 39764 18362 39816 18368
rect 39210 18255 39266 18264
rect 39488 18284 39540 18290
rect 39488 18226 39540 18232
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 38844 18216 38896 18222
rect 38844 18158 38896 18164
rect 38856 17678 38884 18158
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 39028 18080 39080 18086
rect 39028 18022 39080 18028
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38948 16794 38976 18022
rect 39040 17270 39068 18022
rect 39120 17672 39172 17678
rect 39120 17614 39172 17620
rect 39028 17264 39080 17270
rect 39028 17206 39080 17212
rect 39132 17134 39160 17614
rect 39212 17536 39264 17542
rect 39212 17478 39264 17484
rect 39486 17504 39542 17513
rect 39120 17128 39172 17134
rect 39120 17070 39172 17076
rect 38936 16788 38988 16794
rect 38936 16730 38988 16736
rect 38844 16720 38896 16726
rect 38844 16662 38896 16668
rect 38856 16590 38884 16662
rect 38844 16584 38896 16590
rect 38844 16526 38896 16532
rect 38936 16584 38988 16590
rect 38936 16526 38988 16532
rect 38844 15360 38896 15366
rect 38844 15302 38896 15308
rect 38856 13394 38884 15302
rect 38948 14822 38976 16526
rect 39120 15904 39172 15910
rect 39120 15846 39172 15852
rect 39028 15020 39080 15026
rect 39028 14962 39080 14968
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 38948 14346 38976 14758
rect 38936 14340 38988 14346
rect 38936 14282 38988 14288
rect 38934 13832 38990 13841
rect 38934 13767 38990 13776
rect 38948 13462 38976 13767
rect 39040 13530 39068 14962
rect 39028 13524 39080 13530
rect 39028 13466 39080 13472
rect 38936 13456 38988 13462
rect 38936 13398 38988 13404
rect 38752 13388 38804 13394
rect 38752 13330 38804 13336
rect 38844 13388 38896 13394
rect 38844 13330 38896 13336
rect 38752 13252 38804 13258
rect 38752 13194 38804 13200
rect 38936 13252 38988 13258
rect 38936 13194 38988 13200
rect 38764 12986 38792 13194
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38752 12980 38804 12986
rect 38752 12922 38804 12928
rect 38948 12918 38976 13194
rect 38936 12912 38988 12918
rect 38936 12854 38988 12860
rect 39132 12374 39160 15846
rect 39224 14521 39252 17478
rect 39486 17439 39542 17448
rect 39500 17338 39528 17439
rect 39396 17332 39448 17338
rect 39396 17274 39448 17280
rect 39488 17332 39540 17338
rect 39488 17274 39540 17280
rect 39304 17196 39356 17202
rect 39408 17184 39436 17274
rect 39580 17196 39632 17202
rect 39408 17156 39580 17184
rect 39304 17138 39356 17144
rect 39580 17138 39632 17144
rect 39316 16794 39344 17138
rect 39304 16788 39356 16794
rect 39304 16730 39356 16736
rect 39488 16652 39540 16658
rect 39488 16594 39540 16600
rect 39302 16144 39358 16153
rect 39500 16114 39528 16594
rect 39302 16079 39304 16088
rect 39356 16079 39358 16088
rect 39488 16108 39540 16114
rect 39304 16050 39356 16056
rect 39488 16050 39540 16056
rect 39580 16040 39632 16046
rect 39580 15982 39632 15988
rect 39592 15026 39620 15982
rect 39776 15910 39804 18362
rect 39764 15904 39816 15910
rect 39764 15846 39816 15852
rect 39776 15065 39804 15846
rect 39762 15056 39818 15065
rect 39304 15020 39356 15026
rect 39304 14962 39356 14968
rect 39580 15020 39632 15026
rect 39762 14991 39818 15000
rect 39580 14962 39632 14968
rect 39316 14822 39344 14962
rect 39486 14920 39542 14929
rect 39486 14855 39542 14864
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 39304 14612 39356 14618
rect 39304 14554 39356 14560
rect 39210 14512 39266 14521
rect 39210 14447 39266 14456
rect 39212 14340 39264 14346
rect 39212 14282 39264 14288
rect 39224 14006 39252 14282
rect 39212 14000 39264 14006
rect 39212 13942 39264 13948
rect 39316 13734 39344 14554
rect 39500 14482 39528 14855
rect 39592 14618 39620 14962
rect 39672 14952 39724 14958
rect 39672 14894 39724 14900
rect 39580 14612 39632 14618
rect 39580 14554 39632 14560
rect 39488 14476 39540 14482
rect 39488 14418 39540 14424
rect 39684 13977 39712 14894
rect 39868 14618 39896 21014
rect 39960 20806 39988 21270
rect 40512 21078 40540 21422
rect 40604 21146 40632 21542
rect 40788 21350 40816 25230
rect 40868 25152 40920 25158
rect 40868 25094 40920 25100
rect 40880 24274 40908 25094
rect 41064 24954 41092 25434
rect 41156 25430 41184 25706
rect 41144 25424 41196 25430
rect 41144 25366 41196 25372
rect 41052 24948 41104 24954
rect 41052 24890 41104 24896
rect 40960 24812 41012 24818
rect 40960 24754 41012 24760
rect 40972 24274 41000 24754
rect 41156 24342 41184 25366
rect 41236 25288 41288 25294
rect 41236 25230 41288 25236
rect 41248 24750 41276 25230
rect 41696 24948 41748 24954
rect 41696 24890 41748 24896
rect 41604 24812 41656 24818
rect 41604 24754 41656 24760
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 41512 24744 41564 24750
rect 41512 24686 41564 24692
rect 41144 24336 41196 24342
rect 41144 24278 41196 24284
rect 40868 24268 40920 24274
rect 40868 24210 40920 24216
rect 40960 24268 41012 24274
rect 40960 24210 41012 24216
rect 41156 23730 41184 24278
rect 41524 24206 41552 24686
rect 41616 24449 41644 24754
rect 41602 24440 41658 24449
rect 41602 24375 41658 24384
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 41236 24064 41288 24070
rect 41236 24006 41288 24012
rect 41144 23724 41196 23730
rect 41144 23666 41196 23672
rect 40868 23520 40920 23526
rect 41248 23497 41276 24006
rect 41524 23866 41552 24142
rect 41616 24070 41644 24375
rect 41708 24184 41736 24890
rect 41696 24178 41748 24184
rect 41696 24120 41748 24126
rect 41604 24064 41656 24070
rect 41604 24006 41656 24012
rect 41512 23860 41564 23866
rect 41512 23802 41564 23808
rect 41892 23769 41920 26318
rect 43444 26308 43496 26314
rect 43444 26250 43496 26256
rect 42800 25968 42852 25974
rect 42800 25910 42852 25916
rect 42064 25900 42116 25906
rect 42064 25842 42116 25848
rect 41972 25696 42024 25702
rect 41972 25638 42024 25644
rect 41984 25294 42012 25638
rect 41972 25288 42024 25294
rect 41972 25230 42024 25236
rect 42076 24206 42104 25842
rect 42432 25288 42484 25294
rect 42432 25230 42484 25236
rect 42156 25152 42208 25158
rect 42156 25094 42208 25100
rect 42168 24954 42196 25094
rect 42156 24948 42208 24954
rect 42156 24890 42208 24896
rect 42444 24886 42472 25230
rect 42432 24880 42484 24886
rect 42432 24822 42484 24828
rect 42616 24676 42668 24682
rect 42616 24618 42668 24624
rect 42248 24404 42300 24410
rect 42248 24346 42300 24352
rect 41972 24200 42024 24206
rect 41972 24142 42024 24148
rect 42064 24200 42116 24206
rect 42064 24142 42116 24148
rect 41878 23760 41934 23769
rect 41878 23695 41934 23704
rect 41512 23520 41564 23526
rect 40868 23462 40920 23468
rect 41234 23488 41290 23497
rect 40880 23118 40908 23462
rect 41512 23462 41564 23468
rect 41234 23423 41290 23432
rect 40868 23112 40920 23118
rect 41236 23112 41288 23118
rect 40868 23054 40920 23060
rect 41234 23080 41236 23089
rect 41420 23112 41472 23118
rect 41288 23080 41290 23089
rect 41144 23044 41196 23050
rect 41420 23054 41472 23060
rect 41234 23015 41290 23024
rect 41144 22986 41196 22992
rect 40960 22976 41012 22982
rect 40960 22918 41012 22924
rect 40868 22704 40920 22710
rect 40866 22672 40868 22681
rect 40920 22672 40922 22681
rect 40866 22607 40922 22616
rect 40972 22098 41000 22918
rect 41156 22778 41184 22986
rect 41144 22772 41196 22778
rect 41144 22714 41196 22720
rect 41144 22636 41196 22642
rect 41432 22624 41460 23054
rect 41196 22596 41460 22624
rect 41144 22578 41196 22584
rect 41052 22500 41104 22506
rect 41052 22442 41104 22448
rect 40960 22092 41012 22098
rect 40960 22034 41012 22040
rect 40960 21956 41012 21962
rect 40960 21898 41012 21904
rect 40868 21548 40920 21554
rect 40868 21490 40920 21496
rect 40776 21344 40828 21350
rect 40776 21286 40828 21292
rect 40592 21140 40644 21146
rect 40592 21082 40644 21088
rect 40500 21072 40552 21078
rect 40500 21014 40552 21020
rect 40040 20868 40092 20874
rect 40040 20810 40092 20816
rect 39948 20800 40000 20806
rect 39948 20742 40000 20748
rect 39960 20466 39988 20742
rect 39948 20460 40000 20466
rect 39948 20402 40000 20408
rect 39960 17678 39988 20402
rect 40052 19854 40080 20810
rect 40500 20800 40552 20806
rect 40498 20768 40500 20777
rect 40552 20768 40554 20777
rect 40498 20703 40554 20712
rect 40144 20590 40540 20618
rect 40144 20262 40172 20590
rect 40512 20534 40540 20590
rect 40224 20528 40276 20534
rect 40224 20470 40276 20476
rect 40500 20528 40552 20534
rect 40500 20470 40552 20476
rect 40236 20330 40264 20470
rect 40604 20346 40632 21082
rect 40880 20641 40908 21490
rect 40866 20632 40922 20641
rect 40684 20596 40736 20602
rect 40866 20567 40922 20576
rect 40684 20538 40736 20544
rect 40224 20324 40276 20330
rect 40420 20318 40632 20346
rect 40276 20284 40356 20312
rect 40224 20266 40276 20272
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 40040 19848 40092 19854
rect 40040 19790 40092 19796
rect 40144 19334 40172 20198
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40236 19446 40264 19790
rect 40224 19440 40276 19446
rect 40224 19382 40276 19388
rect 40328 19378 40356 20284
rect 40316 19372 40368 19378
rect 40144 19306 40264 19334
rect 40316 19314 40368 19320
rect 40130 18320 40186 18329
rect 40130 18255 40186 18264
rect 40144 17678 40172 18255
rect 39948 17672 40000 17678
rect 40132 17672 40184 17678
rect 40000 17632 40080 17660
rect 39948 17614 40000 17620
rect 40052 16998 40080 17632
rect 40132 17614 40184 17620
rect 40236 17610 40264 19306
rect 40420 18426 40448 20318
rect 40592 20256 40644 20262
rect 40592 20198 40644 20204
rect 40604 19854 40632 20198
rect 40696 19990 40724 20538
rect 40868 20460 40920 20466
rect 40868 20402 40920 20408
rect 40776 20052 40828 20058
rect 40776 19994 40828 20000
rect 40684 19984 40736 19990
rect 40684 19926 40736 19932
rect 40500 19848 40552 19854
rect 40500 19790 40552 19796
rect 40592 19848 40644 19854
rect 40592 19790 40644 19796
rect 40512 19514 40540 19790
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40684 19508 40736 19514
rect 40684 19450 40736 19456
rect 40500 18692 40552 18698
rect 40500 18634 40552 18640
rect 40408 18420 40460 18426
rect 40408 18362 40460 18368
rect 40512 18306 40540 18634
rect 40592 18420 40644 18426
rect 40592 18362 40644 18368
rect 40420 18278 40540 18306
rect 40316 18216 40368 18222
rect 40316 18158 40368 18164
rect 40224 17604 40276 17610
rect 40224 17546 40276 17552
rect 40328 17542 40356 18158
rect 40316 17536 40368 17542
rect 40316 17478 40368 17484
rect 40132 17060 40184 17066
rect 40132 17002 40184 17008
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40052 15450 40080 16934
rect 40144 16590 40172 17002
rect 40328 16658 40356 17478
rect 40420 17116 40448 18278
rect 40500 17740 40552 17746
rect 40500 17682 40552 17688
rect 40512 17270 40540 17682
rect 40500 17264 40552 17270
rect 40500 17206 40552 17212
rect 40420 17088 40540 17116
rect 40408 16992 40460 16998
rect 40408 16934 40460 16940
rect 40316 16652 40368 16658
rect 40316 16594 40368 16600
rect 40132 16584 40184 16590
rect 40132 16526 40184 16532
rect 40316 16176 40368 16182
rect 40316 16118 40368 16124
rect 40222 15736 40278 15745
rect 40222 15671 40224 15680
rect 40276 15671 40278 15680
rect 40224 15642 40276 15648
rect 40132 15564 40184 15570
rect 40132 15506 40184 15512
rect 39960 15422 40080 15450
rect 39960 14906 39988 15422
rect 40040 15360 40092 15366
rect 40040 15302 40092 15308
rect 40052 15026 40080 15302
rect 40040 15020 40092 15026
rect 40040 14962 40092 14968
rect 39960 14878 40080 14906
rect 39856 14612 39908 14618
rect 39856 14554 39908 14560
rect 39868 14385 39896 14554
rect 39854 14376 39910 14385
rect 39854 14311 39910 14320
rect 39670 13968 39726 13977
rect 39670 13903 39726 13912
rect 39304 13728 39356 13734
rect 39304 13670 39356 13676
rect 40052 13530 40080 14878
rect 40040 13524 40092 13530
rect 40040 13466 40092 13472
rect 39212 13456 39264 13462
rect 39212 13398 39264 13404
rect 39120 12368 39172 12374
rect 39120 12310 39172 12316
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38212 11354 38240 11698
rect 39132 11558 39160 12310
rect 39224 12238 39252 13398
rect 40144 13190 40172 15506
rect 40236 15201 40264 15642
rect 40328 15570 40356 16118
rect 40420 16114 40448 16934
rect 40512 16590 40540 17088
rect 40500 16584 40552 16590
rect 40500 16526 40552 16532
rect 40512 16425 40540 16526
rect 40498 16416 40554 16425
rect 40498 16351 40554 16360
rect 40500 16244 40552 16250
rect 40500 16186 40552 16192
rect 40408 16108 40460 16114
rect 40408 16050 40460 16056
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 40222 15192 40278 15201
rect 40222 15127 40278 15136
rect 40222 15056 40278 15065
rect 40222 14991 40278 15000
rect 40236 14958 40264 14991
rect 40224 14952 40276 14958
rect 40408 14952 40460 14958
rect 40224 14894 40276 14900
rect 40328 14912 40408 14940
rect 40328 14074 40356 14912
rect 40408 14894 40460 14900
rect 40316 14068 40368 14074
rect 40316 14010 40368 14016
rect 40406 13968 40462 13977
rect 40406 13903 40462 13912
rect 40316 13864 40368 13870
rect 40316 13806 40368 13812
rect 40328 13569 40356 13806
rect 40314 13560 40370 13569
rect 40314 13495 40370 13504
rect 40316 13320 40368 13326
rect 40316 13262 40368 13268
rect 39672 13184 39724 13190
rect 39672 13126 39724 13132
rect 40132 13184 40184 13190
rect 40132 13126 40184 13132
rect 39684 12850 39712 13126
rect 40328 12986 40356 13262
rect 40420 13258 40448 13903
rect 40512 13394 40540 16186
rect 40500 13388 40552 13394
rect 40500 13330 40552 13336
rect 40408 13252 40460 13258
rect 40408 13194 40460 13200
rect 40500 13184 40552 13190
rect 40500 13126 40552 13132
rect 40512 12986 40540 13126
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40500 12980 40552 12986
rect 40500 12922 40552 12928
rect 39672 12844 39724 12850
rect 39672 12786 39724 12792
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 39224 11762 39252 12174
rect 40604 11830 40632 18362
rect 40696 17882 40724 19450
rect 40788 18766 40816 19994
rect 40880 19825 40908 20402
rect 40866 19816 40922 19825
rect 40866 19751 40922 19760
rect 40868 19372 40920 19378
rect 40972 19360 41000 21898
rect 41064 21570 41092 22442
rect 41156 22030 41184 22578
rect 41144 22024 41196 22030
rect 41144 21966 41196 21972
rect 41236 21888 41288 21894
rect 41236 21830 41288 21836
rect 41064 21542 41184 21570
rect 41052 21412 41104 21418
rect 41052 21354 41104 21360
rect 41064 20466 41092 21354
rect 41156 20602 41184 21542
rect 41248 21146 41276 21830
rect 41326 21584 41382 21593
rect 41326 21519 41328 21528
rect 41380 21519 41382 21528
rect 41328 21490 41380 21496
rect 41236 21140 41288 21146
rect 41236 21082 41288 21088
rect 41144 20596 41196 20602
rect 41144 20538 41196 20544
rect 41052 20460 41104 20466
rect 41052 20402 41104 20408
rect 41064 20330 41092 20402
rect 41248 20398 41276 21082
rect 41236 20392 41288 20398
rect 41236 20334 41288 20340
rect 41052 20324 41104 20330
rect 41052 20266 41104 20272
rect 41144 20256 41196 20262
rect 41144 20198 41196 20204
rect 41156 19922 41184 20198
rect 41144 19916 41196 19922
rect 41144 19858 41196 19864
rect 40920 19332 41000 19360
rect 40868 19314 40920 19320
rect 40776 18760 40828 18766
rect 40776 18702 40828 18708
rect 40684 17876 40736 17882
rect 40684 17818 40736 17824
rect 40696 17202 40724 17818
rect 40776 17332 40828 17338
rect 40776 17274 40828 17280
rect 40684 17196 40736 17202
rect 40684 17138 40736 17144
rect 40788 16658 40816 17274
rect 40776 16652 40828 16658
rect 40776 16594 40828 16600
rect 40788 16250 40816 16594
rect 40776 16244 40828 16250
rect 40776 16186 40828 16192
rect 40880 16182 40908 19314
rect 41052 19236 41104 19242
rect 41052 19178 41104 19184
rect 41064 18766 41092 19178
rect 41156 18902 41184 19858
rect 41524 19854 41552 23462
rect 41788 23044 41840 23050
rect 41788 22986 41840 22992
rect 41800 22642 41828 22986
rect 41788 22636 41840 22642
rect 41788 22578 41840 22584
rect 41696 22500 41748 22506
rect 41748 22460 41828 22488
rect 41696 22442 41748 22448
rect 41800 22166 41828 22460
rect 41696 22160 41748 22166
rect 41696 22102 41748 22108
rect 41788 22160 41840 22166
rect 41788 22102 41840 22108
rect 41602 21856 41658 21865
rect 41602 21791 41658 21800
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 41328 19712 41380 19718
rect 41328 19654 41380 19660
rect 41144 18896 41196 18902
rect 41144 18838 41196 18844
rect 41052 18760 41104 18766
rect 41052 18702 41104 18708
rect 41064 17762 41092 18702
rect 41340 18290 41368 19654
rect 41420 19304 41472 19310
rect 41420 19246 41472 19252
rect 41512 19304 41564 19310
rect 41512 19246 41564 19252
rect 41432 18714 41460 19246
rect 41524 18970 41552 19246
rect 41512 18964 41564 18970
rect 41512 18906 41564 18912
rect 41432 18686 41552 18714
rect 41524 18630 41552 18686
rect 41512 18624 41564 18630
rect 41512 18566 41564 18572
rect 41328 18284 41380 18290
rect 41328 18226 41380 18232
rect 41512 18216 41564 18222
rect 41512 18158 41564 18164
rect 41234 18048 41290 18057
rect 41234 17983 41290 17992
rect 40972 17734 41092 17762
rect 40972 17202 41000 17734
rect 41248 17678 41276 17983
rect 41524 17882 41552 18158
rect 41616 17954 41644 21791
rect 41708 21418 41736 22102
rect 41984 22098 42012 24142
rect 42076 23662 42104 24142
rect 42064 23656 42116 23662
rect 42064 23598 42116 23604
rect 41972 22092 42024 22098
rect 41972 22034 42024 22040
rect 41984 21622 42012 22034
rect 41972 21616 42024 21622
rect 41972 21558 42024 21564
rect 41696 21412 41748 21418
rect 41696 21354 41748 21360
rect 41984 21010 42012 21558
rect 41972 21004 42024 21010
rect 41972 20946 42024 20952
rect 41984 20602 42012 20946
rect 42156 20800 42208 20806
rect 42156 20742 42208 20748
rect 41788 20596 41840 20602
rect 41788 20538 41840 20544
rect 41972 20596 42024 20602
rect 41972 20538 42024 20544
rect 41696 20256 41748 20262
rect 41696 20198 41748 20204
rect 41708 19990 41736 20198
rect 41696 19984 41748 19990
rect 41696 19926 41748 19932
rect 41800 19854 41828 20538
rect 41880 20460 41932 20466
rect 41880 20402 41932 20408
rect 41892 19990 41920 20402
rect 42064 20392 42116 20398
rect 42064 20334 42116 20340
rect 41970 20088 42026 20097
rect 41970 20023 41972 20032
rect 42024 20023 42026 20032
rect 41972 19994 42024 20000
rect 41880 19984 41932 19990
rect 41880 19926 41932 19932
rect 41984 19854 42012 19994
rect 41788 19848 41840 19854
rect 41788 19790 41840 19796
rect 41972 19848 42024 19854
rect 41972 19790 42024 19796
rect 41696 19712 41748 19718
rect 41696 19654 41748 19660
rect 41708 18873 41736 19654
rect 42076 19446 42104 20334
rect 42064 19440 42116 19446
rect 42064 19382 42116 19388
rect 41880 19372 41932 19378
rect 41880 19314 41932 19320
rect 41788 19304 41840 19310
rect 41788 19246 41840 19252
rect 41800 19174 41828 19246
rect 41788 19168 41840 19174
rect 41788 19110 41840 19116
rect 41694 18864 41750 18873
rect 41892 18834 41920 19314
rect 41694 18799 41750 18808
rect 41880 18828 41932 18834
rect 41880 18770 41932 18776
rect 41616 17926 41736 17954
rect 41512 17876 41564 17882
rect 41512 17818 41564 17824
rect 41708 17814 41736 17926
rect 42076 17882 42104 19382
rect 42064 17876 42116 17882
rect 42064 17818 42116 17824
rect 41696 17808 41748 17814
rect 41696 17750 41748 17756
rect 41420 17740 41472 17746
rect 41420 17682 41472 17688
rect 41512 17740 41564 17746
rect 41512 17682 41564 17688
rect 41236 17672 41288 17678
rect 41432 17649 41460 17682
rect 41236 17614 41288 17620
rect 41418 17640 41474 17649
rect 41418 17575 41474 17584
rect 41524 17338 41552 17682
rect 41512 17332 41564 17338
rect 41512 17274 41564 17280
rect 40960 17196 41012 17202
rect 40960 17138 41012 17144
rect 41328 17196 41380 17202
rect 41328 17138 41380 17144
rect 41340 16998 41368 17138
rect 41420 17060 41472 17066
rect 41420 17002 41472 17008
rect 40960 16992 41012 16998
rect 40960 16934 41012 16940
rect 41328 16992 41380 16998
rect 41328 16934 41380 16940
rect 40868 16176 40920 16182
rect 40868 16118 40920 16124
rect 40868 16040 40920 16046
rect 40868 15982 40920 15988
rect 40776 15904 40828 15910
rect 40776 15846 40828 15852
rect 40682 15192 40738 15201
rect 40682 15127 40738 15136
rect 40696 15026 40724 15127
rect 40684 15020 40736 15026
rect 40684 14962 40736 14968
rect 40684 14476 40736 14482
rect 40684 14418 40736 14424
rect 40696 14113 40724 14418
rect 40682 14104 40738 14113
rect 40788 14074 40816 15846
rect 40880 14929 40908 15982
rect 40972 15978 41000 16934
rect 41340 16794 41368 16934
rect 41328 16788 41380 16794
rect 41328 16730 41380 16736
rect 41432 16640 41460 17002
rect 41340 16612 41460 16640
rect 41236 16584 41288 16590
rect 41234 16552 41236 16561
rect 41288 16552 41290 16561
rect 41234 16487 41290 16496
rect 40960 15972 41012 15978
rect 40960 15914 41012 15920
rect 41144 15700 41196 15706
rect 41144 15642 41196 15648
rect 41156 15502 41184 15642
rect 41144 15496 41196 15502
rect 41144 15438 41196 15444
rect 40866 14920 40922 14929
rect 40866 14855 40922 14864
rect 41052 14816 41104 14822
rect 41052 14758 41104 14764
rect 41064 14414 41092 14758
rect 40960 14408 41012 14414
rect 40880 14368 40960 14396
rect 40682 14039 40738 14048
rect 40776 14068 40828 14074
rect 40776 14010 40828 14016
rect 40684 13932 40736 13938
rect 40684 13874 40736 13880
rect 40696 13841 40724 13874
rect 40682 13832 40738 13841
rect 40682 13767 40738 13776
rect 40788 13530 40816 14010
rect 40776 13524 40828 13530
rect 40776 13466 40828 13472
rect 40776 13320 40828 13326
rect 40776 13262 40828 13268
rect 40788 12442 40816 13262
rect 40880 12918 40908 14368
rect 40960 14350 41012 14356
rect 41052 14408 41104 14414
rect 41052 14350 41104 14356
rect 41340 14278 41368 16612
rect 41708 16590 41736 17750
rect 41972 17536 42024 17542
rect 41972 17478 42024 17484
rect 41984 17066 42012 17478
rect 42076 17338 42104 17818
rect 42064 17332 42116 17338
rect 42064 17274 42116 17280
rect 41972 17060 42024 17066
rect 41972 17002 42024 17008
rect 41696 16584 41748 16590
rect 41696 16526 41748 16532
rect 41420 16516 41472 16522
rect 41420 16458 41472 16464
rect 41432 16114 41460 16458
rect 41512 16244 41564 16250
rect 41512 16186 41564 16192
rect 41420 16108 41472 16114
rect 41420 16050 41472 16056
rect 41524 15094 41552 16186
rect 41512 15088 41564 15094
rect 41512 15030 41564 15036
rect 41602 15056 41658 15065
rect 41524 14396 41552 15030
rect 41602 14991 41604 15000
rect 41656 14991 41658 15000
rect 41604 14962 41656 14968
rect 41708 14822 41736 16526
rect 41880 16108 41932 16114
rect 41880 16050 41932 16056
rect 41892 16017 41920 16050
rect 41878 16008 41934 16017
rect 41878 15943 41934 15952
rect 42076 15706 42104 17274
rect 42064 15700 42116 15706
rect 42064 15642 42116 15648
rect 41788 15020 41840 15026
rect 41788 14962 41840 14968
rect 41800 14929 41828 14962
rect 41972 14952 42024 14958
rect 41786 14920 41842 14929
rect 41972 14894 42024 14900
rect 41786 14855 41842 14864
rect 41696 14816 41748 14822
rect 41696 14758 41748 14764
rect 41984 14482 42012 14894
rect 41972 14476 42024 14482
rect 41972 14418 42024 14424
rect 41604 14408 41656 14414
rect 41524 14368 41604 14396
rect 41604 14350 41656 14356
rect 41328 14272 41380 14278
rect 40958 14240 41014 14249
rect 41328 14214 41380 14220
rect 40958 14175 41014 14184
rect 40972 13938 41000 14175
rect 41144 14000 41196 14006
rect 41144 13942 41196 13948
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 40972 13326 41000 13874
rect 41156 13870 41184 13942
rect 41340 13938 41368 14214
rect 42076 14074 42104 15642
rect 42168 15026 42196 20742
rect 42260 20466 42288 24346
rect 42628 24274 42656 24618
rect 42616 24268 42668 24274
rect 42668 24228 42748 24256
rect 42616 24210 42668 24216
rect 42616 24064 42668 24070
rect 42616 24006 42668 24012
rect 42432 23860 42484 23866
rect 42432 23802 42484 23808
rect 42340 22636 42392 22642
rect 42340 22578 42392 22584
rect 42248 20460 42300 20466
rect 42248 20402 42300 20408
rect 42352 20074 42380 22578
rect 42444 20788 42472 23802
rect 42628 22817 42656 24006
rect 42720 23662 42748 24228
rect 42708 23656 42760 23662
rect 42708 23598 42760 23604
rect 42720 23118 42748 23598
rect 42708 23112 42760 23118
rect 42708 23054 42760 23060
rect 42812 22930 42840 25910
rect 43456 25906 43484 26250
rect 43628 25968 43680 25974
rect 43628 25910 43680 25916
rect 43444 25900 43496 25906
rect 43444 25842 43496 25848
rect 43536 25900 43588 25906
rect 43536 25842 43588 25848
rect 43352 25696 43404 25702
rect 43352 25638 43404 25644
rect 43364 25294 43392 25638
rect 43456 25362 43484 25842
rect 43444 25356 43496 25362
rect 43444 25298 43496 25304
rect 43352 25288 43404 25294
rect 43352 25230 43404 25236
rect 42984 25220 43036 25226
rect 42984 25162 43036 25168
rect 42996 24954 43024 25162
rect 43352 25152 43404 25158
rect 43352 25094 43404 25100
rect 42984 24948 43036 24954
rect 42984 24890 43036 24896
rect 43364 23866 43392 25094
rect 43456 24682 43484 25298
rect 43548 24886 43576 25842
rect 43536 24880 43588 24886
rect 43536 24822 43588 24828
rect 43640 24818 43668 25910
rect 44008 25430 44036 26862
rect 44824 26240 44876 26246
rect 44824 26182 44876 26188
rect 44836 25906 44864 26182
rect 44824 25900 44876 25906
rect 44824 25842 44876 25848
rect 46112 25900 46164 25906
rect 46112 25842 46164 25848
rect 43996 25424 44048 25430
rect 43996 25366 44048 25372
rect 43904 25288 43956 25294
rect 43904 25230 43956 25236
rect 43812 25220 43864 25226
rect 43812 25162 43864 25168
rect 43628 24812 43680 24818
rect 43628 24754 43680 24760
rect 43444 24676 43496 24682
rect 43444 24618 43496 24624
rect 43536 24132 43588 24138
rect 43536 24074 43588 24080
rect 43352 23860 43404 23866
rect 43352 23802 43404 23808
rect 43548 23798 43576 24074
rect 43536 23792 43588 23798
rect 43536 23734 43588 23740
rect 43640 23730 43668 24754
rect 43824 24614 43852 25162
rect 43812 24608 43864 24614
rect 43812 24550 43864 24556
rect 43824 23798 43852 24550
rect 43812 23792 43864 23798
rect 43812 23734 43864 23740
rect 43168 23724 43220 23730
rect 43168 23666 43220 23672
rect 43444 23724 43496 23730
rect 43444 23666 43496 23672
rect 43628 23724 43680 23730
rect 43628 23666 43680 23672
rect 42984 23520 43036 23526
rect 42984 23462 43036 23468
rect 42996 23186 43024 23462
rect 42984 23180 43036 23186
rect 42984 23122 43036 23128
rect 42812 22902 42932 22930
rect 42614 22808 42670 22817
rect 42614 22743 42670 22752
rect 42628 22574 42656 22743
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 42800 22568 42852 22574
rect 42800 22510 42852 22516
rect 42812 22030 42840 22510
rect 42800 22024 42852 22030
rect 42720 21984 42800 22012
rect 42720 21842 42748 21984
rect 42800 21966 42852 21972
rect 42904 21978 42932 22902
rect 42996 22710 43024 23122
rect 43180 22982 43208 23666
rect 43352 23248 43404 23254
rect 43352 23190 43404 23196
rect 43168 22976 43220 22982
rect 43168 22918 43220 22924
rect 43364 22710 43392 23190
rect 42984 22704 43036 22710
rect 42984 22646 43036 22652
rect 43352 22704 43404 22710
rect 43352 22646 43404 22652
rect 43076 22432 43128 22438
rect 43076 22374 43128 22380
rect 43088 22273 43116 22374
rect 43074 22264 43130 22273
rect 43074 22199 43130 22208
rect 43168 22228 43220 22234
rect 43168 22170 43220 22176
rect 43180 22001 43208 22170
rect 43352 22024 43404 22030
rect 43166 21992 43222 22001
rect 42904 21962 43116 21978
rect 42904 21956 43128 21962
rect 42904 21950 43076 21956
rect 43352 21966 43404 21972
rect 43166 21927 43222 21936
rect 43076 21898 43128 21904
rect 42720 21814 43024 21842
rect 42708 21344 42760 21350
rect 42708 21286 42760 21292
rect 42892 21344 42944 21350
rect 42892 21286 42944 21292
rect 42720 21146 42748 21286
rect 42708 21140 42760 21146
rect 42708 21082 42760 21088
rect 42524 20936 42576 20942
rect 42904 20924 42932 21286
rect 42576 20896 42932 20924
rect 42524 20878 42576 20884
rect 42524 20800 42576 20806
rect 42444 20760 42524 20788
rect 42524 20742 42576 20748
rect 42800 20800 42852 20806
rect 42800 20742 42852 20748
rect 42432 20460 42484 20466
rect 42432 20402 42484 20408
rect 42260 20046 42380 20074
rect 42260 19145 42288 20046
rect 42340 19984 42392 19990
rect 42340 19926 42392 19932
rect 42246 19136 42302 19145
rect 42246 19071 42302 19080
rect 42260 16590 42288 19071
rect 42248 16584 42300 16590
rect 42248 16526 42300 16532
rect 42156 15020 42208 15026
rect 42156 14962 42208 14968
rect 42156 14816 42208 14822
rect 42156 14758 42208 14764
rect 42168 14482 42196 14758
rect 42156 14476 42208 14482
rect 42156 14418 42208 14424
rect 41880 14068 41932 14074
rect 41880 14010 41932 14016
rect 42064 14068 42116 14074
rect 42064 14010 42116 14016
rect 41328 13932 41380 13938
rect 41328 13874 41380 13880
rect 41144 13864 41196 13870
rect 41144 13806 41196 13812
rect 40960 13320 41012 13326
rect 40960 13262 41012 13268
rect 41052 13252 41104 13258
rect 41052 13194 41104 13200
rect 40868 12912 40920 12918
rect 40868 12854 40920 12860
rect 40960 12844 41012 12850
rect 41064 12832 41092 13194
rect 41156 12918 41184 13806
rect 41236 13728 41288 13734
rect 41236 13670 41288 13676
rect 41512 13728 41564 13734
rect 41512 13670 41564 13676
rect 41144 12912 41196 12918
rect 41144 12854 41196 12860
rect 41248 12850 41276 13670
rect 41524 12850 41552 13670
rect 41892 13326 41920 14010
rect 41970 13968 42026 13977
rect 41970 13903 41972 13912
rect 42024 13903 42026 13912
rect 41972 13874 42024 13880
rect 42156 13728 42208 13734
rect 42156 13670 42208 13676
rect 42062 13560 42118 13569
rect 42062 13495 42118 13504
rect 42076 13394 42104 13495
rect 42064 13388 42116 13394
rect 42064 13330 42116 13336
rect 42168 13326 42196 13670
rect 41880 13320 41932 13326
rect 41880 13262 41932 13268
rect 42156 13320 42208 13326
rect 42156 13262 42208 13268
rect 41892 12918 41920 13262
rect 42260 13190 42288 16526
rect 42352 16522 42380 19926
rect 42444 19378 42472 20402
rect 42432 19372 42484 19378
rect 42432 19314 42484 19320
rect 42432 18964 42484 18970
rect 42432 18906 42484 18912
rect 42444 17678 42472 18906
rect 42536 18698 42564 20742
rect 42616 19848 42668 19854
rect 42616 19790 42668 19796
rect 42524 18692 42576 18698
rect 42524 18634 42576 18640
rect 42536 18222 42564 18634
rect 42524 18216 42576 18222
rect 42524 18158 42576 18164
rect 42524 17876 42576 17882
rect 42524 17818 42576 17824
rect 42432 17672 42484 17678
rect 42432 17614 42484 17620
rect 42536 17610 42564 17818
rect 42628 17610 42656 19790
rect 42708 19372 42760 19378
rect 42708 19314 42760 19320
rect 42720 17678 42748 19314
rect 42812 18834 42840 20742
rect 42904 20466 42932 20896
rect 42892 20460 42944 20466
rect 42892 20402 42944 20408
rect 42904 19786 42932 20402
rect 42892 19780 42944 19786
rect 42892 19722 42944 19728
rect 42800 18828 42852 18834
rect 42800 18770 42852 18776
rect 42800 18420 42852 18426
rect 42800 18362 42852 18368
rect 42812 17814 42840 18362
rect 42904 18290 42932 19722
rect 42996 18358 43024 21814
rect 43088 19514 43116 21898
rect 43076 19508 43128 19514
rect 43076 19450 43128 19456
rect 43180 19446 43208 21927
rect 43260 21548 43312 21554
rect 43260 21490 43312 21496
rect 43272 21418 43300 21490
rect 43260 21412 43312 21418
rect 43260 21354 43312 21360
rect 43364 20466 43392 21966
rect 43456 20602 43484 23666
rect 43536 23520 43588 23526
rect 43536 23462 43588 23468
rect 43548 23254 43576 23462
rect 43536 23248 43588 23254
rect 43536 23190 43588 23196
rect 43548 21622 43576 23190
rect 43824 23050 43852 23734
rect 43916 23089 43944 25230
rect 44008 24410 44036 25366
rect 44836 24818 44864 25842
rect 46124 25294 46152 25842
rect 46112 25288 46164 25294
rect 46112 25230 46164 25236
rect 45468 25220 45520 25226
rect 45468 25162 45520 25168
rect 45480 24886 45508 25162
rect 45468 24880 45520 24886
rect 45388 24840 45468 24868
rect 44272 24812 44324 24818
rect 44272 24754 44324 24760
rect 44824 24812 44876 24818
rect 44876 24772 44956 24800
rect 44824 24754 44876 24760
rect 44088 24676 44140 24682
rect 44088 24618 44140 24624
rect 43996 24404 44048 24410
rect 43996 24346 44048 24352
rect 44008 24206 44036 24346
rect 43996 24200 44048 24206
rect 43996 24142 44048 24148
rect 43902 23080 43958 23089
rect 43812 23044 43864 23050
rect 43902 23015 43958 23024
rect 43812 22986 43864 22992
rect 43628 22976 43680 22982
rect 43628 22918 43680 22924
rect 43640 22098 43668 22918
rect 43628 22092 43680 22098
rect 43628 22034 43680 22040
rect 43720 21956 43772 21962
rect 43720 21898 43772 21904
rect 43536 21616 43588 21622
rect 43536 21558 43588 21564
rect 43548 21010 43576 21558
rect 43732 21486 43760 21898
rect 43824 21554 43852 22986
rect 43916 22964 43944 23015
rect 43996 22976 44048 22982
rect 43916 22936 43996 22964
rect 43996 22918 44048 22924
rect 44008 22438 44036 22918
rect 44100 22574 44128 24618
rect 44284 24274 44312 24754
rect 44272 24268 44324 24274
rect 44272 24210 44324 24216
rect 44180 24132 44232 24138
rect 44180 24074 44232 24080
rect 44192 23730 44220 24074
rect 44180 23724 44232 23730
rect 44180 23666 44232 23672
rect 44088 22568 44140 22574
rect 44088 22510 44140 22516
rect 43996 22432 44048 22438
rect 43996 22374 44048 22380
rect 44008 22030 44036 22374
rect 43996 22024 44048 22030
rect 43996 21966 44048 21972
rect 43812 21548 43864 21554
rect 43812 21490 43864 21496
rect 43720 21480 43772 21486
rect 43720 21422 43772 21428
rect 43628 21412 43680 21418
rect 43628 21354 43680 21360
rect 43536 21004 43588 21010
rect 43536 20946 43588 20952
rect 43640 20890 43668 21354
rect 43824 20942 43852 21490
rect 43548 20862 43668 20890
rect 43812 20936 43864 20942
rect 43812 20878 43864 20884
rect 43444 20596 43496 20602
rect 43444 20538 43496 20544
rect 43352 20460 43404 20466
rect 43352 20402 43404 20408
rect 43444 19848 43496 19854
rect 43350 19816 43406 19825
rect 43444 19790 43496 19796
rect 43350 19751 43406 19760
rect 43364 19718 43392 19751
rect 43352 19712 43404 19718
rect 43272 19672 43352 19700
rect 43272 19514 43300 19672
rect 43352 19654 43404 19660
rect 43260 19508 43312 19514
rect 43260 19450 43312 19456
rect 43168 19440 43220 19446
rect 43168 19382 43220 19388
rect 43272 19378 43300 19450
rect 43456 19446 43484 19790
rect 43352 19440 43404 19446
rect 43352 19382 43404 19388
rect 43444 19440 43496 19446
rect 43444 19382 43496 19388
rect 43260 19372 43312 19378
rect 43260 19314 43312 19320
rect 43074 19272 43130 19281
rect 43074 19207 43130 19216
rect 43088 19174 43116 19207
rect 43076 19168 43128 19174
rect 43076 19110 43128 19116
rect 42984 18352 43036 18358
rect 42984 18294 43036 18300
rect 43272 18290 43300 19314
rect 42892 18284 42944 18290
rect 42892 18226 42944 18232
rect 43260 18284 43312 18290
rect 43260 18226 43312 18232
rect 43168 18080 43220 18086
rect 43168 18022 43220 18028
rect 42800 17808 42852 17814
rect 42800 17750 42852 17756
rect 42892 17808 42944 17814
rect 42892 17750 42944 17756
rect 42708 17672 42760 17678
rect 42708 17614 42760 17620
rect 42524 17604 42576 17610
rect 42524 17546 42576 17552
rect 42616 17604 42668 17610
rect 42616 17546 42668 17552
rect 42800 17536 42852 17542
rect 42720 17484 42800 17490
rect 42720 17478 42852 17484
rect 42720 17462 42840 17478
rect 42616 17196 42668 17202
rect 42616 17138 42668 17144
rect 42340 16516 42392 16522
rect 42340 16458 42392 16464
rect 42628 15638 42656 17138
rect 42616 15632 42668 15638
rect 42522 15600 42578 15609
rect 42616 15574 42668 15580
rect 42522 15535 42578 15544
rect 42536 15502 42564 15535
rect 42524 15496 42576 15502
rect 42524 15438 42576 15444
rect 42432 15156 42484 15162
rect 42432 15098 42484 15104
rect 42444 13326 42472 15098
rect 42720 15026 42748 17462
rect 42904 17202 42932 17750
rect 43180 17678 43208 18022
rect 43168 17672 43220 17678
rect 43168 17614 43220 17620
rect 43258 17640 43314 17649
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 42892 17196 42944 17202
rect 43076 17196 43128 17202
rect 42892 17138 42944 17144
rect 42996 17156 43076 17184
rect 42812 16454 42840 17138
rect 42800 16448 42852 16454
rect 42800 16390 42852 16396
rect 42800 15564 42852 15570
rect 42800 15506 42852 15512
rect 42812 15026 42840 15506
rect 42708 15020 42760 15026
rect 42708 14962 42760 14968
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42708 14884 42760 14890
rect 42708 14826 42760 14832
rect 42616 14408 42668 14414
rect 42616 14350 42668 14356
rect 42628 13938 42656 14350
rect 42616 13932 42668 13938
rect 42616 13874 42668 13880
rect 42720 13870 42748 14826
rect 42708 13864 42760 13870
rect 42708 13806 42760 13812
rect 42812 13394 42840 14962
rect 42892 14952 42944 14958
rect 42996 14940 43024 17156
rect 43076 17138 43128 17144
rect 43180 17082 43208 17614
rect 43258 17575 43314 17584
rect 43364 17592 43392 19382
rect 43444 18896 43496 18902
rect 43442 18864 43444 18873
rect 43548 18884 43576 20862
rect 44008 20806 44036 21966
rect 44100 21622 44128 22510
rect 44284 22030 44312 24210
rect 44548 23860 44600 23866
rect 44548 23802 44600 23808
rect 44560 23497 44588 23802
rect 44928 23662 44956 24772
rect 45008 24064 45060 24070
rect 45008 24006 45060 24012
rect 44916 23656 44968 23662
rect 44916 23598 44968 23604
rect 44928 23526 44956 23598
rect 44916 23520 44968 23526
rect 44546 23488 44602 23497
rect 44916 23462 44968 23468
rect 44546 23423 44602 23432
rect 45020 23322 45048 24006
rect 45008 23316 45060 23322
rect 45008 23258 45060 23264
rect 44640 23044 44692 23050
rect 44640 22986 44692 22992
rect 44652 22642 44680 22986
rect 45020 22642 45048 23258
rect 44640 22636 44692 22642
rect 44640 22578 44692 22584
rect 45008 22636 45060 22642
rect 45008 22578 45060 22584
rect 44272 22024 44324 22030
rect 44272 21966 44324 21972
rect 44456 21956 44508 21962
rect 44456 21898 44508 21904
rect 44088 21616 44140 21622
rect 44088 21558 44140 21564
rect 44468 21554 44496 21898
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 44456 21548 44508 21554
rect 44456 21490 44508 21496
rect 44088 21480 44140 21486
rect 44088 21422 44140 21428
rect 43720 20800 43772 20806
rect 43720 20742 43772 20748
rect 43996 20800 44048 20806
rect 43996 20742 44048 20748
rect 43732 20466 43760 20742
rect 43812 20596 43864 20602
rect 43812 20538 43864 20544
rect 43720 20460 43772 20466
rect 43720 20402 43772 20408
rect 43628 20324 43680 20330
rect 43628 20266 43680 20272
rect 43640 19417 43668 20266
rect 43626 19408 43682 19417
rect 43626 19343 43682 19352
rect 43496 18864 43576 18884
rect 43498 18856 43576 18864
rect 43732 18834 43760 20402
rect 43824 19689 43852 20538
rect 43810 19680 43866 19689
rect 43810 19615 43866 19624
rect 43442 18799 43498 18808
rect 43720 18828 43772 18834
rect 43720 18770 43772 18776
rect 43824 18766 43852 19615
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 43628 18760 43680 18766
rect 43628 18702 43680 18708
rect 43812 18760 43864 18766
rect 43812 18702 43864 18708
rect 43536 18624 43588 18630
rect 43536 18566 43588 18572
rect 43548 18426 43576 18566
rect 43536 18420 43588 18426
rect 43536 18362 43588 18368
rect 43444 18352 43496 18358
rect 43444 18294 43496 18300
rect 43456 17882 43484 18294
rect 43444 17876 43496 17882
rect 43444 17818 43496 17824
rect 43536 17604 43588 17610
rect 43272 17542 43300 17575
rect 43364 17564 43536 17592
rect 43536 17546 43588 17552
rect 43260 17536 43312 17542
rect 43548 17513 43576 17546
rect 43260 17478 43312 17484
rect 43534 17504 43590 17513
rect 43088 17054 43208 17082
rect 43088 16046 43116 17054
rect 43168 16992 43220 16998
rect 43168 16934 43220 16940
rect 43180 16658 43208 16934
rect 43168 16652 43220 16658
rect 43168 16594 43220 16600
rect 43076 16040 43128 16046
rect 43076 15982 43128 15988
rect 42944 14912 43024 14940
rect 42892 14894 42944 14900
rect 42996 14006 43024 14912
rect 42984 14000 43036 14006
rect 42984 13942 43036 13948
rect 43272 13462 43300 17478
rect 43534 17439 43590 17448
rect 43536 17196 43588 17202
rect 43536 17138 43588 17144
rect 43548 17066 43576 17138
rect 43536 17060 43588 17066
rect 43536 17002 43588 17008
rect 43640 16794 43668 18702
rect 43916 18612 43944 19314
rect 43732 18584 43944 18612
rect 43732 18193 43760 18584
rect 44008 18340 44036 20742
rect 44100 19922 44128 21422
rect 44192 20942 44220 21490
rect 44652 21350 44680 22578
rect 44824 21684 44876 21690
rect 44824 21626 44876 21632
rect 44640 21344 44692 21350
rect 44640 21286 44692 21292
rect 44180 20936 44232 20942
rect 44180 20878 44232 20884
rect 44456 20868 44508 20874
rect 44456 20810 44508 20816
rect 44180 20460 44232 20466
rect 44180 20402 44232 20408
rect 44088 19916 44140 19922
rect 44088 19858 44140 19864
rect 44100 19786 44128 19858
rect 44192 19854 44220 20402
rect 44272 20324 44324 20330
rect 44272 20266 44324 20272
rect 44284 19922 44312 20266
rect 44364 20256 44416 20262
rect 44362 20224 44364 20233
rect 44416 20224 44418 20233
rect 44362 20159 44418 20168
rect 44468 19922 44496 20810
rect 44548 20256 44600 20262
rect 44548 20198 44600 20204
rect 44272 19916 44324 19922
rect 44272 19858 44324 19864
rect 44456 19916 44508 19922
rect 44456 19858 44508 19864
rect 44180 19848 44232 19854
rect 44180 19790 44232 19796
rect 44088 19780 44140 19786
rect 44088 19722 44140 19728
rect 44088 19168 44140 19174
rect 44088 19110 44140 19116
rect 44100 18714 44128 19110
rect 44192 18970 44220 19790
rect 44272 19236 44324 19242
rect 44272 19178 44324 19184
rect 44180 18964 44232 18970
rect 44180 18906 44232 18912
rect 44284 18902 44312 19178
rect 44272 18896 44324 18902
rect 44272 18838 44324 18844
rect 44100 18686 44220 18714
rect 43916 18312 44036 18340
rect 43812 18284 43864 18290
rect 43812 18226 43864 18232
rect 43718 18184 43774 18193
rect 43718 18119 43774 18128
rect 43628 16788 43680 16794
rect 43628 16730 43680 16736
rect 43442 16688 43498 16697
rect 43732 16674 43760 18119
rect 43442 16623 43498 16632
rect 43548 16646 43760 16674
rect 43456 16590 43484 16623
rect 43352 16584 43404 16590
rect 43352 16526 43404 16532
rect 43444 16584 43496 16590
rect 43444 16526 43496 16532
rect 43364 16425 43392 16526
rect 43350 16416 43406 16425
rect 43350 16351 43406 16360
rect 43456 16114 43484 16526
rect 43444 16108 43496 16114
rect 43444 16050 43496 16056
rect 43352 14884 43404 14890
rect 43352 14826 43404 14832
rect 43364 14550 43392 14826
rect 43444 14612 43496 14618
rect 43444 14554 43496 14560
rect 43352 14544 43404 14550
rect 43352 14486 43404 14492
rect 43260 13456 43312 13462
rect 43260 13398 43312 13404
rect 42800 13388 42852 13394
rect 42800 13330 42852 13336
rect 43456 13326 43484 14554
rect 43548 14414 43576 16646
rect 43628 16584 43680 16590
rect 43720 16584 43772 16590
rect 43628 16526 43680 16532
rect 43718 16552 43720 16561
rect 43772 16552 43774 16561
rect 43640 16454 43668 16526
rect 43718 16487 43774 16496
rect 43628 16448 43680 16454
rect 43628 16390 43680 16396
rect 43640 16250 43668 16390
rect 43628 16244 43680 16250
rect 43628 16186 43680 16192
rect 43732 16114 43760 16487
rect 43824 16182 43852 18226
rect 43916 16998 43944 18312
rect 43994 17640 44050 17649
rect 44192 17610 44220 18686
rect 44284 18290 44312 18838
rect 44272 18284 44324 18290
rect 44272 18226 44324 18232
rect 43994 17575 43996 17584
rect 44048 17575 44050 17584
rect 44180 17604 44232 17610
rect 43996 17546 44048 17552
rect 44180 17546 44232 17552
rect 43996 17060 44048 17066
rect 43996 17002 44048 17008
rect 43904 16992 43956 16998
rect 43904 16934 43956 16940
rect 43904 16448 43956 16454
rect 43904 16390 43956 16396
rect 43812 16176 43864 16182
rect 43812 16118 43864 16124
rect 43720 16108 43772 16114
rect 43720 16050 43772 16056
rect 43628 15904 43680 15910
rect 43628 15846 43680 15852
rect 43536 14408 43588 14414
rect 43536 14350 43588 14356
rect 43548 13938 43576 14350
rect 43536 13932 43588 13938
rect 43536 13874 43588 13880
rect 43640 13802 43668 15846
rect 43916 15570 43944 16390
rect 43904 15564 43956 15570
rect 43904 15506 43956 15512
rect 43812 15496 43864 15502
rect 43812 15438 43864 15444
rect 43824 14822 43852 15438
rect 43812 14816 43864 14822
rect 43812 14758 43864 14764
rect 43824 14618 43852 14758
rect 43812 14612 43864 14618
rect 43812 14554 43864 14560
rect 43628 13796 43680 13802
rect 43628 13738 43680 13744
rect 44008 13326 44036 17002
rect 44088 16788 44140 16794
rect 44088 16730 44140 16736
rect 44100 16454 44128 16730
rect 44088 16448 44140 16454
rect 44088 16390 44140 16396
rect 44100 15162 44128 16390
rect 44284 16182 44312 18226
rect 44560 18222 44588 20198
rect 44836 20058 44864 21626
rect 45020 21554 45048 22578
rect 45100 22500 45152 22506
rect 45100 22442 45152 22448
rect 45008 21548 45060 21554
rect 45008 21490 45060 21496
rect 44824 20052 44876 20058
rect 44824 19994 44876 20000
rect 44916 19168 44968 19174
rect 44916 19110 44968 19116
rect 44928 18766 44956 19110
rect 44916 18760 44968 18766
rect 44916 18702 44968 18708
rect 44928 18290 44956 18702
rect 44916 18284 44968 18290
rect 44916 18226 44968 18232
rect 44548 18216 44600 18222
rect 44548 18158 44600 18164
rect 44928 17746 44956 18226
rect 44916 17740 44968 17746
rect 44916 17682 44968 17688
rect 44548 17536 44600 17542
rect 44548 17478 44600 17484
rect 44560 16590 44588 17478
rect 44928 17202 44956 17682
rect 45020 17270 45048 21490
rect 45112 21146 45140 22442
rect 45388 22030 45416 24840
rect 45468 24822 45520 24828
rect 45560 24812 45612 24818
rect 45560 24754 45612 24760
rect 45468 24676 45520 24682
rect 45468 24618 45520 24624
rect 45480 24342 45508 24618
rect 45468 24336 45520 24342
rect 45468 24278 45520 24284
rect 45572 23594 45600 24754
rect 46124 24206 46152 25230
rect 46112 24200 46164 24206
rect 46112 24142 46164 24148
rect 46020 24132 46072 24138
rect 46020 24074 46072 24080
rect 45560 23588 45612 23594
rect 45560 23530 45612 23536
rect 45572 23118 45600 23530
rect 45560 23112 45612 23118
rect 45560 23054 45612 23060
rect 45744 22636 45796 22642
rect 45744 22578 45796 22584
rect 45468 22568 45520 22574
rect 45468 22510 45520 22516
rect 45480 22030 45508 22510
rect 45756 22098 45784 22578
rect 45928 22160 45980 22166
rect 45928 22102 45980 22108
rect 45744 22092 45796 22098
rect 45744 22034 45796 22040
rect 45376 22024 45428 22030
rect 45376 21966 45428 21972
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45836 22024 45888 22030
rect 45836 21966 45888 21972
rect 45480 21622 45508 21966
rect 45848 21690 45876 21966
rect 45940 21690 45968 22102
rect 45836 21684 45888 21690
rect 45836 21626 45888 21632
rect 45928 21684 45980 21690
rect 45928 21626 45980 21632
rect 45468 21616 45520 21622
rect 45468 21558 45520 21564
rect 45284 21548 45336 21554
rect 45284 21490 45336 21496
rect 45100 21140 45152 21146
rect 45100 21082 45152 21088
rect 45192 20936 45244 20942
rect 45192 20878 45244 20884
rect 45100 20528 45152 20534
rect 45100 20470 45152 20476
rect 45112 19786 45140 20470
rect 45204 20466 45232 20878
rect 45192 20460 45244 20466
rect 45192 20402 45244 20408
rect 45190 19952 45246 19961
rect 45190 19887 45192 19896
rect 45244 19887 45246 19896
rect 45192 19858 45244 19864
rect 45100 19780 45152 19786
rect 45100 19722 45152 19728
rect 45112 17678 45140 19722
rect 45296 19174 45324 21490
rect 45652 20936 45704 20942
rect 45652 20878 45704 20884
rect 45664 20466 45692 20878
rect 45652 20460 45704 20466
rect 45652 20402 45704 20408
rect 45468 19848 45520 19854
rect 45468 19790 45520 19796
rect 45480 19718 45508 19790
rect 45468 19712 45520 19718
rect 45468 19654 45520 19660
rect 45560 19712 45612 19718
rect 45560 19654 45612 19660
rect 45572 19360 45600 19654
rect 45848 19378 45876 21626
rect 45940 20330 45968 21626
rect 45928 20324 45980 20330
rect 45928 20266 45980 20272
rect 45940 19854 45968 20266
rect 46032 20058 46060 24074
rect 46124 23730 46152 24142
rect 46112 23724 46164 23730
rect 46112 23666 46164 23672
rect 46112 23112 46164 23118
rect 46112 23054 46164 23060
rect 46020 20052 46072 20058
rect 46020 19994 46072 20000
rect 45928 19848 45980 19854
rect 45928 19790 45980 19796
rect 46032 19514 46060 19994
rect 46020 19508 46072 19514
rect 46020 19450 46072 19456
rect 45480 19332 45600 19360
rect 45836 19372 45888 19378
rect 45376 19304 45428 19310
rect 45376 19246 45428 19252
rect 45284 19168 45336 19174
rect 45284 19110 45336 19116
rect 45192 18216 45244 18222
rect 45192 18158 45244 18164
rect 45100 17672 45152 17678
rect 45100 17614 45152 17620
rect 45008 17264 45060 17270
rect 45008 17206 45060 17212
rect 44916 17196 44968 17202
rect 44916 17138 44968 17144
rect 44548 16584 44600 16590
rect 44548 16526 44600 16532
rect 44272 16176 44324 16182
rect 44272 16118 44324 16124
rect 44456 16040 44508 16046
rect 44456 15982 44508 15988
rect 44088 15156 44140 15162
rect 44088 15098 44140 15104
rect 44468 15026 44496 15982
rect 44456 15020 44508 15026
rect 44456 14962 44508 14968
rect 44456 14408 44508 14414
rect 44560 14396 44588 16526
rect 45112 15910 45140 17614
rect 45204 16114 45232 18158
rect 45192 16108 45244 16114
rect 45192 16050 45244 16056
rect 45100 15904 45152 15910
rect 45100 15846 45152 15852
rect 45112 15570 45140 15846
rect 45100 15564 45152 15570
rect 45100 15506 45152 15512
rect 45388 14618 45416 19246
rect 45480 17678 45508 19332
rect 45836 19314 45888 19320
rect 45848 18766 45876 19314
rect 46124 18970 46152 23054
rect 46112 18964 46164 18970
rect 46112 18906 46164 18912
rect 45836 18760 45888 18766
rect 45836 18702 45888 18708
rect 45744 18080 45796 18086
rect 45744 18022 45796 18028
rect 45468 17672 45520 17678
rect 45468 17614 45520 17620
rect 45480 16250 45508 17614
rect 45468 16244 45520 16250
rect 45468 16186 45520 16192
rect 45480 15502 45508 16186
rect 45652 15904 45704 15910
rect 45652 15846 45704 15852
rect 45664 15502 45692 15846
rect 45468 15496 45520 15502
rect 45468 15438 45520 15444
rect 45652 15496 45704 15502
rect 45652 15438 45704 15444
rect 45756 15484 45784 18022
rect 45848 17678 45876 18702
rect 46492 18154 46520 57394
rect 52288 57254 52316 57394
rect 52276 57248 52328 57254
rect 52276 57190 52328 57196
rect 57152 57248 57204 57254
rect 57152 57190 57204 57196
rect 58254 57216 58310 57225
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 52288 33454 52316 57190
rect 52276 33448 52328 33454
rect 52276 33390 52328 33396
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 57164 26858 57192 57190
rect 58254 57151 58310 57160
rect 58268 57050 58296 57151
rect 58256 57044 58308 57050
rect 58256 56986 58308 56992
rect 57612 56704 57664 56710
rect 57612 56646 57664 56652
rect 57244 51808 57296 51814
rect 57244 51750 57296 51756
rect 57256 37233 57284 51750
rect 57336 45824 57388 45830
rect 57336 45766 57388 45772
rect 57242 37224 57298 37233
rect 57242 37159 57298 37168
rect 57152 26852 57204 26858
rect 57152 26794 57204 26800
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 57348 24177 57376 45766
rect 57428 34536 57480 34542
rect 57428 34478 57480 34484
rect 57440 31210 57468 34478
rect 57428 31204 57480 31210
rect 57428 31146 57480 31152
rect 57624 26926 57652 56646
rect 58256 51808 58308 51814
rect 58254 51776 58256 51785
rect 58308 51776 58310 51785
rect 58254 51711 58310 51720
rect 58256 45824 58308 45830
rect 58256 45766 58308 45772
rect 58268 45665 58296 45766
rect 58254 45656 58310 45665
rect 58254 45591 58310 45600
rect 57704 40384 57756 40390
rect 57704 40326 57756 40332
rect 58256 40384 58308 40390
rect 58256 40326 58308 40332
rect 57612 26920 57664 26926
rect 57612 26862 57664 26868
rect 57334 24168 57390 24177
rect 57334 24103 57390 24112
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 46664 21344 46716 21350
rect 46664 21286 46716 21292
rect 46676 19922 46704 21286
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 46664 19916 46716 19922
rect 46664 19858 46716 19864
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 46480 18148 46532 18154
rect 46480 18090 46532 18096
rect 45836 17672 45888 17678
rect 45834 17640 45836 17649
rect 45888 17640 45890 17649
rect 45834 17575 45890 17584
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 57428 17128 57480 17134
rect 57426 17096 57428 17105
rect 57480 17096 57482 17105
rect 57426 17031 57482 17040
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 45836 15496 45888 15502
rect 45756 15456 45836 15484
rect 45376 14612 45428 14618
rect 45376 14554 45428 14560
rect 44508 14368 44588 14396
rect 44456 14350 44508 14356
rect 44272 14272 44324 14278
rect 44272 14214 44324 14220
rect 44180 14068 44232 14074
rect 44180 14010 44232 14016
rect 44088 13932 44140 13938
rect 44192 13920 44220 14010
rect 44284 13938 44312 14214
rect 44456 14000 44508 14006
rect 44362 13968 44418 13977
rect 44140 13892 44220 13920
rect 44088 13874 44140 13880
rect 44192 13326 44220 13892
rect 44272 13932 44324 13938
rect 44456 13942 44508 13948
rect 44362 13903 44364 13912
rect 44272 13874 44324 13880
rect 44416 13903 44418 13912
rect 44364 13874 44416 13880
rect 44468 13802 44496 13942
rect 44560 13920 44588 14368
rect 45480 13938 45508 15438
rect 44640 13932 44692 13938
rect 44560 13892 44640 13920
rect 44640 13874 44692 13880
rect 45468 13932 45520 13938
rect 45468 13874 45520 13880
rect 45664 13802 45692 15438
rect 45756 13870 45784 15456
rect 45836 15438 45888 15444
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 45744 13864 45796 13870
rect 45744 13806 45796 13812
rect 44456 13796 44508 13802
rect 44456 13738 44508 13744
rect 45652 13796 45704 13802
rect 45652 13738 45704 13744
rect 42432 13320 42484 13326
rect 42432 13262 42484 13268
rect 43444 13320 43496 13326
rect 43444 13262 43496 13268
rect 43996 13320 44048 13326
rect 43996 13262 44048 13268
rect 44180 13320 44232 13326
rect 44180 13262 44232 13268
rect 42248 13184 42300 13190
rect 42248 13126 42300 13132
rect 44468 12986 44496 13738
rect 45008 13728 45060 13734
rect 45008 13670 45060 13676
rect 44456 12980 44508 12986
rect 44456 12922 44508 12928
rect 41880 12912 41932 12918
rect 41880 12854 41932 12860
rect 41012 12804 41092 12832
rect 41236 12844 41288 12850
rect 40960 12786 41012 12792
rect 41236 12786 41288 12792
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 41892 12442 41920 12854
rect 45020 12714 45048 13670
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 45008 12708 45060 12714
rect 45008 12650 45060 12656
rect 40776 12436 40828 12442
rect 40776 12378 40828 12384
rect 41880 12436 41932 12442
rect 41880 12378 41932 12384
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 40592 11824 40644 11830
rect 40592 11766 40644 11772
rect 39212 11756 39264 11762
rect 39212 11698 39264 11704
rect 39304 11756 39356 11762
rect 39304 11698 39356 11704
rect 39120 11552 39172 11558
rect 39120 11494 39172 11500
rect 37740 11348 37792 11354
rect 37740 11290 37792 11296
rect 38200 11348 38252 11354
rect 38200 11290 38252 11296
rect 37200 11218 37412 11234
rect 37200 11212 37424 11218
rect 37200 11206 37372 11212
rect 37200 10062 37228 11206
rect 37372 11154 37424 11160
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37292 10810 37320 11086
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37292 9586 37320 10746
rect 37464 10124 37516 10130
rect 37464 10066 37516 10072
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37476 9450 37504 10066
rect 37752 9994 37780 11290
rect 39316 11286 39344 11698
rect 39764 11552 39816 11558
rect 39764 11494 39816 11500
rect 39304 11280 39356 11286
rect 39304 11222 39356 11228
rect 38568 11076 38620 11082
rect 38568 11018 38620 11024
rect 38292 10464 38344 10470
rect 38292 10406 38344 10412
rect 38304 10062 38332 10406
rect 38580 10062 38608 11018
rect 39776 10742 39804 11494
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 39764 10736 39816 10742
rect 39764 10678 39816 10684
rect 39120 10532 39172 10538
rect 39120 10474 39172 10480
rect 39132 10130 39160 10474
rect 39120 10124 39172 10130
rect 39120 10066 39172 10072
rect 38292 10056 38344 10062
rect 38568 10056 38620 10062
rect 38292 9998 38344 10004
rect 38488 10016 38568 10044
rect 37740 9988 37792 9994
rect 37740 9930 37792 9936
rect 38384 9988 38436 9994
rect 38384 9930 38436 9936
rect 37648 9920 37700 9926
rect 37648 9862 37700 9868
rect 37464 9444 37516 9450
rect 37464 9386 37516 9392
rect 37660 8974 37688 9862
rect 37752 9586 37780 9930
rect 38396 9722 38424 9930
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 38488 9518 38516 10016
rect 38568 9998 38620 10004
rect 39132 9518 39160 10066
rect 39776 10062 39804 10678
rect 39764 10056 39816 10062
rect 39764 9998 39816 10004
rect 57520 9920 57572 9926
rect 57520 9862 57572 9868
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 38476 9512 38528 9518
rect 38476 9454 38528 9460
rect 39120 9512 39172 9518
rect 39120 9454 39172 9460
rect 37648 8968 37700 8974
rect 37648 8910 37700 8916
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37660 8566 37688 8910
rect 37648 8560 37700 8566
rect 37648 8502 37700 8508
rect 37844 8362 37872 8910
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 37832 8356 37884 8362
rect 37832 8298 37884 8304
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37568 7886 37596 8230
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 57532 5914 57560 9862
rect 57716 8906 57744 40326
rect 58268 40225 58296 40326
rect 58254 40216 58310 40225
rect 58254 40151 58310 40160
rect 57888 34740 57940 34746
rect 57888 34682 57940 34688
rect 57900 34105 57928 34682
rect 57886 34096 57942 34105
rect 57886 34031 57942 34040
rect 57888 29028 57940 29034
rect 57888 28970 57940 28976
rect 57900 28665 57928 28970
rect 57886 28656 57942 28665
rect 57886 28591 57942 28600
rect 58164 26580 58216 26586
rect 58164 26522 58216 26528
rect 58176 11354 58204 26522
rect 58254 22536 58310 22545
rect 58254 22471 58256 22480
rect 58308 22471 58310 22480
rect 58256 22442 58308 22448
rect 58254 17096 58310 17105
rect 58254 17031 58256 17040
rect 58308 17031 58310 17040
rect 58256 17002 58308 17008
rect 58164 11348 58216 11354
rect 58164 11290 58216 11296
rect 58256 11076 58308 11082
rect 58256 11018 58308 11024
rect 58268 10985 58296 11018
rect 58254 10976 58310 10985
rect 58254 10911 58310 10920
rect 57704 8900 57756 8906
rect 57704 8842 57756 8848
rect 57520 5908 57572 5914
rect 57520 5850 57572 5856
rect 57532 5710 57560 5850
rect 57520 5704 57572 5710
rect 57520 5646 57572 5652
rect 58256 5568 58308 5574
rect 58254 5536 58256 5545
rect 58308 5536 58310 5545
rect 50294 5468 50602 5477
rect 58254 5471 58310 5480
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 44086 2680 44142 2689
rect 37096 2644 37148 2650
rect 44086 2615 44088 2624
rect 37096 2586 37148 2592
rect 44140 2615 44142 2624
rect 44180 2644 44232 2650
rect 44088 2586 44140 2592
rect 44180 2586 44232 2592
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 37108 2446 37136 2586
rect 44192 2530 44220 2586
rect 44008 2514 44220 2530
rect 43996 2508 44220 2514
rect 44048 2502 44220 2508
rect 43996 2450 44048 2456
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 22192 2372 22244 2378
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 18 200 74 800
rect 5170 200 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 2366
rect 22192 2314 22244 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 10980 800 11008 2246
rect 16132 800 16160 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21928 800 21956 2246
rect 27080 800 27108 2246
rect 32876 800 32904 2246
rect 38028 800 38056 2246
rect 43824 800 43852 2382
rect 48964 2304 49016 2310
rect 48964 2246 49016 2252
rect 55128 2304 55180 2310
rect 55128 2246 55180 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 48976 800 49004 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 54772 870 54892 898
rect 54772 800 54800 870
rect 5276 734 5488 762
rect 10966 200 11022 800
rect 16118 200 16174 800
rect 21914 200 21970 800
rect 27066 200 27122 800
rect 32862 200 32918 800
rect 38014 200 38070 800
rect 43810 200 43866 800
rect 48962 200 49018 800
rect 54758 200 54814 800
rect 54864 762 54892 870
rect 55140 762 55168 2246
rect 59924 800 59952 2246
rect 54864 734 55168 762
rect 59910 200 59966 800
<< via2 >>
rect 1674 57840 1730 57896
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 1674 51756 1676 51776
rect 1676 51756 1728 51776
rect 1728 51756 1730 51776
rect 1674 51720 1730 51756
rect 1674 46316 1676 46336
rect 1676 46316 1728 46336
rect 1728 46316 1730 46336
rect 1674 46280 1730 46316
rect 1674 40160 1730 40216
rect 1674 34720 1730 34776
rect 1674 28600 1730 28656
rect 1674 23160 1730 23216
rect 2134 27376 2190 27432
rect 1674 17060 1730 17096
rect 1674 17040 1676 17060
rect 1676 17040 1728 17060
rect 1728 17040 1730 17060
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 30562 56616 30618 56672
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 22098 46980 22154 47016
rect 22098 46960 22100 46980
rect 22100 46960 22152 46980
rect 22152 46960 22154 46980
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 20442 44412 20444 44432
rect 20444 44412 20496 44432
rect 20496 44412 20498 44432
rect 20442 44376 20498 44412
rect 17130 38664 17186 38720
rect 16486 37168 16542 37224
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1674 11620 1730 11656
rect 1674 11600 1676 11620
rect 1676 11600 1728 11620
rect 1728 11600 1730 11620
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1674 5516 1676 5536
rect 1676 5516 1728 5536
rect 1728 5516 1730 5536
rect 1674 5480 1730 5516
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 18602 38664 18658 38720
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19338 41248 19394 41304
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19982 41112 20038 41168
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20442 38664 20498 38720
rect 20626 43716 20682 43752
rect 20626 43696 20628 43716
rect 20628 43696 20680 43716
rect 20680 43696 20682 43716
rect 20718 42880 20774 42936
rect 20626 41248 20682 41304
rect 20902 45484 20958 45520
rect 20902 45464 20904 45484
rect 20904 45464 20956 45484
rect 20956 45464 20958 45484
rect 21454 44920 21510 44976
rect 21362 43832 21418 43888
rect 21178 38292 21180 38312
rect 21180 38292 21232 38312
rect 21232 38292 21234 38312
rect 21178 38256 21234 38292
rect 22742 45772 22744 45792
rect 22744 45772 22796 45792
rect 22796 45772 22798 45792
rect 22742 45736 22798 45772
rect 21822 43716 21878 43752
rect 21822 43696 21824 43716
rect 21824 43696 21876 43716
rect 21876 43696 21878 43716
rect 21362 39480 21418 39536
rect 22466 44820 22468 44840
rect 22468 44820 22520 44840
rect 22520 44820 22522 44840
rect 22466 44784 22522 44820
rect 21730 40468 21732 40488
rect 21732 40468 21784 40488
rect 21784 40468 21786 40488
rect 21730 40432 21786 40468
rect 21730 39344 21786 39400
rect 21454 37304 21510 37360
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 23294 45328 23350 45384
rect 22834 44396 22890 44432
rect 22834 44376 22836 44396
rect 22836 44376 22888 44396
rect 22888 44376 22890 44396
rect 22650 44240 22706 44296
rect 22190 41792 22246 41848
rect 22466 42608 22522 42664
rect 22282 40296 22338 40352
rect 22190 39888 22246 39944
rect 22006 39208 22062 39264
rect 22466 41384 22522 41440
rect 22466 41132 22522 41168
rect 22466 41112 22468 41132
rect 22468 41112 22520 41132
rect 22520 41112 22522 41132
rect 22374 39616 22430 39672
rect 22282 38664 22338 38720
rect 22742 42644 22744 42664
rect 22744 42644 22796 42664
rect 22796 42644 22798 42664
rect 22742 42608 22798 42644
rect 24030 44920 24086 44976
rect 22834 35808 22890 35864
rect 23294 40704 23350 40760
rect 23294 39752 23350 39808
rect 23386 39244 23388 39264
rect 23388 39244 23440 39264
rect 23440 39244 23442 39264
rect 23386 39208 23442 39244
rect 23478 39072 23534 39128
rect 24674 44920 24730 44976
rect 24398 44240 24454 44296
rect 23662 38936 23718 38992
rect 24398 42472 24454 42528
rect 24490 42336 24546 42392
rect 24398 40432 24454 40488
rect 23938 38664 23994 38720
rect 25318 44240 25374 44296
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 25502 45736 25558 45792
rect 25594 44920 25650 44976
rect 25410 43288 25466 43344
rect 25318 41556 25320 41576
rect 25320 41556 25372 41576
rect 25372 41556 25374 41576
rect 25318 41520 25374 41556
rect 24858 39616 24914 39672
rect 24214 35808 24270 35864
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 25134 39208 25190 39264
rect 25226 38256 25282 38312
rect 25042 37032 25098 37088
rect 25778 42472 25834 42528
rect 27526 44820 27528 44840
rect 27528 44820 27580 44840
rect 27580 44820 27582 44840
rect 27526 44784 27582 44820
rect 26514 44240 26570 44296
rect 25410 38664 25466 38720
rect 26054 40976 26110 41032
rect 26514 41248 26570 41304
rect 26514 40976 26570 41032
rect 26146 37984 26202 38040
rect 25686 35536 25742 35592
rect 25502 32408 25558 32464
rect 26514 39364 26570 39400
rect 26514 39344 26516 39364
rect 26516 39344 26568 39364
rect 26568 39344 26570 39364
rect 27158 42880 27214 42936
rect 26974 41384 27030 41440
rect 27158 41012 27160 41032
rect 27160 41012 27212 41032
rect 27212 41012 27214 41032
rect 27158 40976 27214 41012
rect 27526 41928 27582 41984
rect 27618 41792 27674 41848
rect 27342 41556 27344 41576
rect 27344 41556 27396 41576
rect 27396 41556 27398 41576
rect 27342 41520 27398 41556
rect 26974 39616 27030 39672
rect 26882 39480 26938 39536
rect 26514 39072 26570 39128
rect 26606 38800 26662 38856
rect 27618 41248 27674 41304
rect 27526 39888 27582 39944
rect 27526 39788 27528 39808
rect 27528 39788 27580 39808
rect 27580 39788 27582 39808
rect 27526 39752 27582 39788
rect 27802 39752 27858 39808
rect 27710 39616 27766 39672
rect 26330 34856 26386 34912
rect 27066 35536 27122 35592
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 17682 2508 17738 2544
rect 17682 2488 17684 2508
rect 17684 2488 17736 2508
rect 17736 2488 17738 2508
rect 24674 30776 24730 30832
rect 26238 30388 26294 30424
rect 26238 30368 26240 30388
rect 26240 30368 26292 30388
rect 26292 30368 26294 30388
rect 27618 39092 27674 39128
rect 27618 39072 27620 39092
rect 27620 39072 27672 39092
rect 27672 39072 27674 39092
rect 27802 38836 27804 38856
rect 27804 38836 27856 38856
rect 27856 38836 27858 38856
rect 27802 38800 27858 38836
rect 28078 41420 28080 41440
rect 28080 41420 28132 41440
rect 28132 41420 28134 41440
rect 28078 41384 28134 41420
rect 28262 41928 28318 41984
rect 28262 41248 28318 41304
rect 28170 40724 28226 40760
rect 28170 40704 28172 40724
rect 28172 40704 28224 40724
rect 28224 40704 28226 40724
rect 28170 40024 28226 40080
rect 28170 39208 28226 39264
rect 28078 38936 28134 38992
rect 27710 34448 27766 34504
rect 27526 34312 27582 34368
rect 28446 42336 28502 42392
rect 28630 45464 28686 45520
rect 28814 41384 28870 41440
rect 28722 41248 28778 41304
rect 28630 40160 28686 40216
rect 28446 38956 28502 38992
rect 28446 38936 28448 38956
rect 28448 38936 28500 38956
rect 28500 38936 28502 38956
rect 28446 38664 28502 38720
rect 29458 44104 29514 44160
rect 29274 41132 29330 41168
rect 29274 41112 29276 41132
rect 29276 41112 29328 41132
rect 29328 41112 29330 41132
rect 28998 40044 29054 40080
rect 28998 40024 29000 40044
rect 29000 40024 29052 40044
rect 29052 40024 29054 40044
rect 28722 38800 28778 38856
rect 29090 39072 29146 39128
rect 28538 37304 28594 37360
rect 29274 38800 29330 38856
rect 29182 35692 29238 35728
rect 29182 35672 29184 35692
rect 29184 35672 29236 35692
rect 29236 35672 29238 35692
rect 28814 34856 28870 34912
rect 29734 42880 29790 42936
rect 29550 39888 29606 39944
rect 29642 39344 29698 39400
rect 27250 32444 27252 32464
rect 27252 32444 27304 32464
rect 27304 32444 27306 32464
rect 27250 32408 27306 32444
rect 29458 35148 29514 35184
rect 29458 35128 29460 35148
rect 29460 35128 29512 35148
rect 29512 35128 29514 35148
rect 28538 31320 28594 31376
rect 28262 30368 28318 30424
rect 30470 39208 30526 39264
rect 30286 37340 30288 37360
rect 30288 37340 30340 37360
rect 30340 37340 30342 37360
rect 30286 37304 30342 37340
rect 30286 37068 30288 37088
rect 30288 37068 30340 37088
rect 30340 37068 30342 37088
rect 30286 37032 30342 37068
rect 30562 37032 30618 37088
rect 30930 37304 30986 37360
rect 31114 38700 31116 38720
rect 31116 38700 31168 38720
rect 31168 38700 31170 38720
rect 31114 38664 31170 38700
rect 30470 35672 30526 35728
rect 31758 39888 31814 39944
rect 31666 38800 31722 38856
rect 31574 38392 31630 38448
rect 31942 41384 31998 41440
rect 32770 44104 32826 44160
rect 32586 42472 32642 42528
rect 32034 38800 32090 38856
rect 31942 38392 31998 38448
rect 33690 43308 33746 43344
rect 33690 43288 33692 43308
rect 33692 43288 33744 43308
rect 33744 43288 33746 43308
rect 32770 41520 32826 41576
rect 33874 45772 33876 45792
rect 33876 45772 33928 45792
rect 33928 45772 33930 45792
rect 33874 45736 33930 45772
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 33874 44104 33930 44160
rect 32218 35672 32274 35728
rect 32310 29044 32312 29064
rect 32312 29044 32364 29064
rect 32364 29044 32366 29064
rect 32310 29008 32366 29044
rect 33690 41132 33746 41168
rect 33690 41112 33692 41132
rect 33692 41112 33744 41132
rect 33744 41112 33746 41132
rect 33966 41384 34022 41440
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34978 43852 35034 43888
rect 34978 43832 34980 43852
rect 34980 43832 35032 43852
rect 35032 43832 35034 43852
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34610 41520 34666 41576
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34058 35128 34114 35184
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 30470 26444 30526 26480
rect 30470 26424 30472 26444
rect 30472 26424 30524 26444
rect 30524 26424 30526 26444
rect 27434 24132 27490 24168
rect 27434 24112 27436 24132
rect 27436 24112 27488 24132
rect 27488 24112 27490 24132
rect 31390 25064 31446 25120
rect 28262 14864 28318 14920
rect 31666 20848 31722 20904
rect 31206 14068 31262 14104
rect 31206 14048 31208 14068
rect 31208 14048 31260 14068
rect 31260 14048 31262 14068
rect 33598 29008 33654 29064
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 32586 21664 32642 21720
rect 32126 17720 32182 17776
rect 32862 18808 32918 18864
rect 33506 21664 33562 21720
rect 33874 22072 33930 22128
rect 33230 17584 33286 17640
rect 33782 19896 33838 19952
rect 33874 19216 33930 19272
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34242 16496 34298 16552
rect 34426 14184 34482 14240
rect 34242 13776 34298 13832
rect 35346 21800 35402 21856
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 36818 26732 36820 26752
rect 36820 26732 36872 26752
rect 36872 26732 36874 26752
rect 36818 26696 36874 26732
rect 35714 21800 35770 21856
rect 35714 21292 35716 21312
rect 35716 21292 35768 21312
rect 35768 21292 35770 21312
rect 35714 21256 35770 21292
rect 35438 20712 35494 20768
rect 35622 20576 35678 20632
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35530 18708 35532 18728
rect 35532 18708 35584 18728
rect 35584 18708 35586 18728
rect 35530 18672 35586 18708
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35346 15136 35402 15192
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35622 15952 35678 16008
rect 35898 18808 35954 18864
rect 37002 23604 37004 23624
rect 37004 23604 37056 23624
rect 37056 23604 37058 23624
rect 37002 23568 37058 23604
rect 36634 19372 36690 19408
rect 36634 19352 36636 19372
rect 36636 19352 36688 19372
rect 36688 19352 36690 19372
rect 36726 17620 36728 17640
rect 36728 17620 36780 17640
rect 36780 17620 36782 17640
rect 36726 17584 36782 17620
rect 36634 16088 36690 16144
rect 36174 14456 36230 14512
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 36726 13388 36782 13424
rect 36726 13368 36728 13388
rect 36728 13368 36780 13388
rect 36780 13368 36782 13388
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 37002 17584 37058 17640
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37462 32000 37518 32056
rect 38382 27396 38438 27432
rect 38382 27376 38384 27396
rect 38384 27376 38436 27396
rect 38436 27376 38438 27396
rect 37830 24404 37886 24440
rect 37830 24384 37832 24404
rect 37832 24384 37884 24404
rect 37884 24384 37886 24404
rect 37738 21800 37794 21856
rect 37462 20868 37518 20904
rect 37462 20848 37464 20868
rect 37464 20848 37516 20868
rect 37516 20848 37518 20868
rect 37462 20576 37518 20632
rect 38014 21528 38070 21584
rect 37830 20168 37886 20224
rect 37830 19624 37886 19680
rect 37554 17584 37610 17640
rect 37922 18672 37978 18728
rect 38106 21256 38162 21312
rect 38014 18128 38070 18184
rect 37830 17312 37886 17368
rect 38106 17740 38162 17776
rect 38106 17720 38108 17740
rect 38108 17720 38160 17740
rect 38160 17720 38162 17740
rect 38106 17332 38162 17368
rect 38106 17312 38108 17332
rect 38108 17312 38160 17332
rect 38160 17312 38162 17332
rect 37922 13932 37978 13968
rect 37922 13912 37924 13932
rect 37924 13912 37976 13932
rect 37976 13912 37978 13932
rect 38474 21664 38530 21720
rect 38382 18284 38438 18320
rect 38382 18264 38384 18284
rect 38384 18264 38436 18284
rect 38436 18264 38438 18284
rect 38566 18808 38622 18864
rect 38658 17992 38714 18048
rect 38566 14884 38622 14920
rect 38566 14864 38568 14884
rect 38568 14864 38620 14884
rect 38620 14864 38622 14884
rect 38290 13912 38346 13968
rect 38566 14456 38622 14512
rect 38658 14320 38714 14376
rect 38474 13776 38530 13832
rect 39394 23704 39450 23760
rect 39118 22752 39174 22808
rect 39302 22652 39304 22672
rect 39304 22652 39356 22672
rect 39356 22652 39358 22672
rect 39302 22616 39358 22652
rect 40130 22752 40186 22808
rect 40038 22480 40094 22536
rect 40038 22072 40094 22128
rect 40222 21972 40224 21992
rect 40224 21972 40276 21992
rect 40276 21972 40278 21992
rect 40222 21936 40278 21972
rect 39670 21528 39726 21584
rect 39578 19080 39634 19136
rect 39210 18264 39266 18320
rect 38934 13776 38990 13832
rect 39486 17448 39542 17504
rect 39302 16108 39358 16144
rect 39302 16088 39304 16108
rect 39304 16088 39356 16108
rect 39356 16088 39358 16108
rect 39762 15000 39818 15056
rect 39486 14864 39542 14920
rect 39210 14456 39266 14512
rect 41602 24384 41658 24440
rect 41878 23704 41934 23760
rect 41234 23432 41290 23488
rect 41234 23060 41236 23080
rect 41236 23060 41288 23080
rect 41288 23060 41290 23080
rect 41234 23024 41290 23060
rect 40866 22652 40868 22672
rect 40868 22652 40920 22672
rect 40920 22652 40922 22672
rect 40866 22616 40922 22652
rect 40498 20748 40500 20768
rect 40500 20748 40552 20768
rect 40552 20748 40554 20768
rect 40498 20712 40554 20748
rect 40866 20576 40922 20632
rect 40130 18264 40186 18320
rect 40222 15700 40278 15736
rect 40222 15680 40224 15700
rect 40224 15680 40276 15700
rect 40276 15680 40278 15700
rect 39854 14320 39910 14376
rect 39670 13912 39726 13968
rect 40498 16360 40554 16416
rect 40222 15136 40278 15192
rect 40222 15000 40278 15056
rect 40406 13912 40462 13968
rect 40314 13504 40370 13560
rect 40866 19760 40922 19816
rect 41326 21548 41382 21584
rect 41326 21528 41328 21548
rect 41328 21528 41380 21548
rect 41380 21528 41382 21548
rect 41602 21800 41658 21856
rect 41234 17992 41290 18048
rect 41970 20052 42026 20088
rect 41970 20032 41972 20052
rect 41972 20032 42024 20052
rect 42024 20032 42026 20052
rect 41694 18808 41750 18864
rect 41418 17584 41474 17640
rect 40682 15136 40738 15192
rect 40682 14048 40738 14104
rect 41234 16532 41236 16552
rect 41236 16532 41288 16552
rect 41288 16532 41290 16552
rect 41234 16496 41290 16532
rect 40866 14864 40922 14920
rect 40682 13776 40738 13832
rect 41602 15020 41658 15056
rect 41602 15000 41604 15020
rect 41604 15000 41656 15020
rect 41656 15000 41658 15020
rect 41878 15952 41934 16008
rect 41786 14864 41842 14920
rect 40958 14184 41014 14240
rect 42614 22752 42670 22808
rect 43074 22208 43130 22264
rect 43166 21936 43222 21992
rect 42246 19080 42302 19136
rect 41970 13932 42026 13968
rect 41970 13912 41972 13932
rect 41972 13912 42024 13932
rect 42024 13912 42026 13932
rect 42062 13504 42118 13560
rect 43902 23024 43958 23080
rect 43350 19760 43406 19816
rect 43074 19216 43130 19272
rect 42522 15544 42578 15600
rect 43258 17584 43314 17640
rect 44546 23432 44602 23488
rect 43626 19352 43682 19408
rect 43442 18844 43444 18864
rect 43444 18844 43496 18864
rect 43496 18844 43498 18864
rect 43442 18808 43498 18844
rect 43810 19624 43866 19680
rect 43534 17448 43590 17504
rect 44362 20204 44364 20224
rect 44364 20204 44416 20224
rect 44416 20204 44418 20224
rect 44362 20168 44418 20204
rect 43718 18128 43774 18184
rect 43442 16632 43498 16688
rect 43350 16360 43406 16416
rect 43718 16532 43720 16552
rect 43720 16532 43772 16552
rect 43772 16532 43774 16552
rect 43718 16496 43774 16532
rect 43994 17604 44050 17640
rect 43994 17584 43996 17604
rect 43996 17584 44048 17604
rect 44048 17584 44050 17604
rect 45190 19916 45246 19952
rect 45190 19896 45192 19916
rect 45192 19896 45244 19916
rect 45244 19896 45246 19916
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 58254 57160 58310 57216
rect 57242 37168 57298 37224
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 58254 51756 58256 51776
rect 58256 51756 58308 51776
rect 58308 51756 58310 51776
rect 58254 51720 58310 51756
rect 58254 45600 58310 45656
rect 57334 24112 57390 24168
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 45834 17620 45836 17640
rect 45836 17620 45888 17640
rect 45888 17620 45890 17640
rect 45834 17584 45890 17620
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 57426 17076 57428 17096
rect 57428 17076 57480 17096
rect 57480 17076 57482 17096
rect 57426 17040 57482 17076
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 44362 13932 44418 13968
rect 44362 13912 44364 13932
rect 44364 13912 44416 13932
rect 44416 13912 44418 13932
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 58254 40160 58310 40216
rect 57886 34040 57942 34096
rect 57886 28600 57942 28656
rect 58254 22500 58310 22536
rect 58254 22480 58256 22500
rect 58256 22480 58308 22500
rect 58308 22480 58310 22500
rect 58254 17060 58310 17096
rect 58254 17040 58256 17060
rect 58256 17040 58308 17060
rect 58308 17040 58310 17060
rect 58254 10920 58310 10976
rect 58254 5516 58256 5536
rect 58256 5516 58308 5536
rect 58308 5516 58310 5536
rect 58254 5480 58310 5516
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 44086 2644 44142 2680
rect 44086 2624 44088 2644
rect 44088 2624 44140 2644
rect 44140 2624 44142 2644
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 200 57898 800 57928
rect 1669 57898 1735 57901
rect 200 57896 1735 57898
rect 200 57840 1674 57896
rect 1730 57840 1735 57896
rect 200 57838 1735 57840
rect 200 57808 800 57838
rect 1669 57835 1735 57838
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 58249 57218 58315 57221
rect 59200 57218 59800 57248
rect 58249 57216 59800 57218
rect 58249 57160 58254 57216
rect 58310 57160 59800 57216
rect 58249 57158 59800 57160
rect 58249 57155 58315 57158
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 59800 57158
rect 34930 57087 35246 57088
rect 30557 56676 30623 56677
rect 30557 56672 30604 56676
rect 30668 56674 30674 56676
rect 30557 56616 30562 56672
rect 30557 56612 30604 56616
rect 30668 56614 30714 56674
rect 30668 56612 30674 56614
rect 30557 56611 30623 56612
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 200 51778 800 51808
rect 1669 51778 1735 51781
rect 200 51776 1735 51778
rect 200 51720 1674 51776
rect 1730 51720 1735 51776
rect 200 51718 1735 51720
rect 200 51688 800 51718
rect 1669 51715 1735 51718
rect 58249 51778 58315 51781
rect 59200 51778 59800 51808
rect 58249 51776 59800 51778
rect 58249 51720 58254 51776
rect 58310 51720 59800 51776
rect 58249 51718 59800 51720
rect 58249 51715 58315 51718
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 59800 51718
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 22093 47020 22159 47021
rect 22093 47016 22140 47020
rect 22204 47018 22210 47020
rect 22093 46960 22098 47016
rect 22093 46956 22140 46960
rect 22204 46958 22250 47018
rect 22204 46956 22210 46958
rect 22093 46955 22159 46956
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 200 46338 800 46368
rect 1669 46338 1735 46341
rect 200 46336 1735 46338
rect 200 46280 1674 46336
rect 1730 46280 1735 46336
rect 200 46278 1735 46280
rect 200 46248 800 46278
rect 1669 46275 1735 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 22737 45794 22803 45797
rect 25497 45794 25563 45797
rect 22737 45792 25563 45794
rect 22737 45736 22742 45792
rect 22798 45736 25502 45792
rect 25558 45736 25563 45792
rect 22737 45734 25563 45736
rect 22737 45731 22803 45734
rect 25497 45731 25563 45734
rect 33726 45732 33732 45796
rect 33796 45794 33802 45796
rect 33869 45794 33935 45797
rect 33796 45792 33935 45794
rect 33796 45736 33874 45792
rect 33930 45736 33935 45792
rect 33796 45734 33935 45736
rect 33796 45732 33802 45734
rect 33869 45731 33935 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58249 45658 58315 45661
rect 59200 45658 59800 45688
rect 58249 45656 59800 45658
rect 58249 45600 58254 45656
rect 58310 45600 59800 45656
rect 58249 45598 59800 45600
rect 58249 45595 58315 45598
rect 59200 45568 59800 45598
rect 20897 45522 20963 45525
rect 28625 45522 28691 45525
rect 20897 45520 28691 45522
rect 20897 45464 20902 45520
rect 20958 45464 28630 45520
rect 28686 45464 28691 45520
rect 20897 45462 28691 45464
rect 20897 45459 20963 45462
rect 28625 45459 28691 45462
rect 23289 45386 23355 45389
rect 23422 45386 23428 45388
rect 23289 45384 23428 45386
rect 23289 45328 23294 45384
rect 23350 45328 23428 45384
rect 23289 45326 23428 45328
rect 23289 45323 23355 45326
rect 23422 45324 23428 45326
rect 23492 45324 23498 45388
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 21449 44978 21515 44981
rect 24025 44978 24091 44981
rect 21449 44976 24091 44978
rect 21449 44920 21454 44976
rect 21510 44920 24030 44976
rect 24086 44920 24091 44976
rect 21449 44918 24091 44920
rect 21449 44915 21515 44918
rect 24025 44915 24091 44918
rect 24669 44978 24735 44981
rect 25589 44978 25655 44981
rect 33726 44978 33732 44980
rect 24669 44976 33732 44978
rect 24669 44920 24674 44976
rect 24730 44920 25594 44976
rect 25650 44920 33732 44976
rect 24669 44918 33732 44920
rect 24669 44915 24735 44918
rect 25589 44915 25655 44918
rect 33726 44916 33732 44918
rect 33796 44916 33802 44980
rect 22461 44842 22527 44845
rect 27521 44842 27587 44845
rect 22461 44840 27587 44842
rect 22461 44784 22466 44840
rect 22522 44784 27526 44840
rect 27582 44784 27587 44840
rect 22461 44782 27587 44784
rect 22461 44779 22527 44782
rect 27521 44779 27587 44782
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 20437 44434 20503 44437
rect 22829 44434 22895 44437
rect 20437 44432 22895 44434
rect 20437 44376 20442 44432
rect 20498 44376 22834 44432
rect 22890 44376 22895 44432
rect 20437 44374 22895 44376
rect 20437 44371 20503 44374
rect 22829 44371 22895 44374
rect 22645 44298 22711 44301
rect 24393 44300 24459 44301
rect 22870 44298 22876 44300
rect 22645 44296 22876 44298
rect 22645 44240 22650 44296
rect 22706 44240 22876 44296
rect 22645 44238 22876 44240
rect 22645 44235 22711 44238
rect 22870 44236 22876 44238
rect 22940 44236 22946 44300
rect 24342 44298 24348 44300
rect 24302 44238 24348 44298
rect 24412 44296 24459 44300
rect 24454 44240 24459 44296
rect 24342 44236 24348 44238
rect 24412 44236 24459 44240
rect 24894 44236 24900 44300
rect 24964 44298 24970 44300
rect 25313 44298 25379 44301
rect 24964 44296 25379 44298
rect 24964 44240 25318 44296
rect 25374 44240 25379 44296
rect 24964 44238 25379 44240
rect 24964 44236 24970 44238
rect 24393 44235 24459 44236
rect 25313 44235 25379 44238
rect 26509 44300 26575 44301
rect 26509 44296 26556 44300
rect 26620 44298 26626 44300
rect 26509 44240 26514 44296
rect 26509 44236 26556 44240
rect 26620 44238 26666 44298
rect 26620 44236 26626 44238
rect 26509 44235 26575 44236
rect 29453 44162 29519 44165
rect 32765 44162 32831 44165
rect 33869 44162 33935 44165
rect 29453 44160 33935 44162
rect 29453 44104 29458 44160
rect 29514 44104 32770 44160
rect 32826 44104 33874 44160
rect 33930 44104 33935 44160
rect 29453 44102 33935 44104
rect 29453 44099 29519 44102
rect 32765 44099 32831 44102
rect 33869 44099 33935 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 21357 43890 21423 43893
rect 34973 43890 35039 43893
rect 21357 43888 35039 43890
rect 21357 43832 21362 43888
rect 21418 43832 34978 43888
rect 35034 43832 35039 43888
rect 21357 43830 35039 43832
rect 21357 43827 21423 43830
rect 34973 43827 35039 43830
rect 20621 43754 20687 43757
rect 21817 43754 21883 43757
rect 20621 43752 21883 43754
rect 20621 43696 20626 43752
rect 20682 43696 21822 43752
rect 21878 43696 21883 43752
rect 20621 43694 21883 43696
rect 20621 43691 20687 43694
rect 21817 43691 21883 43694
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 25405 43346 25471 43349
rect 33685 43346 33751 43349
rect 25405 43344 33751 43346
rect 25405 43288 25410 43344
rect 25466 43288 33690 43344
rect 33746 43288 33751 43344
rect 25405 43286 33751 43288
rect 25405 43283 25471 43286
rect 33685 43283 33751 43286
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 20713 42938 20779 42941
rect 27153 42938 27219 42941
rect 20713 42936 27219 42938
rect 20713 42880 20718 42936
rect 20774 42880 27158 42936
rect 27214 42880 27219 42936
rect 20713 42878 27219 42880
rect 20713 42875 20779 42878
rect 27153 42875 27219 42878
rect 28942 42876 28948 42940
rect 29012 42938 29018 42940
rect 29729 42938 29795 42941
rect 29012 42936 29795 42938
rect 29012 42880 29734 42936
rect 29790 42880 29795 42936
rect 29012 42878 29795 42880
rect 29012 42876 29018 42878
rect 29729 42875 29795 42878
rect 22461 42666 22527 42669
rect 22737 42666 22803 42669
rect 22461 42664 22803 42666
rect 22461 42608 22466 42664
rect 22522 42608 22742 42664
rect 22798 42608 22803 42664
rect 22461 42606 22803 42608
rect 22461 42603 22527 42606
rect 22737 42603 22803 42606
rect 24393 42530 24459 42533
rect 25773 42530 25839 42533
rect 32581 42530 32647 42533
rect 24393 42528 32647 42530
rect 24393 42472 24398 42528
rect 24454 42472 25778 42528
rect 25834 42472 32586 42528
rect 32642 42472 32647 42528
rect 24393 42470 32647 42472
rect 24393 42467 24459 42470
rect 25773 42467 25839 42470
rect 32581 42467 32647 42470
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 24485 42394 24551 42397
rect 28441 42394 28507 42397
rect 24485 42392 28507 42394
rect 24485 42336 24490 42392
rect 24546 42336 28446 42392
rect 28502 42336 28507 42392
rect 24485 42334 28507 42336
rect 24485 42331 24551 42334
rect 28441 42331 28507 42334
rect 27521 41988 27587 41989
rect 27470 41986 27476 41988
rect 27430 41926 27476 41986
rect 27540 41984 27587 41988
rect 27582 41928 27587 41984
rect 27470 41924 27476 41926
rect 27540 41924 27587 41928
rect 27521 41923 27587 41924
rect 28257 41986 28323 41989
rect 28390 41986 28396 41988
rect 28257 41984 28396 41986
rect 28257 41928 28262 41984
rect 28318 41928 28396 41984
rect 28257 41926 28396 41928
rect 28257 41923 28323 41926
rect 28390 41924 28396 41926
rect 28460 41924 28466 41988
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 22185 41850 22251 41853
rect 27613 41850 27679 41853
rect 22185 41848 27679 41850
rect 22185 41792 22190 41848
rect 22246 41792 27618 41848
rect 27674 41792 27679 41848
rect 22185 41790 27679 41792
rect 22185 41787 22251 41790
rect 27613 41787 27679 41790
rect 25313 41578 25379 41581
rect 27337 41578 27403 41581
rect 25313 41576 27403 41578
rect 25313 41520 25318 41576
rect 25374 41520 27342 41576
rect 27398 41520 27403 41576
rect 25313 41518 27403 41520
rect 25313 41515 25379 41518
rect 27337 41515 27403 41518
rect 32765 41578 32831 41581
rect 34605 41578 34671 41581
rect 32765 41576 34671 41578
rect 32765 41520 32770 41576
rect 32826 41520 34610 41576
rect 34666 41520 34671 41576
rect 32765 41518 34671 41520
rect 32765 41515 32831 41518
rect 34605 41515 34671 41518
rect 22461 41442 22527 41445
rect 26969 41442 27035 41445
rect 22461 41440 27035 41442
rect 22461 41384 22466 41440
rect 22522 41384 26974 41440
rect 27030 41384 27035 41440
rect 22461 41382 27035 41384
rect 22461 41379 22527 41382
rect 26969 41379 27035 41382
rect 28073 41442 28139 41445
rect 28809 41442 28875 41445
rect 28073 41440 28875 41442
rect 28073 41384 28078 41440
rect 28134 41384 28814 41440
rect 28870 41384 28875 41440
rect 28073 41382 28875 41384
rect 28073 41379 28139 41382
rect 28809 41379 28875 41382
rect 31937 41442 32003 41445
rect 33961 41442 34027 41445
rect 31937 41440 34027 41442
rect 31937 41384 31942 41440
rect 31998 41384 33966 41440
rect 34022 41384 34027 41440
rect 31937 41382 34027 41384
rect 31937 41379 32003 41382
rect 33961 41379 34027 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 19333 41306 19399 41309
rect 20621 41306 20687 41309
rect 26509 41306 26575 41309
rect 27613 41306 27679 41309
rect 19333 41304 19442 41306
rect 19333 41248 19338 41304
rect 19394 41248 19442 41304
rect 19333 41243 19442 41248
rect 20621 41304 27679 41306
rect 20621 41248 20626 41304
rect 20682 41248 26514 41304
rect 26570 41248 27618 41304
rect 27674 41248 27679 41304
rect 20621 41246 27679 41248
rect 20621 41243 20687 41246
rect 26509 41243 26575 41246
rect 27613 41243 27679 41246
rect 28257 41306 28323 41309
rect 28717 41306 28783 41309
rect 28257 41304 28783 41306
rect 28257 41248 28262 41304
rect 28318 41248 28722 41304
rect 28778 41248 28783 41304
rect 28257 41246 28783 41248
rect 28257 41243 28323 41246
rect 28717 41243 28783 41246
rect 19382 41170 19442 41243
rect 19977 41170 20043 41173
rect 19382 41168 20043 41170
rect 19382 41112 19982 41168
rect 20038 41112 20043 41168
rect 19382 41110 20043 41112
rect 19977 41107 20043 41110
rect 22461 41170 22527 41173
rect 29126 41170 29132 41172
rect 22461 41168 29132 41170
rect 22461 41112 22466 41168
rect 22522 41112 29132 41168
rect 22461 41110 29132 41112
rect 22461 41107 22527 41110
rect 29126 41108 29132 41110
rect 29196 41170 29202 41172
rect 29269 41170 29335 41173
rect 33685 41172 33751 41173
rect 33685 41170 33732 41172
rect 29196 41168 29335 41170
rect 29196 41112 29274 41168
rect 29330 41112 29335 41168
rect 29196 41110 29335 41112
rect 33640 41168 33732 41170
rect 33640 41112 33690 41168
rect 33640 41110 33732 41112
rect 29196 41108 29202 41110
rect 29269 41107 29335 41110
rect 33685 41108 33732 41110
rect 33796 41108 33802 41172
rect 33685 41107 33751 41108
rect 26049 41034 26115 41037
rect 26509 41034 26575 41037
rect 26049 41032 26575 41034
rect 26049 40976 26054 41032
rect 26110 40976 26514 41032
rect 26570 40976 26575 41032
rect 26049 40974 26575 40976
rect 26049 40971 26115 40974
rect 26509 40971 26575 40974
rect 27153 41034 27219 41037
rect 27286 41034 27292 41036
rect 27153 41032 27292 41034
rect 27153 40976 27158 41032
rect 27214 40976 27292 41032
rect 27153 40974 27292 40976
rect 27153 40971 27219 40974
rect 27286 40972 27292 40974
rect 27356 40972 27362 41036
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 23289 40762 23355 40765
rect 28165 40762 28231 40765
rect 23289 40760 28231 40762
rect 23289 40704 23294 40760
rect 23350 40704 28170 40760
rect 28226 40704 28231 40760
rect 23289 40702 28231 40704
rect 23289 40699 23355 40702
rect 28165 40699 28231 40702
rect 21725 40490 21791 40493
rect 24393 40490 24459 40493
rect 21725 40488 24459 40490
rect 21725 40432 21730 40488
rect 21786 40432 24398 40488
rect 24454 40432 24459 40488
rect 21725 40430 24459 40432
rect 21725 40427 21791 40430
rect 24393 40427 24459 40430
rect 22277 40354 22343 40357
rect 27838 40354 27844 40356
rect 22277 40352 27844 40354
rect 22277 40296 22282 40352
rect 22338 40296 27844 40352
rect 22277 40294 27844 40296
rect 22277 40291 22343 40294
rect 27838 40292 27844 40294
rect 27908 40292 27914 40356
rect 19570 40288 19886 40289
rect 200 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 1669 40218 1735 40221
rect 200 40216 1735 40218
rect 200 40160 1674 40216
rect 1730 40160 1735 40216
rect 200 40158 1735 40160
rect 200 40128 800 40158
rect 1669 40155 1735 40158
rect 27654 40156 27660 40220
rect 27724 40218 27730 40220
rect 28625 40218 28691 40221
rect 27724 40216 28691 40218
rect 27724 40160 28630 40216
rect 28686 40160 28691 40216
rect 27724 40158 28691 40160
rect 27724 40156 27730 40158
rect 28625 40155 28691 40158
rect 58249 40218 58315 40221
rect 59200 40218 59800 40248
rect 58249 40216 59800 40218
rect 58249 40160 58254 40216
rect 58310 40160 59800 40216
rect 58249 40158 59800 40160
rect 58249 40155 58315 40158
rect 59200 40128 59800 40158
rect 28165 40082 28231 40085
rect 28993 40082 29059 40085
rect 28165 40080 29059 40082
rect 28165 40024 28170 40080
rect 28226 40024 28998 40080
rect 29054 40024 29059 40080
rect 28165 40022 29059 40024
rect 28165 40019 28231 40022
rect 28993 40019 29059 40022
rect 22185 39948 22251 39949
rect 22134 39946 22140 39948
rect 22094 39886 22140 39946
rect 22204 39944 22251 39948
rect 22246 39888 22251 39944
rect 22134 39884 22140 39886
rect 22204 39884 22251 39888
rect 22185 39883 22251 39884
rect 27521 39946 27587 39949
rect 29545 39946 29611 39949
rect 31753 39946 31819 39949
rect 27521 39944 27860 39946
rect 27521 39888 27526 39944
rect 27582 39888 27860 39944
rect 27521 39886 27860 39888
rect 27521 39883 27587 39886
rect 27800 39813 27860 39886
rect 29545 39944 31819 39946
rect 29545 39888 29550 39944
rect 29606 39888 31758 39944
rect 31814 39888 31819 39944
rect 29545 39886 31819 39888
rect 29545 39883 29611 39886
rect 31753 39883 31819 39886
rect 23289 39810 23355 39813
rect 24894 39810 24900 39812
rect 23289 39808 24900 39810
rect 23289 39752 23294 39808
rect 23350 39752 24900 39808
rect 23289 39750 24900 39752
rect 23289 39747 23355 39750
rect 24894 39748 24900 39750
rect 24964 39748 24970 39812
rect 26550 39748 26556 39812
rect 26620 39810 26626 39812
rect 27521 39810 27587 39813
rect 26620 39808 27587 39810
rect 26620 39752 27526 39808
rect 27582 39752 27587 39808
rect 26620 39750 27587 39752
rect 26620 39748 26626 39750
rect 27521 39747 27587 39750
rect 27797 39808 27863 39813
rect 27797 39752 27802 39808
rect 27858 39752 27863 39808
rect 27797 39747 27863 39752
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 22369 39674 22435 39677
rect 24853 39674 24919 39677
rect 22369 39672 24919 39674
rect 22369 39616 22374 39672
rect 22430 39616 24858 39672
rect 24914 39616 24919 39672
rect 22369 39614 24919 39616
rect 22369 39611 22435 39614
rect 24853 39611 24919 39614
rect 26969 39674 27035 39677
rect 27705 39674 27771 39677
rect 26969 39672 27771 39674
rect 26969 39616 26974 39672
rect 27030 39616 27710 39672
rect 27766 39616 27771 39672
rect 26969 39614 27771 39616
rect 26969 39611 27035 39614
rect 27705 39611 27771 39614
rect 21357 39538 21423 39541
rect 26877 39538 26943 39541
rect 21357 39536 26943 39538
rect 21357 39480 21362 39536
rect 21418 39480 26882 39536
rect 26938 39480 26943 39536
rect 21357 39478 26943 39480
rect 21357 39475 21423 39478
rect 26877 39475 26943 39478
rect 21725 39402 21791 39405
rect 26509 39402 26575 39405
rect 29637 39402 29703 39405
rect 21725 39400 29703 39402
rect 21725 39344 21730 39400
rect 21786 39344 26514 39400
rect 26570 39344 29642 39400
rect 29698 39344 29703 39400
rect 21725 39342 29703 39344
rect 21725 39339 21791 39342
rect 26509 39339 26575 39342
rect 29637 39339 29703 39342
rect 22001 39266 22067 39269
rect 23381 39266 23447 39269
rect 22001 39264 23447 39266
rect 22001 39208 22006 39264
rect 22062 39208 23386 39264
rect 23442 39208 23447 39264
rect 22001 39206 23447 39208
rect 22001 39203 22067 39206
rect 23381 39203 23447 39206
rect 25129 39266 25195 39269
rect 28165 39266 28231 39269
rect 30465 39266 30531 39269
rect 25129 39264 28231 39266
rect 25129 39208 25134 39264
rect 25190 39208 28170 39264
rect 28226 39208 28231 39264
rect 25129 39206 28231 39208
rect 25129 39203 25195 39206
rect 28165 39203 28231 39206
rect 30422 39264 30531 39266
rect 30422 39208 30470 39264
rect 30526 39208 30531 39264
rect 30422 39203 30531 39208
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 23473 39130 23539 39133
rect 26509 39130 26575 39133
rect 27613 39130 27679 39133
rect 23473 39128 27679 39130
rect 23473 39072 23478 39128
rect 23534 39072 26514 39128
rect 26570 39072 27618 39128
rect 27674 39072 27679 39128
rect 23473 39070 27679 39072
rect 23473 39067 23539 39070
rect 26509 39067 26575 39070
rect 27613 39067 27679 39070
rect 29085 39130 29151 39133
rect 30422 39130 30482 39203
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 29085 39128 30482 39130
rect 29085 39072 29090 39128
rect 29146 39072 30482 39128
rect 29085 39070 30482 39072
rect 29085 39067 29151 39070
rect 23422 38932 23428 38996
rect 23492 38994 23498 38996
rect 23657 38994 23723 38997
rect 28073 38994 28139 38997
rect 28441 38994 28507 38997
rect 23492 38992 28507 38994
rect 23492 38936 23662 38992
rect 23718 38936 28078 38992
rect 28134 38936 28446 38992
rect 28502 38936 28507 38992
rect 23492 38934 28507 38936
rect 23492 38932 23498 38934
rect 23657 38931 23723 38934
rect 28073 38931 28139 38934
rect 28441 38931 28507 38934
rect 26601 38860 26667 38861
rect 26550 38796 26556 38860
rect 26620 38858 26667 38860
rect 27797 38860 27863 38861
rect 27797 38858 27844 38860
rect 26620 38856 26712 38858
rect 26662 38800 26712 38856
rect 26620 38798 26712 38800
rect 27752 38856 27844 38858
rect 27908 38858 27914 38860
rect 28717 38858 28783 38861
rect 29269 38858 29335 38861
rect 27908 38856 29335 38858
rect 27752 38800 27802 38856
rect 27908 38800 28722 38856
rect 28778 38800 29274 38856
rect 29330 38800 29335 38856
rect 27752 38798 27844 38800
rect 26620 38796 26667 38798
rect 26601 38795 26667 38796
rect 27797 38796 27844 38798
rect 27908 38798 29335 38800
rect 27908 38796 27914 38798
rect 27797 38795 27863 38796
rect 28717 38795 28783 38798
rect 29269 38795 29335 38798
rect 31661 38858 31727 38861
rect 32029 38858 32095 38861
rect 31661 38856 32095 38858
rect 31661 38800 31666 38856
rect 31722 38800 32034 38856
rect 32090 38800 32095 38856
rect 31661 38798 32095 38800
rect 31661 38795 31727 38798
rect 32029 38795 32095 38798
rect 17125 38722 17191 38725
rect 18597 38722 18663 38725
rect 17125 38720 18663 38722
rect 17125 38664 17130 38720
rect 17186 38664 18602 38720
rect 18658 38664 18663 38720
rect 17125 38662 18663 38664
rect 17125 38659 17191 38662
rect 18597 38659 18663 38662
rect 20437 38722 20503 38725
rect 22277 38722 22343 38725
rect 20437 38720 22343 38722
rect 20437 38664 20442 38720
rect 20498 38664 22282 38720
rect 22338 38664 22343 38720
rect 20437 38662 22343 38664
rect 20437 38659 20503 38662
rect 22277 38659 22343 38662
rect 23933 38722 23999 38725
rect 24710 38722 24716 38724
rect 23933 38720 24716 38722
rect 23933 38664 23938 38720
rect 23994 38664 24716 38720
rect 23933 38662 24716 38664
rect 23933 38659 23999 38662
rect 24710 38660 24716 38662
rect 24780 38660 24786 38724
rect 25405 38722 25471 38725
rect 27286 38722 27292 38724
rect 25405 38720 27292 38722
rect 25405 38664 25410 38720
rect 25466 38664 27292 38720
rect 25405 38662 27292 38664
rect 25405 38659 25471 38662
rect 27286 38660 27292 38662
rect 27356 38722 27362 38724
rect 28441 38722 28507 38725
rect 27356 38720 28507 38722
rect 27356 38664 28446 38720
rect 28502 38664 28507 38720
rect 27356 38662 28507 38664
rect 27356 38660 27362 38662
rect 28441 38659 28507 38662
rect 31109 38724 31175 38725
rect 31109 38720 31156 38724
rect 31220 38722 31226 38724
rect 31109 38664 31114 38720
rect 31109 38660 31156 38664
rect 31220 38662 31266 38722
rect 31220 38660 31226 38662
rect 31109 38659 31175 38660
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 31569 38450 31635 38453
rect 31937 38450 32003 38453
rect 31569 38448 32003 38450
rect 31569 38392 31574 38448
rect 31630 38392 31942 38448
rect 31998 38392 32003 38448
rect 31569 38390 32003 38392
rect 31569 38387 31635 38390
rect 31937 38387 32003 38390
rect 21173 38314 21239 38317
rect 25221 38314 25287 38317
rect 21173 38312 25287 38314
rect 21173 38256 21178 38312
rect 21234 38256 25226 38312
rect 25282 38256 25287 38312
rect 21173 38254 25287 38256
rect 21173 38251 21239 38254
rect 25221 38251 25287 38254
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 26141 38042 26207 38045
rect 28942 38042 28948 38044
rect 26141 38040 28948 38042
rect 26141 37984 26146 38040
rect 26202 37984 28948 38040
rect 26141 37982 28948 37984
rect 26141 37979 26207 37982
rect 28942 37980 28948 37982
rect 29012 37980 29018 38044
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 21449 37362 21515 37365
rect 28533 37362 28599 37365
rect 21449 37360 28599 37362
rect 21449 37304 21454 37360
rect 21510 37304 28538 37360
rect 28594 37304 28599 37360
rect 21449 37302 28599 37304
rect 21449 37299 21515 37302
rect 28533 37299 28599 37302
rect 30281 37362 30347 37365
rect 30925 37362 30991 37365
rect 30281 37360 30991 37362
rect 30281 37304 30286 37360
rect 30342 37304 30930 37360
rect 30986 37304 30991 37360
rect 30281 37302 30991 37304
rect 30281 37299 30347 37302
rect 30925 37299 30991 37302
rect 16481 37226 16547 37229
rect 57237 37226 57303 37229
rect 16481 37224 57303 37226
rect 16481 37168 16486 37224
rect 16542 37168 57242 37224
rect 57298 37168 57303 37224
rect 16481 37166 57303 37168
rect 16481 37163 16547 37166
rect 57237 37163 57303 37166
rect 25037 37090 25103 37093
rect 27654 37090 27660 37092
rect 25037 37088 27660 37090
rect 25037 37032 25042 37088
rect 25098 37032 27660 37088
rect 25037 37030 27660 37032
rect 25037 37027 25103 37030
rect 27654 37028 27660 37030
rect 27724 37028 27730 37092
rect 30281 37090 30347 37093
rect 30557 37090 30623 37093
rect 30281 37088 30623 37090
rect 30281 37032 30286 37088
rect 30342 37032 30562 37088
rect 30618 37032 30623 37088
rect 30281 37030 30623 37032
rect 30281 37027 30347 37030
rect 30557 37027 30623 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 22829 35868 22895 35869
rect 22829 35866 22876 35868
rect 22784 35864 22876 35866
rect 22784 35808 22834 35864
rect 22784 35806 22876 35808
rect 22829 35804 22876 35806
rect 22940 35804 22946 35868
rect 24209 35866 24275 35869
rect 24342 35866 24348 35868
rect 24209 35864 24348 35866
rect 24209 35808 24214 35864
rect 24270 35808 24348 35864
rect 24209 35806 24348 35808
rect 22829 35803 22895 35804
rect 24209 35803 24275 35806
rect 24342 35804 24348 35806
rect 24412 35804 24418 35868
rect 29177 35732 29243 35733
rect 29126 35668 29132 35732
rect 29196 35730 29243 35732
rect 30465 35730 30531 35733
rect 32213 35730 32279 35733
rect 29196 35728 29288 35730
rect 29238 35672 29288 35728
rect 29196 35670 29288 35672
rect 30465 35728 32279 35730
rect 30465 35672 30470 35728
rect 30526 35672 32218 35728
rect 32274 35672 32279 35728
rect 30465 35670 32279 35672
rect 29196 35668 29243 35670
rect 29177 35667 29243 35668
rect 30465 35667 30531 35670
rect 32213 35667 32279 35670
rect 25681 35594 25747 35597
rect 27061 35594 27127 35597
rect 25681 35592 27127 35594
rect 25681 35536 25686 35592
rect 25742 35536 27066 35592
rect 27122 35536 27127 35592
rect 25681 35534 27127 35536
rect 25681 35531 25747 35534
rect 27061 35531 27127 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 29453 35186 29519 35189
rect 34053 35186 34119 35189
rect 29453 35184 34119 35186
rect 29453 35128 29458 35184
rect 29514 35128 34058 35184
rect 34114 35128 34119 35184
rect 29453 35126 34119 35128
rect 29453 35123 29519 35126
rect 34053 35123 34119 35126
rect 26325 34914 26391 34917
rect 28809 34914 28875 34917
rect 26325 34912 28875 34914
rect 26325 34856 26330 34912
rect 26386 34856 28814 34912
rect 28870 34856 28875 34912
rect 26325 34854 28875 34856
rect 26325 34851 26391 34854
rect 28809 34851 28875 34854
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 1669 34778 1735 34781
rect 200 34776 1735 34778
rect 200 34720 1674 34776
rect 1730 34720 1735 34776
rect 200 34718 1735 34720
rect 200 34688 800 34718
rect 1669 34715 1735 34718
rect 27470 34444 27476 34508
rect 27540 34506 27546 34508
rect 27705 34506 27771 34509
rect 27540 34504 27771 34506
rect 27540 34448 27710 34504
rect 27766 34448 27771 34504
rect 27540 34446 27771 34448
rect 27540 34444 27546 34446
rect 27705 34443 27771 34446
rect 27521 34370 27587 34373
rect 28390 34370 28396 34372
rect 27521 34368 28396 34370
rect 27521 34312 27526 34368
rect 27582 34312 28396 34368
rect 27521 34310 28396 34312
rect 27521 34307 27587 34310
rect 28390 34308 28396 34310
rect 28460 34308 28466 34372
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 57881 34098 57947 34101
rect 59200 34098 59800 34128
rect 57881 34096 59800 34098
rect 57881 34040 57886 34096
rect 57942 34040 59800 34096
rect 57881 34038 59800 34040
rect 57881 34035 57947 34038
rect 59200 34008 59800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 25497 32466 25563 32469
rect 27245 32466 27311 32469
rect 25497 32464 27311 32466
rect 25497 32408 25502 32464
rect 25558 32408 27250 32464
rect 27306 32408 27311 32464
rect 25497 32406 27311 32408
rect 25497 32403 25563 32406
rect 27245 32403 27311 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 37457 32058 37523 32061
rect 37590 32058 37596 32060
rect 37457 32056 37596 32058
rect 37457 32000 37462 32056
rect 37518 32000 37596 32056
rect 37457 31998 37596 32000
rect 37457 31995 37523 31998
rect 37590 31996 37596 31998
rect 37660 31996 37666 32060
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 28533 31378 28599 31381
rect 31150 31378 31156 31380
rect 28533 31376 31156 31378
rect 28533 31320 28538 31376
rect 28594 31320 31156 31376
rect 28533 31318 31156 31320
rect 28533 31315 28599 31318
rect 31150 31316 31156 31318
rect 31220 31316 31226 31380
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 24669 30836 24735 30837
rect 24669 30834 24716 30836
rect 24624 30832 24716 30834
rect 24624 30776 24674 30832
rect 24624 30774 24716 30776
rect 24669 30772 24716 30774
rect 24780 30772 24786 30836
rect 24669 30771 24735 30772
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 26233 30426 26299 30429
rect 28257 30426 28323 30429
rect 26233 30424 28323 30426
rect 26233 30368 26238 30424
rect 26294 30368 28262 30424
rect 28318 30368 28323 30424
rect 26233 30366 28323 30368
rect 26233 30363 26299 30366
rect 28257 30363 28323 30366
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 32305 29066 32371 29069
rect 33593 29066 33659 29069
rect 32305 29064 33659 29066
rect 32305 29008 32310 29064
rect 32366 29008 33598 29064
rect 33654 29008 33659 29064
rect 32305 29006 33659 29008
rect 32305 29003 32371 29006
rect 33593 29003 33659 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1669 28658 1735 28661
rect 200 28656 1735 28658
rect 200 28600 1674 28656
rect 1730 28600 1735 28656
rect 200 28598 1735 28600
rect 200 28568 800 28598
rect 1669 28595 1735 28598
rect 57881 28658 57947 28661
rect 59200 28658 59800 28688
rect 57881 28656 59800 28658
rect 57881 28600 57886 28656
rect 57942 28600 59800 28656
rect 57881 28598 59800 28600
rect 57881 28595 57947 28598
rect 59200 28568 59800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 2129 27434 2195 27437
rect 38377 27434 38443 27437
rect 2129 27432 38443 27434
rect 2129 27376 2134 27432
rect 2190 27376 38382 27432
rect 38438 27376 38443 27432
rect 2129 27374 38443 27376
rect 2129 27371 2195 27374
rect 38377 27371 38443 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 36813 26756 36879 26757
rect 36813 26754 36860 26756
rect 36768 26752 36860 26754
rect 36768 26696 36818 26752
rect 36768 26694 36860 26696
rect 36813 26692 36860 26694
rect 36924 26692 36930 26756
rect 36813 26691 36879 26692
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 30465 26482 30531 26485
rect 30598 26482 30604 26484
rect 30465 26480 30604 26482
rect 30465 26424 30470 26480
rect 30526 26424 30604 26480
rect 30465 26422 30604 26424
rect 30465 26419 30531 26422
rect 30598 26420 30604 26422
rect 30668 26420 30674 26484
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 31385 25122 31451 25125
rect 31518 25122 31524 25124
rect 31385 25120 31524 25122
rect 31385 25064 31390 25120
rect 31446 25064 31524 25120
rect 31385 25062 31524 25064
rect 31385 25059 31451 25062
rect 31518 25060 31524 25062
rect 31588 25060 31594 25124
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 37825 24442 37891 24445
rect 41597 24442 41663 24445
rect 37825 24440 41663 24442
rect 37825 24384 37830 24440
rect 37886 24384 41602 24440
rect 41658 24384 41663 24440
rect 37825 24382 41663 24384
rect 37825 24379 37891 24382
rect 41597 24379 41663 24382
rect 27429 24170 27495 24173
rect 57329 24170 57395 24173
rect 27429 24168 57395 24170
rect 27429 24112 27434 24168
rect 27490 24112 57334 24168
rect 57390 24112 57395 24168
rect 27429 24110 57395 24112
rect 27429 24107 27495 24110
rect 57329 24107 57395 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 39389 23762 39455 23765
rect 41873 23762 41939 23765
rect 38610 23760 41939 23762
rect 38610 23704 39394 23760
rect 39450 23704 41878 23760
rect 41934 23704 41939 23760
rect 38610 23702 41939 23704
rect 31518 23564 31524 23628
rect 31588 23626 31594 23628
rect 36997 23626 37063 23629
rect 38610 23626 38670 23702
rect 39389 23699 39455 23702
rect 41873 23699 41939 23702
rect 31588 23624 38670 23626
rect 31588 23568 37002 23624
rect 37058 23568 38670 23624
rect 31588 23566 38670 23568
rect 31588 23564 31594 23566
rect 36997 23563 37063 23566
rect 39982 23428 39988 23492
rect 40052 23490 40058 23492
rect 41229 23490 41295 23493
rect 40052 23488 41295 23490
rect 40052 23432 41234 23488
rect 41290 23432 41295 23488
rect 40052 23430 41295 23432
rect 40052 23428 40058 23430
rect 41229 23427 41295 23430
rect 44541 23492 44607 23493
rect 44541 23488 44588 23492
rect 44652 23490 44658 23492
rect 44541 23432 44546 23488
rect 44541 23428 44588 23432
rect 44652 23430 44698 23490
rect 44652 23428 44658 23430
rect 44541 23427 44607 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 41229 23082 41295 23085
rect 43897 23082 43963 23085
rect 41229 23080 43963 23082
rect 41229 23024 41234 23080
rect 41290 23024 43902 23080
rect 43958 23024 43963 23080
rect 41229 23022 43963 23024
rect 41229 23019 41295 23022
rect 43897 23019 43963 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 39113 22810 39179 22813
rect 40125 22810 40191 22813
rect 42609 22810 42675 22813
rect 39113 22808 42675 22810
rect 39113 22752 39118 22808
rect 39174 22752 40130 22808
rect 40186 22752 42614 22808
rect 42670 22752 42675 22808
rect 39113 22750 42675 22752
rect 39113 22747 39179 22750
rect 40125 22747 40191 22750
rect 42609 22747 42675 22750
rect 39297 22674 39363 22677
rect 40861 22674 40927 22677
rect 39297 22672 40927 22674
rect 39297 22616 39302 22672
rect 39358 22616 40866 22672
rect 40922 22616 40927 22672
rect 39297 22614 40927 22616
rect 39297 22611 39363 22614
rect 40861 22611 40927 22614
rect 40033 22538 40099 22541
rect 40166 22538 40172 22540
rect 40033 22536 40172 22538
rect 40033 22480 40038 22536
rect 40094 22480 40172 22536
rect 40033 22478 40172 22480
rect 40033 22475 40099 22478
rect 40166 22476 40172 22478
rect 40236 22476 40242 22540
rect 58249 22538 58315 22541
rect 59200 22538 59800 22568
rect 58249 22536 59800 22538
rect 58249 22480 58254 22536
rect 58310 22480 59800 22536
rect 58249 22478 59800 22480
rect 58249 22475 58315 22478
rect 59200 22448 59800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 43069 22268 43135 22269
rect 43069 22264 43116 22268
rect 43180 22266 43186 22268
rect 43069 22208 43074 22264
rect 43069 22204 43116 22208
rect 43180 22206 43226 22266
rect 43180 22204 43186 22206
rect 43069 22203 43135 22204
rect 33869 22130 33935 22133
rect 40033 22130 40099 22133
rect 33869 22128 40099 22130
rect 33869 22072 33874 22128
rect 33930 22072 40038 22128
rect 40094 22072 40099 22128
rect 33869 22070 40099 22072
rect 33869 22067 33935 22070
rect 40033 22067 40099 22070
rect 40217 21994 40283 21997
rect 43161 21994 43227 21997
rect 40217 21992 43227 21994
rect 40217 21936 40222 21992
rect 40278 21936 43166 21992
rect 43222 21936 43227 21992
rect 40217 21934 43227 21936
rect 40217 21931 40283 21934
rect 43161 21931 43227 21934
rect 35341 21858 35407 21861
rect 35709 21858 35775 21861
rect 35341 21856 35775 21858
rect 35341 21800 35346 21856
rect 35402 21800 35714 21856
rect 35770 21800 35775 21856
rect 35341 21798 35775 21800
rect 35341 21795 35407 21798
rect 35709 21795 35775 21798
rect 37733 21858 37799 21861
rect 41597 21858 41663 21861
rect 37733 21856 41663 21858
rect 37733 21800 37738 21856
rect 37794 21800 41602 21856
rect 41658 21800 41663 21856
rect 37733 21798 41663 21800
rect 37733 21795 37799 21798
rect 41597 21795 41663 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 32581 21722 32647 21725
rect 33501 21722 33567 21725
rect 38469 21722 38535 21725
rect 32581 21720 38535 21722
rect 32581 21664 32586 21720
rect 32642 21664 33506 21720
rect 33562 21664 38474 21720
rect 38530 21664 38535 21720
rect 32581 21662 38535 21664
rect 32581 21659 32647 21662
rect 33501 21659 33567 21662
rect 38469 21659 38535 21662
rect 38009 21586 38075 21589
rect 39665 21586 39731 21589
rect 41321 21586 41387 21589
rect 38009 21584 41387 21586
rect 38009 21528 38014 21584
rect 38070 21528 39670 21584
rect 39726 21528 41326 21584
rect 41382 21528 41387 21584
rect 38009 21526 41387 21528
rect 38009 21523 38075 21526
rect 39665 21523 39731 21526
rect 41321 21523 41387 21526
rect 35709 21314 35775 21317
rect 38101 21314 38167 21317
rect 35709 21312 38167 21314
rect 35709 21256 35714 21312
rect 35770 21256 38106 21312
rect 38162 21256 38167 21312
rect 35709 21254 38167 21256
rect 35709 21251 35775 21254
rect 38101 21251 38167 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 31661 20906 31727 20909
rect 37457 20906 37523 20909
rect 31661 20904 37523 20906
rect 31661 20848 31666 20904
rect 31722 20848 37462 20904
rect 37518 20848 37523 20904
rect 31661 20846 37523 20848
rect 31661 20843 31727 20846
rect 37457 20843 37523 20846
rect 35433 20770 35499 20773
rect 40493 20772 40559 20773
rect 40493 20770 40540 20772
rect 35433 20768 40540 20770
rect 35433 20712 35438 20768
rect 35494 20712 40498 20768
rect 35433 20710 40540 20712
rect 35433 20707 35499 20710
rect 40493 20708 40540 20710
rect 40604 20708 40610 20772
rect 40493 20707 40559 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 35617 20634 35683 20637
rect 37457 20634 37523 20637
rect 40861 20634 40927 20637
rect 35617 20632 35818 20634
rect 35617 20576 35622 20632
rect 35678 20576 35818 20632
rect 35617 20574 35818 20576
rect 35617 20571 35683 20574
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 35758 20090 35818 20574
rect 37457 20632 40927 20634
rect 37457 20576 37462 20632
rect 37518 20576 40866 20632
rect 40922 20576 40927 20632
rect 37457 20574 40927 20576
rect 37457 20571 37523 20574
rect 40861 20571 40927 20574
rect 37825 20226 37891 20229
rect 44214 20226 44220 20228
rect 37825 20224 44220 20226
rect 37825 20168 37830 20224
rect 37886 20168 44220 20224
rect 37825 20166 44220 20168
rect 37825 20163 37891 20166
rect 44214 20164 44220 20166
rect 44284 20226 44290 20228
rect 44357 20226 44423 20229
rect 44284 20224 44423 20226
rect 44284 20168 44362 20224
rect 44418 20168 44423 20224
rect 44284 20166 44423 20168
rect 44284 20164 44290 20166
rect 44357 20163 44423 20166
rect 41965 20090 42031 20093
rect 35758 20088 42031 20090
rect 35758 20032 41970 20088
rect 42026 20032 42031 20088
rect 35758 20030 42031 20032
rect 41965 20027 42031 20030
rect 33777 19954 33843 19957
rect 44398 19954 44404 19956
rect 33777 19952 44404 19954
rect 33777 19896 33782 19952
rect 33838 19896 44404 19952
rect 33777 19894 44404 19896
rect 33777 19891 33843 19894
rect 44398 19892 44404 19894
rect 44468 19954 44474 19956
rect 45185 19954 45251 19957
rect 44468 19952 45251 19954
rect 44468 19896 45190 19952
rect 45246 19896 45251 19952
rect 44468 19894 45251 19896
rect 44468 19892 44474 19894
rect 45185 19891 45251 19894
rect 40861 19818 40927 19821
rect 43345 19818 43411 19821
rect 40861 19816 43411 19818
rect 40861 19760 40866 19816
rect 40922 19760 43350 19816
rect 43406 19760 43411 19816
rect 40861 19758 43411 19760
rect 40861 19755 40927 19758
rect 43345 19755 43411 19758
rect 37825 19682 37891 19685
rect 43805 19682 43871 19685
rect 37825 19680 43871 19682
rect 37825 19624 37830 19680
rect 37886 19624 43810 19680
rect 43866 19624 43871 19680
rect 37825 19622 43871 19624
rect 37825 19619 37891 19622
rect 43805 19619 43871 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 36629 19412 36695 19413
rect 43621 19412 43687 19413
rect 36629 19410 36676 19412
rect 36548 19408 36676 19410
rect 36740 19410 36746 19412
rect 39982 19410 39988 19412
rect 36548 19352 36634 19408
rect 36548 19350 36676 19352
rect 36629 19348 36676 19350
rect 36740 19350 39988 19410
rect 36740 19348 36746 19350
rect 39982 19348 39988 19350
rect 40052 19348 40058 19412
rect 43621 19408 43668 19412
rect 43732 19410 43738 19412
rect 43621 19352 43626 19408
rect 43621 19348 43668 19352
rect 43732 19350 43778 19410
rect 43732 19348 43738 19350
rect 36629 19347 36695 19348
rect 43621 19347 43687 19348
rect 33869 19274 33935 19277
rect 43069 19274 43135 19277
rect 33869 19272 43135 19274
rect 33869 19216 33874 19272
rect 33930 19216 43074 19272
rect 43130 19216 43135 19272
rect 33869 19214 43135 19216
rect 33869 19211 33935 19214
rect 43069 19211 43135 19214
rect 39573 19138 39639 19141
rect 42241 19138 42307 19141
rect 39573 19136 42307 19138
rect 39573 19080 39578 19136
rect 39634 19080 42246 19136
rect 42302 19080 42307 19136
rect 39573 19078 42307 19080
rect 39573 19075 39639 19078
rect 42241 19075 42307 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 32857 18866 32923 18869
rect 35893 18866 35959 18869
rect 32857 18864 35959 18866
rect 32857 18808 32862 18864
rect 32918 18808 35898 18864
rect 35954 18808 35959 18864
rect 32857 18806 35959 18808
rect 32857 18803 32923 18806
rect 35893 18803 35959 18806
rect 38561 18866 38627 18869
rect 41689 18866 41755 18869
rect 38561 18864 41755 18866
rect 38561 18808 38566 18864
rect 38622 18808 41694 18864
rect 41750 18808 41755 18864
rect 38561 18806 41755 18808
rect 38561 18803 38627 18806
rect 41689 18803 41755 18806
rect 43294 18804 43300 18868
rect 43364 18866 43370 18868
rect 43437 18866 43503 18869
rect 43364 18864 43503 18866
rect 43364 18808 43442 18864
rect 43498 18808 43503 18864
rect 43364 18806 43503 18808
rect 43364 18804 43370 18806
rect 43437 18803 43503 18806
rect 35525 18730 35591 18733
rect 37917 18730 37983 18733
rect 35525 18728 37983 18730
rect 35525 18672 35530 18728
rect 35586 18672 37922 18728
rect 37978 18672 37983 18728
rect 35525 18670 37983 18672
rect 35525 18667 35591 18670
rect 37917 18667 37983 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 38377 18322 38443 18325
rect 39205 18322 39271 18325
rect 40125 18322 40191 18325
rect 38377 18320 40191 18322
rect 38377 18264 38382 18320
rect 38438 18264 39210 18320
rect 39266 18264 40130 18320
rect 40186 18264 40191 18320
rect 38377 18262 40191 18264
rect 38377 18259 38443 18262
rect 39205 18259 39271 18262
rect 40125 18259 40191 18262
rect 38009 18186 38075 18189
rect 43713 18186 43779 18189
rect 38009 18184 43779 18186
rect 38009 18128 38014 18184
rect 38070 18128 43718 18184
rect 43774 18128 43779 18184
rect 38009 18126 43779 18128
rect 38009 18123 38075 18126
rect 43713 18123 43779 18126
rect 38653 18050 38719 18053
rect 41229 18050 41295 18053
rect 38653 18048 41295 18050
rect 38653 17992 38658 18048
rect 38714 17992 41234 18048
rect 41290 17992 41295 18048
rect 38653 17990 41295 17992
rect 38653 17987 38719 17990
rect 41229 17987 41295 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 32121 17778 32187 17781
rect 38101 17778 38167 17781
rect 32121 17776 38167 17778
rect 32121 17720 32126 17776
rect 32182 17720 38106 17776
rect 38162 17720 38167 17776
rect 32121 17718 38167 17720
rect 32121 17715 32187 17718
rect 38101 17715 38167 17718
rect 33225 17642 33291 17645
rect 36721 17642 36787 17645
rect 36997 17642 37063 17645
rect 33225 17640 37063 17642
rect 33225 17584 33230 17640
rect 33286 17584 36726 17640
rect 36782 17584 37002 17640
rect 37058 17584 37063 17640
rect 33225 17582 37063 17584
rect 33225 17579 33291 17582
rect 36721 17579 36787 17582
rect 36997 17579 37063 17582
rect 37549 17642 37615 17645
rect 41413 17642 41479 17645
rect 43253 17642 43319 17645
rect 37549 17640 43319 17642
rect 37549 17584 37554 17640
rect 37610 17584 41418 17640
rect 41474 17584 43258 17640
rect 43314 17584 43319 17640
rect 37549 17582 43319 17584
rect 37549 17579 37615 17582
rect 41413 17579 41479 17582
rect 43253 17579 43319 17582
rect 43989 17642 44055 17645
rect 45829 17642 45895 17645
rect 43989 17640 45895 17642
rect 43989 17584 43994 17640
rect 44050 17584 45834 17640
rect 45890 17584 45895 17640
rect 43989 17582 45895 17584
rect 43989 17579 44055 17582
rect 45829 17579 45895 17582
rect 39481 17506 39547 17509
rect 43529 17506 43595 17509
rect 39481 17504 43595 17506
rect 39481 17448 39486 17504
rect 39542 17448 43534 17504
rect 43590 17448 43595 17504
rect 39481 17446 43595 17448
rect 39481 17443 39547 17446
rect 43529 17443 43595 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 37825 17370 37891 17373
rect 38101 17370 38167 17373
rect 37825 17368 38167 17370
rect 37825 17312 37830 17368
rect 37886 17312 38106 17368
rect 38162 17312 38167 17368
rect 37825 17310 38167 17312
rect 37825 17307 37891 17310
rect 38101 17307 38167 17310
rect 200 17098 800 17128
rect 1669 17098 1735 17101
rect 200 17096 1735 17098
rect 200 17040 1674 17096
rect 1730 17040 1735 17096
rect 200 17038 1735 17040
rect 200 17008 800 17038
rect 1669 17035 1735 17038
rect 37590 17036 37596 17100
rect 37660 17098 37666 17100
rect 57421 17098 57487 17101
rect 37660 17096 57487 17098
rect 37660 17040 57426 17096
rect 57482 17040 57487 17096
rect 37660 17038 57487 17040
rect 37660 17036 37666 17038
rect 57421 17035 57487 17038
rect 58249 17098 58315 17101
rect 59200 17098 59800 17128
rect 58249 17096 59800 17098
rect 58249 17040 58254 17096
rect 58310 17040 59800 17096
rect 58249 17038 59800 17040
rect 58249 17035 58315 17038
rect 59200 17008 59800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 43437 16690 43503 16693
rect 44582 16690 44588 16692
rect 43437 16688 44588 16690
rect 43437 16632 43442 16688
rect 43498 16632 44588 16688
rect 43437 16630 44588 16632
rect 43437 16627 43503 16630
rect 44582 16628 44588 16630
rect 44652 16628 44658 16692
rect 34237 16554 34303 16557
rect 41229 16554 41295 16557
rect 43713 16556 43779 16557
rect 43662 16554 43668 16556
rect 34237 16552 43668 16554
rect 43732 16554 43779 16556
rect 43732 16552 43824 16554
rect 34237 16496 34242 16552
rect 34298 16496 41234 16552
rect 41290 16496 43668 16552
rect 43774 16496 43824 16552
rect 34237 16494 43668 16496
rect 34237 16491 34303 16494
rect 41229 16491 41295 16494
rect 43662 16492 43668 16494
rect 43732 16494 43824 16496
rect 43732 16492 43779 16494
rect 43713 16491 43779 16492
rect 40350 16356 40356 16420
rect 40420 16418 40426 16420
rect 40493 16418 40559 16421
rect 40420 16416 40559 16418
rect 40420 16360 40498 16416
rect 40554 16360 40559 16416
rect 40420 16358 40559 16360
rect 40420 16356 40426 16358
rect 40493 16355 40559 16358
rect 43345 16418 43411 16421
rect 44214 16418 44220 16420
rect 43345 16416 44220 16418
rect 43345 16360 43350 16416
rect 43406 16360 44220 16416
rect 43345 16358 44220 16360
rect 43345 16355 43411 16358
rect 44214 16356 44220 16358
rect 44284 16356 44290 16420
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 36629 16146 36695 16149
rect 39297 16146 39363 16149
rect 36629 16144 39363 16146
rect 36629 16088 36634 16144
rect 36690 16088 39302 16144
rect 39358 16088 39363 16144
rect 36629 16086 39363 16088
rect 36629 16083 36695 16086
rect 39297 16083 39363 16086
rect 35617 16010 35683 16013
rect 41873 16010 41939 16013
rect 35617 16008 41939 16010
rect 35617 15952 35622 16008
rect 35678 15952 41878 16008
rect 41934 15952 41939 16008
rect 35617 15950 41939 15952
rect 35617 15947 35683 15950
rect 41873 15947 41939 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 40217 15738 40283 15741
rect 43294 15738 43300 15740
rect 40217 15736 43300 15738
rect 40217 15680 40222 15736
rect 40278 15680 43300 15736
rect 40217 15678 43300 15680
rect 40217 15675 40283 15678
rect 43294 15676 43300 15678
rect 43364 15676 43370 15740
rect 42517 15602 42583 15605
rect 43110 15602 43116 15604
rect 42517 15600 43116 15602
rect 42517 15544 42522 15600
rect 42578 15544 43116 15600
rect 42517 15542 43116 15544
rect 42517 15539 42583 15542
rect 43110 15540 43116 15542
rect 43180 15540 43186 15604
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 35341 15194 35407 15197
rect 40217 15194 40283 15197
rect 35341 15192 40283 15194
rect 35341 15136 35346 15192
rect 35402 15136 40222 15192
rect 40278 15136 40283 15192
rect 35341 15134 40283 15136
rect 35341 15131 35407 15134
rect 40217 15131 40283 15134
rect 40677 15194 40743 15197
rect 44398 15194 44404 15196
rect 40677 15192 44404 15194
rect 40677 15136 40682 15192
rect 40738 15136 44404 15192
rect 40677 15134 44404 15136
rect 40677 15131 40743 15134
rect 44398 15132 44404 15134
rect 44468 15132 44474 15196
rect 39757 15058 39823 15061
rect 40217 15058 40283 15061
rect 39757 15056 40283 15058
rect 39757 15000 39762 15056
rect 39818 15000 40222 15056
rect 40278 15000 40283 15056
rect 39757 14998 40283 15000
rect 39757 14995 39823 14998
rect 40217 14995 40283 14998
rect 40534 14996 40540 15060
rect 40604 15058 40610 15060
rect 41597 15058 41663 15061
rect 40604 15056 41663 15058
rect 40604 15000 41602 15056
rect 41658 15000 41663 15056
rect 40604 14998 41663 15000
rect 40604 14996 40610 14998
rect 41597 14995 41663 14998
rect 28257 14922 28323 14925
rect 38561 14922 38627 14925
rect 28257 14920 38627 14922
rect 28257 14864 28262 14920
rect 28318 14864 38566 14920
rect 38622 14864 38627 14920
rect 28257 14862 38627 14864
rect 28257 14859 28323 14862
rect 38561 14859 38627 14862
rect 39481 14922 39547 14925
rect 40861 14922 40927 14925
rect 41781 14922 41847 14925
rect 39481 14920 41847 14922
rect 39481 14864 39486 14920
rect 39542 14864 40866 14920
rect 40922 14864 41786 14920
rect 41842 14864 41847 14920
rect 39481 14862 41847 14864
rect 39481 14859 39547 14862
rect 40861 14859 40927 14862
rect 41781 14859 41847 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 36169 14514 36235 14517
rect 38561 14514 38627 14517
rect 36169 14512 38627 14514
rect 36169 14456 36174 14512
rect 36230 14456 38566 14512
rect 38622 14456 38627 14512
rect 36169 14454 38627 14456
rect 36169 14451 36235 14454
rect 38561 14451 38627 14454
rect 39205 14514 39271 14517
rect 39205 14512 41016 14514
rect 39205 14456 39210 14512
rect 39266 14456 41016 14512
rect 39205 14454 41016 14456
rect 39205 14451 39271 14454
rect 38653 14378 38719 14381
rect 39849 14378 39915 14381
rect 38653 14376 39915 14378
rect 38653 14320 38658 14376
rect 38714 14320 39854 14376
rect 39910 14320 39915 14376
rect 38653 14318 39915 14320
rect 38653 14315 38719 14318
rect 39849 14315 39915 14318
rect 40956 14245 41016 14454
rect 34421 14242 34487 14245
rect 40166 14242 40172 14244
rect 34421 14240 40172 14242
rect 34421 14184 34426 14240
rect 34482 14184 40172 14240
rect 34421 14182 40172 14184
rect 34421 14179 34487 14182
rect 40166 14180 40172 14182
rect 40236 14180 40242 14244
rect 40953 14240 41019 14245
rect 40953 14184 40958 14240
rect 41014 14184 41019 14240
rect 40953 14179 41019 14184
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 31201 14106 31267 14109
rect 40677 14106 40743 14109
rect 31201 14104 40743 14106
rect 31201 14048 31206 14104
rect 31262 14048 40682 14104
rect 40738 14048 40743 14104
rect 31201 14046 40743 14048
rect 31201 14043 31267 14046
rect 40677 14043 40743 14046
rect 37917 13970 37983 13973
rect 38285 13970 38351 13973
rect 37917 13968 38351 13970
rect 37917 13912 37922 13968
rect 37978 13912 38290 13968
rect 38346 13912 38351 13968
rect 37917 13910 38351 13912
rect 37917 13907 37983 13910
rect 38285 13907 38351 13910
rect 39665 13970 39731 13973
rect 40401 13970 40467 13973
rect 41965 13970 42031 13973
rect 44357 13970 44423 13973
rect 39665 13968 44423 13970
rect 39665 13912 39670 13968
rect 39726 13912 40406 13968
rect 40462 13912 41970 13968
rect 42026 13912 44362 13968
rect 44418 13912 44423 13968
rect 39665 13910 44423 13912
rect 39665 13907 39731 13910
rect 40401 13907 40467 13910
rect 41965 13907 42031 13910
rect 44357 13907 44423 13910
rect 34237 13834 34303 13837
rect 38469 13834 38535 13837
rect 34237 13832 38535 13834
rect 34237 13776 34242 13832
rect 34298 13776 38474 13832
rect 38530 13776 38535 13832
rect 34237 13774 38535 13776
rect 34237 13771 34303 13774
rect 38469 13771 38535 13774
rect 38929 13834 38995 13837
rect 40350 13834 40356 13836
rect 38929 13832 40356 13834
rect 38929 13776 38934 13832
rect 38990 13776 40356 13832
rect 38929 13774 40356 13776
rect 38929 13771 38995 13774
rect 40350 13772 40356 13774
rect 40420 13834 40426 13836
rect 40677 13834 40743 13837
rect 40420 13832 40743 13834
rect 40420 13776 40682 13832
rect 40738 13776 40743 13832
rect 40420 13774 40743 13776
rect 40420 13772 40426 13774
rect 40677 13771 40743 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 40309 13562 40375 13565
rect 42057 13562 42123 13565
rect 40309 13560 42123 13562
rect 40309 13504 40314 13560
rect 40370 13504 42062 13560
rect 42118 13504 42123 13560
rect 40309 13502 42123 13504
rect 40309 13499 40375 13502
rect 42057 13499 42123 13502
rect 36721 13428 36787 13429
rect 36670 13364 36676 13428
rect 36740 13426 36787 13428
rect 36740 13424 36832 13426
rect 36782 13368 36832 13424
rect 36740 13366 36832 13368
rect 36740 13364 36787 13366
rect 36721 13363 36787 13364
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 200 11658 800 11688
rect 1669 11658 1735 11661
rect 200 11656 1735 11658
rect 200 11600 1674 11656
rect 1730 11600 1735 11656
rect 200 11598 1735 11600
rect 200 11568 800 11598
rect 1669 11595 1735 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 58249 10978 58315 10981
rect 59200 10978 59800 11008
rect 58249 10976 59800 10978
rect 58249 10920 58254 10976
rect 58310 10920 59800 10976
rect 58249 10918 59800 10920
rect 58249 10915 58315 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 59800 10918
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 58249 5538 58315 5541
rect 59200 5538 59800 5568
rect 58249 5536 59800 5538
rect 58249 5480 58254 5536
rect 58310 5480 59800 5536
rect 58249 5478 59800 5480
rect 58249 5475 58315 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 59200 5448 59800 5478
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 36854 2620 36860 2684
rect 36924 2682 36930 2684
rect 44081 2682 44147 2685
rect 36924 2680 44147 2682
rect 36924 2624 44086 2680
rect 44142 2624 44147 2680
rect 36924 2622 44147 2624
rect 36924 2620 36930 2622
rect 44081 2619 44147 2622
rect 17677 2546 17743 2549
rect 31518 2546 31524 2548
rect 17677 2544 31524 2546
rect 17677 2488 17682 2544
rect 17738 2488 31524 2544
rect 17677 2486 31524 2488
rect 17677 2483 17743 2486
rect 31518 2484 31524 2486
rect 31588 2484 31594 2548
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 30604 56672 30668 56676
rect 30604 56616 30618 56672
rect 30618 56616 30668 56672
rect 30604 56612 30668 56616
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 22140 47016 22204 47020
rect 22140 46960 22154 47016
rect 22154 46960 22204 47016
rect 22140 46956 22204 46960
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 33732 45732 33796 45796
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 23428 45324 23492 45388
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 33732 44916 33796 44980
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 22876 44236 22940 44300
rect 24348 44296 24412 44300
rect 24348 44240 24398 44296
rect 24398 44240 24412 44296
rect 24348 44236 24412 44240
rect 24900 44236 24964 44300
rect 26556 44296 26620 44300
rect 26556 44240 26570 44296
rect 26570 44240 26620 44296
rect 26556 44236 26620 44240
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 28948 42876 29012 42940
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 27476 41984 27540 41988
rect 27476 41928 27526 41984
rect 27526 41928 27540 41984
rect 27476 41924 27540 41928
rect 28396 41924 28460 41988
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 29132 41108 29196 41172
rect 33732 41168 33796 41172
rect 33732 41112 33746 41168
rect 33746 41112 33796 41168
rect 33732 41108 33796 41112
rect 27292 40972 27356 41036
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 27844 40292 27908 40356
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 27660 40156 27724 40220
rect 22140 39944 22204 39948
rect 22140 39888 22190 39944
rect 22190 39888 22204 39944
rect 22140 39884 22204 39888
rect 24900 39748 24964 39812
rect 26556 39748 26620 39812
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 23428 38932 23492 38996
rect 26556 38856 26620 38860
rect 26556 38800 26606 38856
rect 26606 38800 26620 38856
rect 26556 38796 26620 38800
rect 27844 38856 27908 38860
rect 27844 38800 27858 38856
rect 27858 38800 27908 38856
rect 27844 38796 27908 38800
rect 24716 38660 24780 38724
rect 27292 38660 27356 38724
rect 31156 38720 31220 38724
rect 31156 38664 31170 38720
rect 31170 38664 31220 38720
rect 31156 38660 31220 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 28948 37980 29012 38044
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 27660 37028 27724 37092
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 22876 35864 22940 35868
rect 22876 35808 22890 35864
rect 22890 35808 22940 35864
rect 22876 35804 22940 35808
rect 24348 35804 24412 35868
rect 29132 35728 29196 35732
rect 29132 35672 29182 35728
rect 29182 35672 29196 35728
rect 29132 35668 29196 35672
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 27476 34444 27540 34508
rect 28396 34308 28460 34372
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 37596 31996 37660 32060
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 31156 31316 31220 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 24716 30832 24780 30836
rect 24716 30776 24730 30832
rect 24730 30776 24780 30832
rect 24716 30772 24780 30776
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 36860 26752 36924 26756
rect 36860 26696 36874 26752
rect 36874 26696 36924 26752
rect 36860 26692 36924 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 30604 26420 30668 26484
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 31524 25060 31588 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 31524 23564 31588 23628
rect 39988 23428 40052 23492
rect 44588 23488 44652 23492
rect 44588 23432 44602 23488
rect 44602 23432 44652 23488
rect 44588 23428 44652 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 40172 22476 40236 22540
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 43116 22264 43180 22268
rect 43116 22208 43130 22264
rect 43130 22208 43180 22264
rect 43116 22204 43180 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 40540 20768 40604 20772
rect 40540 20712 40554 20768
rect 40554 20712 40604 20768
rect 40540 20708 40604 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 44220 20164 44284 20228
rect 44404 19892 44468 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 36676 19408 36740 19412
rect 36676 19352 36690 19408
rect 36690 19352 36740 19408
rect 36676 19348 36740 19352
rect 39988 19348 40052 19412
rect 43668 19408 43732 19412
rect 43668 19352 43682 19408
rect 43682 19352 43732 19408
rect 43668 19348 43732 19352
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 43300 18804 43364 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 37596 17036 37660 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 44588 16628 44652 16692
rect 43668 16552 43732 16556
rect 43668 16496 43718 16552
rect 43718 16496 43732 16552
rect 43668 16492 43732 16496
rect 40356 16356 40420 16420
rect 44220 16356 44284 16420
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 43300 15676 43364 15740
rect 43116 15540 43180 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 44404 15132 44468 15196
rect 40540 14996 40604 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 40172 14180 40236 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 40356 13772 40420 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 36676 13424 36740 13428
rect 36676 13368 36726 13424
rect 36726 13368 36740 13424
rect 36676 13364 36740 13368
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 36860 2620 36924 2684
rect 31524 2484 31588 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 30603 56676 30669 56677
rect 30603 56612 30604 56676
rect 30668 56612 30669 56676
rect 30603 56611 30669 56612
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 22139 47020 22205 47021
rect 22139 46956 22140 47020
rect 22204 46956 22205 47020
rect 22139 46955 22205 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 22142 39949 22202 46955
rect 23427 45388 23493 45389
rect 23427 45324 23428 45388
rect 23492 45324 23493 45388
rect 23427 45323 23493 45324
rect 22875 44300 22941 44301
rect 22875 44236 22876 44300
rect 22940 44236 22941 44300
rect 22875 44235 22941 44236
rect 22139 39948 22205 39949
rect 22139 39884 22140 39948
rect 22204 39884 22205 39948
rect 22139 39883 22205 39884
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 22878 35869 22938 44235
rect 23430 38997 23490 45323
rect 24347 44300 24413 44301
rect 24347 44236 24348 44300
rect 24412 44236 24413 44300
rect 24347 44235 24413 44236
rect 24899 44300 24965 44301
rect 24899 44236 24900 44300
rect 24964 44236 24965 44300
rect 24899 44235 24965 44236
rect 26555 44300 26621 44301
rect 26555 44236 26556 44300
rect 26620 44236 26621 44300
rect 26555 44235 26621 44236
rect 23427 38996 23493 38997
rect 23427 38932 23428 38996
rect 23492 38932 23493 38996
rect 23427 38931 23493 38932
rect 24350 35869 24410 44235
rect 24902 39813 24962 44235
rect 26558 39813 26618 44235
rect 28947 42940 29013 42941
rect 28947 42876 28948 42940
rect 29012 42876 29013 42940
rect 28947 42875 29013 42876
rect 27475 41988 27541 41989
rect 27475 41924 27476 41988
rect 27540 41924 27541 41988
rect 27475 41923 27541 41924
rect 28395 41988 28461 41989
rect 28395 41924 28396 41988
rect 28460 41924 28461 41988
rect 28395 41923 28461 41924
rect 27291 41036 27357 41037
rect 27291 40972 27292 41036
rect 27356 40972 27357 41036
rect 27291 40971 27357 40972
rect 24899 39812 24965 39813
rect 24899 39748 24900 39812
rect 24964 39748 24965 39812
rect 24899 39747 24965 39748
rect 26555 39812 26621 39813
rect 26555 39748 26556 39812
rect 26620 39748 26621 39812
rect 26555 39747 26621 39748
rect 26558 38861 26618 39747
rect 26555 38860 26621 38861
rect 26555 38796 26556 38860
rect 26620 38796 26621 38860
rect 26555 38795 26621 38796
rect 27294 38725 27354 40971
rect 24715 38724 24781 38725
rect 24715 38660 24716 38724
rect 24780 38660 24781 38724
rect 24715 38659 24781 38660
rect 27291 38724 27357 38725
rect 27291 38660 27292 38724
rect 27356 38660 27357 38724
rect 27291 38659 27357 38660
rect 22875 35868 22941 35869
rect 22875 35804 22876 35868
rect 22940 35804 22941 35868
rect 22875 35803 22941 35804
rect 24347 35868 24413 35869
rect 24347 35804 24348 35868
rect 24412 35804 24413 35868
rect 24347 35803 24413 35804
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 24718 30837 24778 38659
rect 27478 34509 27538 41923
rect 27843 40356 27909 40357
rect 27843 40292 27844 40356
rect 27908 40292 27909 40356
rect 27843 40291 27909 40292
rect 27659 40220 27725 40221
rect 27659 40156 27660 40220
rect 27724 40156 27725 40220
rect 27659 40155 27725 40156
rect 27662 37093 27722 40155
rect 27846 38861 27906 40291
rect 27843 38860 27909 38861
rect 27843 38796 27844 38860
rect 27908 38796 27909 38860
rect 27843 38795 27909 38796
rect 27659 37092 27725 37093
rect 27659 37028 27660 37092
rect 27724 37028 27725 37092
rect 27659 37027 27725 37028
rect 27475 34508 27541 34509
rect 27475 34444 27476 34508
rect 27540 34444 27541 34508
rect 27475 34443 27541 34444
rect 28398 34373 28458 41923
rect 28950 38045 29010 42875
rect 29131 41172 29197 41173
rect 29131 41108 29132 41172
rect 29196 41108 29197 41172
rect 29131 41107 29197 41108
rect 28947 38044 29013 38045
rect 28947 37980 28948 38044
rect 29012 37980 29013 38044
rect 28947 37979 29013 37980
rect 29134 35733 29194 41107
rect 29131 35732 29197 35733
rect 29131 35668 29132 35732
rect 29196 35668 29197 35732
rect 29131 35667 29197 35668
rect 28395 34372 28461 34373
rect 28395 34308 28396 34372
rect 28460 34308 28461 34372
rect 28395 34307 28461 34308
rect 24715 30836 24781 30837
rect 24715 30772 24716 30836
rect 24780 30772 24781 30836
rect 24715 30771 24781 30772
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 30606 26485 30666 56611
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 33731 45796 33797 45797
rect 33731 45732 33732 45796
rect 33796 45732 33797 45796
rect 33731 45731 33797 45732
rect 33734 44981 33794 45731
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 33731 44980 33797 44981
rect 33731 44916 33732 44980
rect 33796 44916 33797 44980
rect 33731 44915 33797 44916
rect 33734 41173 33794 44915
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 33731 41172 33797 41173
rect 33731 41108 33732 41172
rect 33796 41108 33797 41172
rect 33731 41107 33797 41108
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 31155 38724 31221 38725
rect 31155 38660 31156 38724
rect 31220 38660 31221 38724
rect 31155 38659 31221 38660
rect 31158 31381 31218 38659
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 31155 31380 31221 31381
rect 31155 31316 31156 31380
rect 31220 31316 31221 31380
rect 31155 31315 31221 31316
rect 34928 31040 35248 32064
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 37595 32060 37661 32061
rect 37595 31996 37596 32060
rect 37660 31996 37661 32060
rect 37595 31995 37661 31996
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 36859 26756 36925 26757
rect 36859 26692 36860 26756
rect 36924 26692 36925 26756
rect 36859 26691 36925 26692
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 30603 26484 30669 26485
rect 30603 26420 30604 26484
rect 30668 26420 30669 26484
rect 30603 26419 30669 26420
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 31523 25124 31589 25125
rect 31523 25060 31524 25124
rect 31588 25060 31589 25124
rect 31523 25059 31589 25060
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 31526 23629 31586 25059
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 31523 23628 31589 23629
rect 31523 23564 31524 23628
rect 31588 23564 31589 23628
rect 31523 23563 31589 23564
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 31526 2549 31586 23563
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 36675 19412 36741 19413
rect 36675 19348 36676 19412
rect 36740 19348 36741 19412
rect 36675 19347 36741 19348
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 36678 13429 36738 19347
rect 36675 13428 36741 13429
rect 36675 13364 36676 13428
rect 36740 13364 36741 13428
rect 36675 13363 36741 13364
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 31523 2548 31589 2549
rect 31523 2484 31524 2548
rect 31588 2484 31589 2548
rect 31523 2483 31589 2484
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 36862 2685 36922 26691
rect 37598 17101 37658 31995
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 39987 23492 40053 23493
rect 39987 23428 39988 23492
rect 40052 23428 40053 23492
rect 39987 23427 40053 23428
rect 44587 23492 44653 23493
rect 44587 23428 44588 23492
rect 44652 23428 44653 23492
rect 44587 23427 44653 23428
rect 39990 19413 40050 23427
rect 40171 22540 40237 22541
rect 40171 22476 40172 22540
rect 40236 22476 40237 22540
rect 40171 22475 40237 22476
rect 39987 19412 40053 19413
rect 39987 19348 39988 19412
rect 40052 19348 40053 19412
rect 39987 19347 40053 19348
rect 37595 17100 37661 17101
rect 37595 17036 37596 17100
rect 37660 17036 37661 17100
rect 37595 17035 37661 17036
rect 40174 14245 40234 22475
rect 43115 22268 43181 22269
rect 43115 22204 43116 22268
rect 43180 22204 43181 22268
rect 43115 22203 43181 22204
rect 40539 20772 40605 20773
rect 40539 20708 40540 20772
rect 40604 20708 40605 20772
rect 40539 20707 40605 20708
rect 40355 16420 40421 16421
rect 40355 16356 40356 16420
rect 40420 16356 40421 16420
rect 40355 16355 40421 16356
rect 40171 14244 40237 14245
rect 40171 14180 40172 14244
rect 40236 14180 40237 14244
rect 40171 14179 40237 14180
rect 40358 13837 40418 16355
rect 40542 15061 40602 20707
rect 43118 15605 43178 22203
rect 44219 20228 44285 20229
rect 44219 20164 44220 20228
rect 44284 20164 44285 20228
rect 44219 20163 44285 20164
rect 43667 19412 43733 19413
rect 43667 19348 43668 19412
rect 43732 19348 43733 19412
rect 43667 19347 43733 19348
rect 43299 18868 43365 18869
rect 43299 18804 43300 18868
rect 43364 18804 43365 18868
rect 43299 18803 43365 18804
rect 43302 15741 43362 18803
rect 43670 16557 43730 19347
rect 43667 16556 43733 16557
rect 43667 16492 43668 16556
rect 43732 16492 43733 16556
rect 43667 16491 43733 16492
rect 44222 16421 44282 20163
rect 44403 19956 44469 19957
rect 44403 19892 44404 19956
rect 44468 19892 44469 19956
rect 44403 19891 44469 19892
rect 44219 16420 44285 16421
rect 44219 16356 44220 16420
rect 44284 16356 44285 16420
rect 44219 16355 44285 16356
rect 43299 15740 43365 15741
rect 43299 15676 43300 15740
rect 43364 15676 43365 15740
rect 43299 15675 43365 15676
rect 43115 15604 43181 15605
rect 43115 15540 43116 15604
rect 43180 15540 43181 15604
rect 43115 15539 43181 15540
rect 44406 15197 44466 19891
rect 44590 16693 44650 23427
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 44587 16692 44653 16693
rect 44587 16628 44588 16692
rect 44652 16628 44653 16692
rect 44587 16627 44653 16628
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 44403 15196 44469 15197
rect 44403 15132 44404 15196
rect 44468 15132 44469 15196
rect 44403 15131 44469 15132
rect 40539 15060 40605 15061
rect 40539 14996 40540 15060
rect 40604 14996 40605 15060
rect 40539 14995 40605 14996
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 40355 13836 40421 13837
rect 40355 13772 40356 13836
rect 40420 13772 40421 13836
rect 40355 13771 40421 13772
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 36859 2684 36925 2685
rect 36859 2620 36860 2684
rect 36924 2620 36925 2684
rect 36859 2619 36925 2620
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1666464484
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A2
timestamp 1666464484
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B1
timestamp 1666464484
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A_N
timestamp 1666464484
transform 1 0 40572 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1666464484
transform 1 0 42688 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A_N
timestamp 1666464484
transform 1 0 36800 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B
timestamp 1666464484
transform 1 0 39376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A2
timestamp 1666464484
transform 1 0 41860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B1
timestamp 1666464484
transform 1 0 41584 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1666464484
transform -1 0 40848 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1666464484
transform -1 0 42964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1666464484
transform 1 0 27416 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1666464484
transform 1 0 29716 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1666464484
transform 1 0 22356 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1666464484
transform 1 0 35512 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B1
timestamp 1666464484
transform 1 0 21344 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1666464484
transform 1 0 33856 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1666464484
transform -1 0 31372 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1666464484
transform 1 0 34040 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1666464484
transform 1 0 34592 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1666464484
transform 1 0 31556 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__C
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B
timestamp 1666464484
transform -1 0 26404 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1666464484
transform 1 0 36248 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B
timestamp 1666464484
transform 1 0 30176 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1666464484
transform 1 0 34132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1666464484
transform -1 0 31188 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1666464484
transform 1 0 28244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A_N
timestamp 1666464484
transform -1 0 31556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__S
timestamp 1666464484
transform 1 0 26772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__S
timestamp 1666464484
transform -1 0 26404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1666464484
transform 1 0 18768 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__S
timestamp 1666464484
transform -1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1666464484
transform -1 0 29072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B
timestamp 1666464484
transform 1 0 26312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1666464484
transform 1 0 27784 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1666464484
transform 1 0 25668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1666464484
transform -1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1666464484
transform -1 0 26128 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1666464484
transform 1 0 34868 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1666464484
transform 1 0 32476 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A2
timestamp 1666464484
transform 1 0 34868 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B1_N
timestamp 1666464484
transform 1 0 34132 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1666464484
transform 1 0 21344 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B
timestamp 1666464484
transform 1 0 35696 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1666464484
transform 1 0 27876 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1666464484
transform 1 0 17664 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1666464484
transform -1 0 29072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A2
timestamp 1666464484
transform -1 0 19412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1666464484
transform 1 0 19688 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1666464484
transform 1 0 25760 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1666464484
transform 1 0 21068 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A1
timestamp 1666464484
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1666464484
transform 1 0 27600 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B
timestamp 1666464484
transform -1 0 19872 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B
timestamp 1666464484
transform 1 0 35880 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1
timestamp 1666464484
transform 1 0 34684 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A2
timestamp 1666464484
transform -1 0 23828 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B1
timestamp 1666464484
transform 1 0 23920 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 1666464484
transform 1 0 20516 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1666464484
transform 1 0 30176 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1666464484
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1666464484
transform 1 0 18676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1666464484
transform 1 0 19688 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A3
timestamp 1666464484
transform 1 0 20884 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1666464484
transform -1 0 20700 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1666464484
transform 1 0 28980 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__B
timestamp 1666464484
transform 1 0 29072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1666464484
transform 1 0 19044 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1666464484
transform 1 0 18216 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1666464484
transform 1 0 25852 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A1
timestamp 1666464484
transform 1 0 26404 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B1
timestamp 1666464484
transform 1 0 30268 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B
timestamp 1666464484
transform -1 0 29440 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__B2
timestamp 1666464484
transform 1 0 25208 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1666464484
transform -1 0 16560 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B
timestamp 1666464484
transform -1 0 29900 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__B1
timestamp 1666464484
transform 1 0 31556 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1666464484
transform 1 0 31464 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1666464484
transform 1 0 27968 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B
timestamp 1666464484
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1666464484
transform 1 0 28888 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 1666464484
transform 1 0 26128 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A
timestamp 1666464484
transform 1 0 20332 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A2
timestamp 1666464484
transform -1 0 23092 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B1
timestamp 1666464484
transform 1 0 23920 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B1
timestamp 1666464484
transform 1 0 23736 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A
timestamp 1666464484
transform -1 0 29348 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B1
timestamp 1666464484
transform 1 0 23184 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1666464484
transform -1 0 19320 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1666464484
transform -1 0 20976 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A1
timestamp 1666464484
transform -1 0 18768 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B2
timestamp 1666464484
transform -1 0 17940 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1666464484
transform 1 0 31648 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A1
timestamp 1666464484
transform -1 0 24932 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A
timestamp 1666464484
transform 1 0 23552 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1666464484
transform -1 0 26864 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__C_N
timestamp 1666464484
transform 1 0 17112 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A3
timestamp 1666464484
transform -1 0 18676 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A1
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B1
timestamp 1666464484
transform -1 0 28336 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A
timestamp 1666464484
transform -1 0 25668 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1666464484
transform -1 0 29164 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B
timestamp 1666464484
transform 1 0 31188 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A1
timestamp 1666464484
transform 1 0 28796 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1666464484
transform 1 0 19412 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A2
timestamp 1666464484
transform -1 0 20148 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A1
timestamp 1666464484
transform -1 0 17848 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1666464484
transform -1 0 17388 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1666464484
transform -1 0 17388 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A
timestamp 1666464484
transform 1 0 26220 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A
timestamp 1666464484
transform 1 0 33212 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__C1
timestamp 1666464484
transform -1 0 34868 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A1
timestamp 1666464484
transform 1 0 26496 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A3
timestamp 1666464484
transform 1 0 24932 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1666464484
transform 1 0 30728 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__B
timestamp 1666464484
transform 1 0 20240 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1666464484
transform 1 0 21344 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__B1
timestamp 1666464484
transform -1 0 19872 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1666464484
transform -1 0 23828 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A1
timestamp 1666464484
transform -1 0 21160 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1666464484
transform 1 0 26404 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B
timestamp 1666464484
transform 1 0 24564 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A2
timestamp 1666464484
transform 1 0 28244 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A2
timestamp 1666464484
transform -1 0 27692 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1666464484
transform 1 0 25852 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1666464484
transform -1 0 19780 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1666464484
transform 1 0 21160 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A
timestamp 1666464484
transform 1 0 19964 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1666464484
transform 1 0 31740 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__B
timestamp 1666464484
transform -1 0 33396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__B1
timestamp 1666464484
transform -1 0 25760 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A1
timestamp 1666464484
transform 1 0 21620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A2
timestamp 1666464484
transform 1 0 21344 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B1_N
timestamp 1666464484
transform 1 0 21344 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A3
timestamp 1666464484
transform 1 0 32016 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1666464484
transform 1 0 29440 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__C1
timestamp 1666464484
transform 1 0 31280 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__C1
timestamp 1666464484
transform 1 0 29716 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__C
timestamp 1666464484
transform 1 0 31648 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A2
timestamp 1666464484
transform -1 0 22264 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__B1
timestamp 1666464484
transform 1 0 22724 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A
timestamp 1666464484
transform 1 0 23828 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__B
timestamp 1666464484
transform 1 0 24656 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A
timestamp 1666464484
transform 1 0 30360 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__B
timestamp 1666464484
transform 1 0 30728 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__C1
timestamp 1666464484
transform 1 0 29348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A2
timestamp 1666464484
transform 1 0 30912 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__C1
timestamp 1666464484
transform 1 0 23184 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A
timestamp 1666464484
transform 1 0 30084 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A1
timestamp 1666464484
transform 1 0 24196 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A2
timestamp 1666464484
transform -1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A1
timestamp 1666464484
transform -1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A1
timestamp 1666464484
transform 1 0 31280 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__A1
timestamp 1666464484
transform 1 0 34224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__C1
timestamp 1666464484
transform -1 0 33120 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__A
timestamp 1666464484
transform 1 0 31280 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__B1
timestamp 1666464484
transform 1 0 33580 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A3
timestamp 1666464484
transform -1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__C1
timestamp 1666464484
transform 1 0 34408 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A
timestamp 1666464484
transform -1 0 35052 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__A
timestamp 1666464484
transform 1 0 34040 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__A1
timestamp 1666464484
transform -1 0 35052 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__B1
timestamp 1666464484
transform -1 0 27324 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A3
timestamp 1666464484
transform -1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__A1
timestamp 1666464484
transform 1 0 34224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__C1
timestamp 1666464484
transform -1 0 34684 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A
timestamp 1666464484
transform -1 0 35880 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__A
timestamp 1666464484
transform -1 0 29624 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__A
timestamp 1666464484
transform -1 0 42044 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__A
timestamp 1666464484
transform -1 0 46368 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A
timestamp 1666464484
transform 1 0 44436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__A1
timestamp 1666464484
transform 1 0 46000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__A
timestamp 1666464484
transform 1 0 41400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__B
timestamp 1666464484
transform -1 0 40204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__B_N
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__A
timestamp 1666464484
transform -1 0 37168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__A3
timestamp 1666464484
transform -1 0 40204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__B1_N
timestamp 1666464484
transform 1 0 45908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__A1_N
timestamp 1666464484
transform 1 0 45632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__A
timestamp 1666464484
transform 1 0 37996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__B1
timestamp 1666464484
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__A1
timestamp 1666464484
transform 1 0 41952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__A3
timestamp 1666464484
transform 1 0 44436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1608__B1
timestamp 1666464484
transform -1 0 46368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__A
timestamp 1666464484
transform -1 0 45356 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1617__A
timestamp 1666464484
transform 1 0 45172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1619__C1
timestamp 1666464484
transform 1 0 45632 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__A
timestamp 1666464484
transform 1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1630__B1
timestamp 1666464484
transform -1 0 46460 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1632__A
timestamp 1666464484
transform 1 0 44252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1635__B1
timestamp 1666464484
transform -1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1637__A
timestamp 1666464484
transform 1 0 32476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1638__A1
timestamp 1666464484
transform 1 0 33028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1645__A
timestamp 1666464484
transform -1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__C1
timestamp 1666464484
transform 1 0 44344 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1651__A1
timestamp 1666464484
transform -1 0 38456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__A1
timestamp 1666464484
transform -1 0 41768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1655__A1
timestamp 1666464484
transform -1 0 41032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1655__B1
timestamp 1666464484
transform -1 0 41952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1660__A2
timestamp 1666464484
transform -1 0 31924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1660__B1
timestamp 1666464484
transform -1 0 27048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1661__B
timestamp 1666464484
transform 1 0 27876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1661__C
timestamp 1666464484
transform 1 0 27324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1662__A
timestamp 1666464484
transform 1 0 29716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1664__A
timestamp 1666464484
transform -1 0 42044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1665__A1
timestamp 1666464484
transform -1 0 46368 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1669__A
timestamp 1666464484
transform -1 0 42780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1681__C1
timestamp 1666464484
transform 1 0 32016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1689__A
timestamp 1666464484
transform 1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1694__A
timestamp 1666464484
transform 1 0 36156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__C
timestamp 1666464484
transform -1 0 41308 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1715__A1
timestamp 1666464484
transform 1 0 43240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1719__B1
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1720__B
timestamp 1666464484
transform -1 0 33304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1722__B1
timestamp 1666464484
transform -1 0 37996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1724__A
timestamp 1666464484
transform 1 0 41768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1734__A
timestamp 1666464484
transform -1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1737__B1
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1747__D_N
timestamp 1666464484
transform 1 0 34224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1749__A
timestamp 1666464484
transform 1 0 41952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1751__A
timestamp 1666464484
transform 1 0 40940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1754__A3
timestamp 1666464484
transform 1 0 38272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1759__B
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1764__A1
timestamp 1666464484
transform 1 0 36616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1764__A2
timestamp 1666464484
transform 1 0 35328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1773__A
timestamp 1666464484
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1776__A
timestamp 1666464484
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1792__A2
timestamp 1666464484
transform -1 0 33212 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1795__B2
timestamp 1666464484
transform 1 0 33856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__A_N
timestamp 1666464484
transform -1 0 28704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__C_N
timestamp 1666464484
transform 1 0 41032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1828__A
timestamp 1666464484
transform -1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1838__A1
timestamp 1666464484
transform 1 0 41216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1844__B2
timestamp 1666464484
transform -1 0 40204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1855__A
timestamp 1666464484
transform 1 0 28520 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1862__A
timestamp 1666464484
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1863__C
timestamp 1666464484
transform 1 0 36616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__A
timestamp 1666464484
transform 1 0 32568 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1875__A1
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__C1
timestamp 1666464484
transform -1 0 29808 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1884__A1
timestamp 1666464484
transform 1 0 38548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1894__C1
timestamp 1666464484
transform 1 0 31464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1906__A1
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1923__A
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__A1
timestamp 1666464484
transform 1 0 33396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1939__A
timestamp 1666464484
transform 1 0 29072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1940__A1
timestamp 1666464484
transform 1 0 27416 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1942__A2
timestamp 1666464484
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1943__B2
timestamp 1666464484
transform 1 0 34224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1946__B1
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1956__A1
timestamp 1666464484
transform 1 0 34868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1971__A1
timestamp 1666464484
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1972__A
timestamp 1666464484
transform 1 0 26312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1975__B
timestamp 1666464484
transform 1 0 28336 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1977__B
timestamp 1666464484
transform -1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1979__A
timestamp 1666464484
transform 1 0 34960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1979__B
timestamp 1666464484
transform 1 0 33028 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__A
timestamp 1666464484
transform -1 0 33488 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__C
timestamp 1666464484
transform 1 0 32752 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1982__B
timestamp 1666464484
transform 1 0 36708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1984__A1
timestamp 1666464484
transform 1 0 38088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1984__B2
timestamp 1666464484
transform -1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1985__B
timestamp 1666464484
transform 1 0 37904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1986__A2
timestamp 1666464484
transform -1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1991__A1
timestamp 1666464484
transform 1 0 35880 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1992__A
timestamp 1666464484
transform 1 0 32568 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1993__A
timestamp 1666464484
transform -1 0 36616 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1994__A1
timestamp 1666464484
transform 1 0 32660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1995__B
timestamp 1666464484
transform -1 0 36248 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1996__A
timestamp 1666464484
transform -1 0 35972 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1997__A1
timestamp 1666464484
transform -1 0 34316 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1997__A2
timestamp 1666464484
transform -1 0 36432 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1997__A3
timestamp 1666464484
transform 1 0 34868 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2000__C
timestamp 1666464484
transform 1 0 35512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2001__A2
timestamp 1666464484
transform 1 0 32660 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2005__A1
timestamp 1666464484
transform -1 0 36708 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2006__A
timestamp 1666464484
transform -1 0 34960 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2007__A2
timestamp 1666464484
transform 1 0 32108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2008__A
timestamp 1666464484
transform -1 0 27508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2009__A
timestamp 1666464484
transform 1 0 26496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2012__CLK
timestamp 1666464484
transform 1 0 27232 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2013__CLK
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2016__CLK
timestamp 1666464484
transform 1 0 29072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2016__RESET_B
timestamp 1666464484
transform 1 0 28520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2024__CLK
timestamp 1666464484
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2024__RESET_B
timestamp 1666464484
transform 1 0 28980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2027__SET_B
timestamp 1666464484
transform -1 0 35696 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2028__RESET_B
timestamp 1666464484
transform -1 0 35052 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2029__RESET_B
timestamp 1666464484
transform 1 0 35696 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2030__SET_B
timestamp 1666464484
transform 1 0 36064 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2031__SET_B
timestamp 1666464484
transform 1 0 35972 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2033__D
timestamp 1666464484
transform 1 0 24564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2034__CLK
timestamp 1666464484
transform -1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2034__RESET_B
timestamp 1666464484
transform 1 0 30452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__CLK
timestamp 1666464484
transform -1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__D
timestamp 1666464484
transform -1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__RESET_B
timestamp 1666464484
transform -1 0 28244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout44_A
timestamp 1666464484
transform 1 0 35144 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_A
timestamp 1666464484
transform -1 0 39100 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout46_A
timestamp 1666464484
transform -1 0 24288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_A
timestamp 1666464484
transform 1 0 31832 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout48_A
timestamp 1666464484
transform -1 0 23276 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_A
timestamp 1666464484
transform 1 0 27324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout50_A
timestamp 1666464484
transform 1 0 37444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout51_A
timestamp 1666464484
transform -1 0 36708 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 29992 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 2668 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 43516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 57684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_A
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output7_A
timestamp 1666464484
transform 1 0 2300 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1666464484
transform 1 0 57408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_A
timestamp 1666464484
transform 1 0 54832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1666464484
transform -1 0 57684 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output13_A
timestamp 1666464484
transform 1 0 45908 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output14_A
timestamp 1666464484
transform 1 0 2300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output15_A
timestamp 1666464484
transform -1 0 57684 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output16_A
timestamp 1666464484
transform -1 0 2484 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output17_A
timestamp 1666464484
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output18_A
timestamp 1666464484
transform -1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output19_A
timestamp 1666464484
transform -1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output21_A
timestamp 1666464484
transform 1 0 52256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform -1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output23_A
timestamp 1666464484
transform 1 0 57408 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_A
timestamp 1666464484
transform -1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_A
timestamp 1666464484
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1666464484
transform -1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1666464484
transform 1 0 57408 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1666464484
transform 1 0 9844 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 1666464484
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1666464484
transform 1 0 48484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 40756 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1666464484
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 1666464484
transform 1 0 2300 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1666464484
transform -1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1666464484
transform 1 0 27876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1666464484
transform -1 0 57684 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1666464484
transform 1 0 57408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1666464484
transform 1 0 25300 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1666464484
transform 1 0 37536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1666464484
transform -1 0 2484 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output42_A
timestamp 1666464484
transform 1 0 1932 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1666464484
transform -1 0 57592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1666464484
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_231
timestamp 1666464484
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1666464484
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1666464484
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1666464484
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1666464484
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1666464484
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_350
timestamp 1666464484
transform 1 0 33304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1666464484
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1666464484
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1666464484
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_406
timestamp 1666464484
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1666464484
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1666464484
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_457
timestamp 1666464484
transform 1 0 43148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666464484
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1666464484
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1666464484
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_513
timestamp 1666464484
transform 1 0 48300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_517
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_525
timestamp 1666464484
transform 1 0 49404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1666464484
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_573
timestamp 1666464484
transform 1 0 53820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_581
timestamp 1666464484
transform 1 0 54556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1666464484
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_595
timestamp 1666464484
transform 1 0 55844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_607
timestamp 1666464484
transform 1 0 56948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_611
timestamp 1666464484
transform 1 0 57316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1666464484
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1666464484
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1666464484
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1666464484
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1666464484
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1666464484
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1666464484
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1666464484
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1666464484
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1666464484
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1666464484
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1666464484
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1666464484
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1666464484
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1666464484
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1666464484
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1666464484
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1666464484
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1666464484
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1666464484
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1666464484
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1666464484
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1666464484
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1666464484
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1666464484
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666464484
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1666464484
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1666464484
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1666464484
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1666464484
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1666464484
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1666464484
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1666464484
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1666464484
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1666464484
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1666464484
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1666464484
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1666464484
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1666464484
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1666464484
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1666464484
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1666464484
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1666464484
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1666464484
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666464484
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666464484
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666464484
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666464484
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666464484
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666464484
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666464484
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1666464484
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1666464484
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1666464484
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1666464484
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1666464484
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1666464484
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1666464484
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1666464484
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666464484
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666464484
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666464484
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666464484
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666464484
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666464484
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666464484
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1666464484
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1666464484
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1666464484
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1666464484
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1666464484
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1666464484
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1666464484
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666464484
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666464484
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666464484
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666464484
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666464484
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666464484
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666464484
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1666464484
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1666464484
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1666464484
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1666464484
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1666464484
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1666464484
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_615
timestamp 1666464484
transform 1 0 57684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1666464484
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666464484
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666464484
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1666464484
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1666464484
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1666464484
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666464484
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1666464484
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1666464484
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1666464484
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1666464484
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_325
timestamp 1666464484
transform 1 0 31004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1666464484
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_357
timestamp 1666464484
transform 1 0 33948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_369
timestamp 1666464484
transform 1 0 35052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_381
timestamp 1666464484
transform 1 0 36156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1666464484
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666464484
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1666464484
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1666464484
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1666464484
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1666464484
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_295
timestamp 1666464484
transform 1 0 28244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_319
timestamp 1666464484
transform 1 0 30452 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_331
timestamp 1666464484
transform 1 0 31556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_343
timestamp 1666464484
transform 1 0 32660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_351
timestamp 1666464484
transform 1 0 33396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1666464484
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666464484
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666464484
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666464484
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1666464484
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1666464484
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1666464484
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_287
timestamp 1666464484
transform 1 0 27508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_328
timestamp 1666464484
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_347
timestamp 1666464484
transform 1 0 33028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_357
timestamp 1666464484
transform 1 0 33948 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_371
timestamp 1666464484
transform 1 0 35236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1666464484
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_402
timestamp 1666464484
transform 1 0 38088 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_414
timestamp 1666464484
transform 1 0 39192 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_426
timestamp 1666464484
transform 1 0 40296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_438
timestamp 1666464484
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1666464484
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1666464484
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1666464484
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1666464484
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_273
timestamp 1666464484
transform 1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1666464484
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_285
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1666464484
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_315
timestamp 1666464484
transform 1 0 30084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1666464484
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_335
timestamp 1666464484
transform 1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_341
timestamp 1666464484
transform 1 0 32476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_349
timestamp 1666464484
transform 1 0 33212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_353
timestamp 1666464484
transform 1 0 33580 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1666464484
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_371
timestamp 1666464484
transform 1 0 35236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_379
timestamp 1666464484
transform 1 0 35972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_391
timestamp 1666464484
transform 1 0 37076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_395
timestamp 1666464484
transform 1 0 37444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1666464484
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666464484
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1666464484
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1666464484
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1666464484
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1666464484
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1666464484
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_303
timestamp 1666464484
transform 1 0 28980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_309
timestamp 1666464484
transform 1 0 29532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_315
timestamp 1666464484
transform 1 0 30084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_321
timestamp 1666464484
transform 1 0 30636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1666464484
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_343
timestamp 1666464484
transform 1 0 32660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_363
timestamp 1666464484
transform 1 0 34500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_370
timestamp 1666464484
transform 1 0 35144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_377
timestamp 1666464484
transform 1 0 35788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1666464484
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_399
timestamp 1666464484
transform 1 0 37812 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_412
timestamp 1666464484
transform 1 0 39008 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_424
timestamp 1666464484
transform 1 0 40112 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_436
timestamp 1666464484
transform 1 0 41216 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666464484
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666464484
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1666464484
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1666464484
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1666464484
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1666464484
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_281
timestamp 1666464484
transform 1 0 26956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_287
timestamp 1666464484
transform 1 0 27508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_294
timestamp 1666464484
transform 1 0 28152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_300
timestamp 1666464484
transform 1 0 28704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1666464484
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_318
timestamp 1666464484
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_332
timestamp 1666464484
transform 1 0 31648 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_344
timestamp 1666464484
transform 1 0 32752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_350
timestamp 1666464484
transform 1 0 33304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1666464484
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_373
timestamp 1666464484
transform 1 0 35420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_382
timestamp 1666464484
transform 1 0 36248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_395
timestamp 1666464484
transform 1 0 37444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_410
timestamp 1666464484
transform 1 0 38824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1666464484
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_430
timestamp 1666464484
transform 1 0 40664 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_442
timestamp 1666464484
transform 1 0 41768 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_454
timestamp 1666464484
transform 1 0 42872 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_466
timestamp 1666464484
transform 1 0 43976 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1666464484
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666464484
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1666464484
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1666464484
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1666464484
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_303
timestamp 1666464484
transform 1 0 28980 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1666464484
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_344
timestamp 1666464484
transform 1 0 32752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_353
timestamp 1666464484
transform 1 0 33580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_368
timestamp 1666464484
transform 1 0 34960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_375
timestamp 1666464484
transform 1 0 35604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_379
timestamp 1666464484
transform 1 0 35972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_397
timestamp 1666464484
transform 1 0 37628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_409
timestamp 1666464484
transform 1 0 38732 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_418
timestamp 1666464484
transform 1 0 39560 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_430
timestamp 1666464484
transform 1 0 40664 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_442
timestamp 1666464484
transform 1 0 41768 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666464484
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666464484
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1666464484
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1666464484
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1666464484
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1666464484
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1666464484
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1666464484
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1666464484
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1666464484
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_320
timestamp 1666464484
transform 1 0 30544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1666464484
transform 1 0 31648 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_336
timestamp 1666464484
transform 1 0 32016 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_341
timestamp 1666464484
transform 1 0 32476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_347
timestamp 1666464484
transform 1 0 33028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666464484
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1666464484
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1666464484
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1666464484
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_387
timestamp 1666464484
transform 1 0 36708 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1666464484
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666464484
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_415
timestamp 1666464484
transform 1 0 39284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666464484
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666464484
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666464484
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1666464484
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_615
timestamp 1666464484
transform 1 0 57684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_623
timestamp 1666464484
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_257
timestamp 1666464484
transform 1 0 24748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1666464484
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1666464484
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_292
timestamp 1666464484
transform 1 0 27968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_300
timestamp 1666464484
transform 1 0 28704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_306
timestamp 1666464484
transform 1 0 29256 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_312
timestamp 1666464484
transform 1 0 29808 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1666464484
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_322
timestamp 1666464484
transform 1 0 30728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1666464484
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1666464484
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_346
timestamp 1666464484
transform 1 0 32936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_354
timestamp 1666464484
transform 1 0 33672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_367
timestamp 1666464484
transform 1 0 34868 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_373
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_379
timestamp 1666464484
transform 1 0 35972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1666464484
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_411
timestamp 1666464484
transform 1 0 38916 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_421
timestamp 1666464484
transform 1 0 39836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1666464484
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1666464484
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1666464484
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1666464484
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1666464484
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1666464484
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1666464484
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_318
timestamp 1666464484
transform 1 0 30360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1666464484
transform 1 0 31648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_338
timestamp 1666464484
transform 1 0 32200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_349
timestamp 1666464484
transform 1 0 33212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1666464484
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_378
timestamp 1666464484
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1666464484
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1666464484
transform 1 0 37168 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_399
timestamp 1666464484
transform 1 0 37812 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_411
timestamp 1666464484
transform 1 0 38916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666464484
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_429
timestamp 1666464484
transform 1 0 40572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_434
timestamp 1666464484
transform 1 0 41032 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_442
timestamp 1666464484
transform 1 0 41768 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_454
timestamp 1666464484
transform 1 0 42872 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1666464484
transform 1 0 43976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1666464484
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1666464484
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1666464484
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1666464484
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1666464484
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1666464484
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_289
timestamp 1666464484
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1666464484
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_318
timestamp 1666464484
transform 1 0 30360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_327
timestamp 1666464484
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1666464484
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_346
timestamp 1666464484
transform 1 0 32936 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_358
timestamp 1666464484
transform 1 0 34040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_366
timestamp 1666464484
transform 1 0 34776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_372
timestamp 1666464484
transform 1 0 35328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_379
timestamp 1666464484
transform 1 0 35972 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1666464484
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_400
timestamp 1666464484
transform 1 0 37904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_406
timestamp 1666464484
transform 1 0 38456 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_421
timestamp 1666464484
transform 1 0 39836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_438
timestamp 1666464484
transform 1 0 41400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1666464484
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_453
timestamp 1666464484
transform 1 0 42780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_465
timestamp 1666464484
transform 1 0 43884 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_477
timestamp 1666464484
transform 1 0 44988 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_489
timestamp 1666464484
transform 1 0 46092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_501
timestamp 1666464484
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1666464484
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_241
timestamp 1666464484
transform 1 0 23276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1666464484
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_275
timestamp 1666464484
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1666464484
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_297
timestamp 1666464484
transform 1 0 28428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1666464484
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_313
timestamp 1666464484
transform 1 0 29900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1666464484
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1666464484
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1666464484
transform 1 0 31372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_335
timestamp 1666464484
transform 1 0 31924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_341
timestamp 1666464484
transform 1 0 32476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_346
timestamp 1666464484
transform 1 0 32936 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_352
timestamp 1666464484
transform 1 0 33488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1666464484
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_376
timestamp 1666464484
transform 1 0 35696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_391
timestamp 1666464484
transform 1 0 37076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_395
timestamp 1666464484
transform 1 0 37444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_404
timestamp 1666464484
transform 1 0 38272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1666464484
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_432
timestamp 1666464484
transform 1 0 40848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_440
timestamp 1666464484
transform 1 0 41584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_451
timestamp 1666464484
transform 1 0 42596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_462
timestamp 1666464484
transform 1 0 43608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666464484
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1666464484
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_233
timestamp 1666464484
transform 1 0 22540 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1666464484
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_248
timestamp 1666464484
transform 1 0 23920 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_257
timestamp 1666464484
transform 1 0 24748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_267
timestamp 1666464484
transform 1 0 25668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1666464484
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1666464484
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_295
timestamp 1666464484
transform 1 0 28244 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_302
timestamp 1666464484
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_315
timestamp 1666464484
transform 1 0 30084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_323
timestamp 1666464484
transform 1 0 30820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1666464484
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_343
timestamp 1666464484
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_351
timestamp 1666464484
transform 1 0 33396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_359
timestamp 1666464484
transform 1 0 34132 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_362
timestamp 1666464484
transform 1 0 34408 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_373
timestamp 1666464484
transform 1 0 35420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1666464484
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_397
timestamp 1666464484
transform 1 0 37628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_402
timestamp 1666464484
transform 1 0 38088 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_408
timestamp 1666464484
transform 1 0 38640 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_412
timestamp 1666464484
transform 1 0 39008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_420
timestamp 1666464484
transform 1 0 39744 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_428
timestamp 1666464484
transform 1 0 40480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_435
timestamp 1666464484
transform 1 0 41124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1666464484
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_456
timestamp 1666464484
transform 1 0 43056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_464
timestamp 1666464484
transform 1 0 43792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_473
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1666464484
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_486
timestamp 1666464484
transform 1 0 45816 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_498
timestamp 1666464484
transform 1 0 46920 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1666464484
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1666464484
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1666464484
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1666464484
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1666464484
transform 1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1666464484
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1666464484
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1666464484
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1666464484
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_303
timestamp 1666464484
transform 1 0 28980 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1666464484
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_315
timestamp 1666464484
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_325
timestamp 1666464484
transform 1 0 31004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_332
timestamp 1666464484
transform 1 0 31648 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_340
timestamp 1666464484
transform 1 0 32384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_347
timestamp 1666464484
transform 1 0 33028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_355
timestamp 1666464484
transform 1 0 33764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1666464484
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_369
timestamp 1666464484
transform 1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_381
timestamp 1666464484
transform 1 0 36156 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_387
timestamp 1666464484
transform 1 0 36708 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_393
timestamp 1666464484
transform 1 0 37260 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_404
timestamp 1666464484
transform 1 0 38272 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_417
timestamp 1666464484
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_425
timestamp 1666464484
transform 1 0 40204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_450
timestamp 1666464484
transform 1 0 42504 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1666464484
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_481
timestamp 1666464484
transform 1 0 45356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_493
timestamp 1666464484
transform 1 0 46460 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_505
timestamp 1666464484
transform 1 0 47564 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_517
timestamp 1666464484
transform 1 0 48668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_529
timestamp 1666464484
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1666464484
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_259
timestamp 1666464484
transform 1 0 24932 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1666464484
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1666464484
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_288
timestamp 1666464484
transform 1 0 27600 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_304
timestamp 1666464484
transform 1 0 29072 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_308
timestamp 1666464484
transform 1 0 29440 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1666464484
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_320
timestamp 1666464484
transform 1 0 30544 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_328
timestamp 1666464484
transform 1 0 31280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1666464484
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_349
timestamp 1666464484
transform 1 0 33212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_356
timestamp 1666464484
transform 1 0 33856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_362
timestamp 1666464484
transform 1 0 34408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_366
timestamp 1666464484
transform 1 0 34776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_376
timestamp 1666464484
transform 1 0 35696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1666464484
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_397
timestamp 1666464484
transform 1 0 37628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1666464484
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1666464484
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_426
timestamp 1666464484
transform 1 0 40296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_434
timestamp 1666464484
transform 1 0 41032 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1666464484
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_461
timestamp 1666464484
transform 1 0 43516 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_472
timestamp 1666464484
transform 1 0 44528 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_484
timestamp 1666464484
transform 1 0 45632 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_496
timestamp 1666464484
transform 1 0 46736 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1666464484
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_241
timestamp 1666464484
transform 1 0 23276 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_285
timestamp 1666464484
transform 1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_291
timestamp 1666464484
transform 1 0 27876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_299
timestamp 1666464484
transform 1 0 28612 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1666464484
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_322
timestamp 1666464484
transform 1 0 30728 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_328
timestamp 1666464484
transform 1 0 31280 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_336
timestamp 1666464484
transform 1 0 32016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_346
timestamp 1666464484
transform 1 0 32936 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_352
timestamp 1666464484
transform 1 0 33488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1666464484
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_372
timestamp 1666464484
transform 1 0 35328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_389
timestamp 1666464484
transform 1 0 36892 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_400
timestamp 1666464484
transform 1 0 37904 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_406
timestamp 1666464484
transform 1 0 38456 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1666464484
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_430
timestamp 1666464484
transform 1 0 40664 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_436
timestamp 1666464484
transform 1 0 41216 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666464484
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_487
timestamp 1666464484
transform 1 0 45908 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_493
timestamp 1666464484
transform 1 0 46460 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_505
timestamp 1666464484
transform 1 0 47564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_517
timestamp 1666464484
transform 1 0 48668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_529
timestamp 1666464484
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1666464484
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1666464484
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1666464484
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_291
timestamp 1666464484
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_295
timestamp 1666464484
transform 1 0 28244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_302
timestamp 1666464484
transform 1 0 28888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1666464484
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_322
timestamp 1666464484
transform 1 0 30728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_344
timestamp 1666464484
transform 1 0 32752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_356
timestamp 1666464484
transform 1 0 33856 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_368
timestamp 1666464484
transform 1 0 34960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_375
timestamp 1666464484
transform 1 0 35604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_383
timestamp 1666464484
transform 1 0 36340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_401
timestamp 1666464484
transform 1 0 37996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_421
timestamp 1666464484
transform 1 0 39836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_431
timestamp 1666464484
transform 1 0 40756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_444
timestamp 1666464484
transform 1 0 41952 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_461
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_470
timestamp 1666464484
transform 1 0 44344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_480
timestamp 1666464484
transform 1 0 45264 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_486
timestamp 1666464484
transform 1 0 45816 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1666464484
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1666464484
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_259
timestamp 1666464484
transform 1 0 24932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_267
timestamp 1666464484
transform 1 0 25668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_275
timestamp 1666464484
transform 1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1666464484
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_297
timestamp 1666464484
transform 1 0 28428 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_321
timestamp 1666464484
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_329
timestamp 1666464484
transform 1 0 31372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_343
timestamp 1666464484
transform 1 0 32660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_351
timestamp 1666464484
transform 1 0 33396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1666464484
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_394
timestamp 1666464484
transform 1 0 37352 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_408
timestamp 1666464484
transform 1 0 38640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1666464484
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_430
timestamp 1666464484
transform 1 0 40664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_441
timestamp 1666464484
transform 1 0 41676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_445
timestamp 1666464484
transform 1 0 42044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_451
timestamp 1666464484
transform 1 0 42596 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_466
timestamp 1666464484
transform 1 0 43976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_473
timestamp 1666464484
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_481
timestamp 1666464484
transform 1 0 45356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_493
timestamp 1666464484
transform 1 0 46460 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_505
timestamp 1666464484
transform 1 0 47564 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_517
timestamp 1666464484
transform 1 0 48668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_529
timestamp 1666464484
transform 1 0 49772 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1666464484
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1666464484
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1666464484
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_233
timestamp 1666464484
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_258
timestamp 1666464484
transform 1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1666464484
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_289
timestamp 1666464484
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_322
timestamp 1666464484
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1666464484
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_343
timestamp 1666464484
transform 1 0 32660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_353
timestamp 1666464484
transform 1 0 33580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_357
timestamp 1666464484
transform 1 0 33948 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_365
timestamp 1666464484
transform 1 0 34684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_374
timestamp 1666464484
transform 1 0 35512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_381
timestamp 1666464484
transform 1 0 36156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1666464484
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_399
timestamp 1666464484
transform 1 0 37812 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_405
timestamp 1666464484
transform 1 0 38364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_408
timestamp 1666464484
transform 1 0 38640 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_417
timestamp 1666464484
transform 1 0 39468 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_426
timestamp 1666464484
transform 1 0 40296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_434
timestamp 1666464484
transform 1 0 41032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_440
timestamp 1666464484
transform 1 0 41584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1666464484
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_459
timestamp 1666464484
transform 1 0 43332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_472
timestamp 1666464484
transform 1 0 44528 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_483
timestamp 1666464484
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1666464484
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1666464484
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_609
timestamp 1666464484
transform 1 0 57132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1666464484
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_623
timestamp 1666464484
transform 1 0 58420 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_258
timestamp 1666464484
transform 1 0 24840 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_264
timestamp 1666464484
transform 1 0 25392 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1666464484
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1666464484
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_282
timestamp 1666464484
transform 1 0 27048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_295
timestamp 1666464484
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_318
timestamp 1666464484
transform 1 0 30360 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_330
timestamp 1666464484
transform 1 0 31464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_338
timestamp 1666464484
transform 1 0 32200 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_344
timestamp 1666464484
transform 1 0 32752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_347
timestamp 1666464484
transform 1 0 33028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1666464484
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_381
timestamp 1666464484
transform 1 0 36156 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_387
timestamp 1666464484
transform 1 0 36708 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_396
timestamp 1666464484
transform 1 0 37536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_406
timestamp 1666464484
transform 1 0 38456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1666464484
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_428
timestamp 1666464484
transform 1 0 40480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_432
timestamp 1666464484
transform 1 0 40848 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_440
timestamp 1666464484
transform 1 0 41584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_446
timestamp 1666464484
transform 1 0 42136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_455
timestamp 1666464484
transform 1 0 42964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_464
timestamp 1666464484
transform 1 0 43792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1666464484
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_482
timestamp 1666464484
transform 1 0 45448 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666464484
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1666464484
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_256
timestamp 1666464484
transform 1 0 24656 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_262
timestamp 1666464484
transform 1 0 25208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1666464484
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_290
timestamp 1666464484
transform 1 0 27784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_298
timestamp 1666464484
transform 1 0 28520 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_304
timestamp 1666464484
transform 1 0 29072 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_321
timestamp 1666464484
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_325
timestamp 1666464484
transform 1 0 31004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_330
timestamp 1666464484
transform 1 0 31464 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_345
timestamp 1666464484
transform 1 0 32844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_352
timestamp 1666464484
transform 1 0 33488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_358
timestamp 1666464484
transform 1 0 34040 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_364
timestamp 1666464484
transform 1 0 34592 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_370
timestamp 1666464484
transform 1 0 35144 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_383
timestamp 1666464484
transform 1 0 36340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1666464484
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_401
timestamp 1666464484
transform 1 0 37996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_412
timestamp 1666464484
transform 1 0 39008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_425
timestamp 1666464484
transform 1 0 40204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_429
timestamp 1666464484
transform 1 0 40572 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_437
timestamp 1666464484
transform 1 0 41308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_445
timestamp 1666464484
transform 1 0 42044 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_460
timestamp 1666464484
transform 1 0 43424 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_467
timestamp 1666464484
transform 1 0 44068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_473
timestamp 1666464484
transform 1 0 44620 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_484
timestamp 1666464484
transform 1 0 45632 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_496
timestamp 1666464484
transform 1 0 46736 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1666464484
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1666464484
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1666464484
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1666464484
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_260
timestamp 1666464484
transform 1 0 25024 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_271
timestamp 1666464484
transform 1 0 26036 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_283
timestamp 1666464484
transform 1 0 27140 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_287
timestamp 1666464484
transform 1 0 27508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1666464484
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1666464484
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_321
timestamp 1666464484
transform 1 0 30636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_330
timestamp 1666464484
transform 1 0 31464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_339
timestamp 1666464484
transform 1 0 32292 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_353
timestamp 1666464484
transform 1 0 33580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1666464484
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_375
timestamp 1666464484
transform 1 0 35604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_386
timestamp 1666464484
transform 1 0 36616 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_400
timestamp 1666464484
transform 1 0 37904 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1666464484
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_409
timestamp 1666464484
transform 1 0 38732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1666464484
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_425
timestamp 1666464484
transform 1 0 40204 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_437
timestamp 1666464484
transform 1 0 41308 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_441
timestamp 1666464484
transform 1 0 41676 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_444
timestamp 1666464484
transform 1 0 41952 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_453
timestamp 1666464484
transform 1 0 42780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_465
timestamp 1666464484
transform 1 0 43884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1666464484
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_486
timestamp 1666464484
transform 1 0 45816 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_492
timestamp 1666464484
transform 1 0 46368 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_504
timestamp 1666464484
transform 1 0 47472 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_516
timestamp 1666464484
transform 1 0 48576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_528
timestamp 1666464484
transform 1 0 49680 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1666464484
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1666464484
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_254
timestamp 1666464484
transform 1 0 24472 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_260
timestamp 1666464484
transform 1 0 25024 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_268
timestamp 1666464484
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_286
timestamp 1666464484
transform 1 0 27416 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_294
timestamp 1666464484
transform 1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_302
timestamp 1666464484
transform 1 0 28888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_313
timestamp 1666464484
transform 1 0 29900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_320
timestamp 1666464484
transform 1 0 30544 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_328
timestamp 1666464484
transform 1 0 31280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1666464484
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1666464484
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_353
timestamp 1666464484
transform 1 0 33580 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_366
timestamp 1666464484
transform 1 0 34776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_377
timestamp 1666464484
transform 1 0 35788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1666464484
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_403
timestamp 1666464484
transform 1 0 38180 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_409
timestamp 1666464484
transform 1 0 38732 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_418
timestamp 1666464484
transform 1 0 39560 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_426
timestamp 1666464484
transform 1 0 40296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_430
timestamp 1666464484
transform 1 0 40664 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_440
timestamp 1666464484
transform 1 0 41584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1666464484
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_455
timestamp 1666464484
transform 1 0 42964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_459
timestamp 1666464484
transform 1 0 43332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_471
timestamp 1666464484
transform 1 0 44436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_477
timestamp 1666464484
transform 1 0 44988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_484
timestamp 1666464484
transform 1 0 45632 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_490
timestamp 1666464484
transform 1 0 46184 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1666464484
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1666464484
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1666464484
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1666464484
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_261
timestamp 1666464484
transform 1 0 25116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1666464484
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_280
timestamp 1666464484
transform 1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_291
timestamp 1666464484
transform 1 0 27876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1666464484
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_323
timestamp 1666464484
transform 1 0 30820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1666464484
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_344
timestamp 1666464484
transform 1 0 32752 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_356
timestamp 1666464484
transform 1 0 33856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1666464484
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_371
timestamp 1666464484
transform 1 0 35236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_374
timestamp 1666464484
transform 1 0 35512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_382
timestamp 1666464484
transform 1 0 36248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_388
timestamp 1666464484
transform 1 0 36800 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_392
timestamp 1666464484
transform 1 0 37168 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_396
timestamp 1666464484
transform 1 0 37536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1666464484
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_407
timestamp 1666464484
transform 1 0 38548 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1666464484
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_430
timestamp 1666464484
transform 1 0 40664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_436
timestamp 1666464484
transform 1 0 41216 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_453
timestamp 1666464484
transform 1 0 42780 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_465
timestamp 1666464484
transform 1 0 43884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1666464484
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_486
timestamp 1666464484
transform 1 0 45816 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_492
timestamp 1666464484
transform 1 0 46368 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_504
timestamp 1666464484
transform 1 0 47472 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_516
timestamp 1666464484
transform 1 0 48576 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_528
timestamp 1666464484
transform 1 0 49680 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1666464484
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1666464484
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_246
timestamp 1666464484
transform 1 0 23736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1666464484
transform 1 0 24472 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1666464484
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1666464484
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_290
timestamp 1666464484
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_298
timestamp 1666464484
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_304
timestamp 1666464484
transform 1 0 29072 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_312
timestamp 1666464484
transform 1 0 29808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_319
timestamp 1666464484
transform 1 0 30452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_325
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1666464484
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_347
timestamp 1666464484
transform 1 0 33028 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_353
timestamp 1666464484
transform 1 0 33580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1666464484
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_364
timestamp 1666464484
transform 1 0 34592 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_369
timestamp 1666464484
transform 1 0 35052 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_379
timestamp 1666464484
transform 1 0 35972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_386
timestamp 1666464484
transform 1 0 36616 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_399
timestamp 1666464484
transform 1 0 37812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_405
timestamp 1666464484
transform 1 0 38364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_412
timestamp 1666464484
transform 1 0 39008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_419
timestamp 1666464484
transform 1 0 39652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_423
timestamp 1666464484
transform 1 0 40020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_429
timestamp 1666464484
transform 1 0 40572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_436
timestamp 1666464484
transform 1 0 41216 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_445
timestamp 1666464484
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_456
timestamp 1666464484
transform 1 0 43056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_460
timestamp 1666464484
transform 1 0 43424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_466
timestamp 1666464484
transform 1 0 43976 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_475
timestamp 1666464484
transform 1 0 44804 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_486
timestamp 1666464484
transform 1 0 45816 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_498
timestamp 1666464484
transform 1 0 46920 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1666464484
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1666464484
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1666464484
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_241
timestamp 1666464484
transform 1 0 23276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1666464484
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_264
timestamp 1666464484
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_272
timestamp 1666464484
transform 1 0 26128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_280
timestamp 1666464484
transform 1 0 26864 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1666464484
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_294
timestamp 1666464484
transform 1 0 28152 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_318
timestamp 1666464484
transform 1 0 30360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_330
timestamp 1666464484
transform 1 0 31464 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1666464484
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_343
timestamp 1666464484
transform 1 0 32660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_349
timestamp 1666464484
transform 1 0 33212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666464484
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666464484
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_373
timestamp 1666464484
transform 1 0 35420 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_379
timestamp 1666464484
transform 1 0 35972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_391
timestamp 1666464484
transform 1 0 37076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_397
timestamp 1666464484
transform 1 0 37628 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_406
timestamp 1666464484
transform 1 0 38456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1666464484
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_429
timestamp 1666464484
transform 1 0 40572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_435
timestamp 1666464484
transform 1 0 41124 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_445
timestamp 1666464484
transform 1 0 42044 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_457
timestamp 1666464484
transform 1 0 43148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_466
timestamp 1666464484
transform 1 0 43976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_472
timestamp 1666464484
transform 1 0 44528 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_486
timestamp 1666464484
transform 1 0 45816 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_492
timestamp 1666464484
transform 1 0 46368 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_504
timestamp 1666464484
transform 1 0 47472 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_516
timestamp 1666464484
transform 1 0 48576 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_528
timestamp 1666464484
transform 1 0 49680 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1666464484
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1666464484
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1666464484
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1666464484
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_250
timestamp 1666464484
transform 1 0 24104 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_262
timestamp 1666464484
transform 1 0 25208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_289
timestamp 1666464484
transform 1 0 27692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1666464484
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1666464484
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_321
timestamp 1666464484
transform 1 0 30636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1666464484
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_343
timestamp 1666464484
transform 1 0 32660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1666464484
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_362
timestamp 1666464484
transform 1 0 34408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_369
timestamp 1666464484
transform 1 0 35052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_373
timestamp 1666464484
transform 1 0 35420 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_377
timestamp 1666464484
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_399
timestamp 1666464484
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_410
timestamp 1666464484
transform 1 0 38824 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_423
timestamp 1666464484
transform 1 0 40020 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_436
timestamp 1666464484
transform 1 0 41216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1666464484
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_457
timestamp 1666464484
transform 1 0 43148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_466
timestamp 1666464484
transform 1 0 43976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_472
timestamp 1666464484
transform 1 0 44528 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_481
timestamp 1666464484
transform 1 0 45356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_489
timestamp 1666464484
transform 1 0 46092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666464484
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1666464484
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_217
timestamp 1666464484
transform 1 0 21068 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_239
timestamp 1666464484
transform 1 0 23092 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1666464484
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_262
timestamp 1666464484
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1666464484
transform 1 0 26036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_275
timestamp 1666464484
transform 1 0 26404 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_283
timestamp 1666464484
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_295
timestamp 1666464484
transform 1 0 28244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666464484
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_317
timestamp 1666464484
transform 1 0 30268 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1666464484
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_335
timestamp 1666464484
transform 1 0 31924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_350
timestamp 1666464484
transform 1 0 33304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1666464484
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_371
timestamp 1666464484
transform 1 0 35236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_375
timestamp 1666464484
transform 1 0 35604 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_382
timestamp 1666464484
transform 1 0 36248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_388
timestamp 1666464484
transform 1 0 36800 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_399
timestamp 1666464484
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_410
timestamp 1666464484
transform 1 0 38824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1666464484
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_426
timestamp 1666464484
transform 1 0 40296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1666464484
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_438
timestamp 1666464484
transform 1 0 41400 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_450
timestamp 1666464484
transform 1 0 42504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_461
timestamp 1666464484
transform 1 0 43516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_470
timestamp 1666464484
transform 1 0 44344 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_487
timestamp 1666464484
transform 1 0 45908 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_499
timestamp 1666464484
transform 1 0 47012 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_511
timestamp 1666464484
transform 1 0 48116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_523
timestamp 1666464484
transform 1 0 49220 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1666464484
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_233
timestamp 1666464484
transform 1 0 22540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1666464484
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_299
timestamp 1666464484
transform 1 0 28612 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1666464484
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1666464484
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1666464484
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_346
timestamp 1666464484
transform 1 0 32936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 1666464484
transform 1 0 33488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_364
timestamp 1666464484
transform 1 0 34592 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_372
timestamp 1666464484
transform 1 0 35328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_384
timestamp 1666464484
transform 1 0 36432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1666464484
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_397
timestamp 1666464484
transform 1 0 37628 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_406
timestamp 1666464484
transform 1 0 38456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_418
timestamp 1666464484
transform 1 0 39560 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_429
timestamp 1666464484
transform 1 0 40572 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_438
timestamp 1666464484
transform 1 0 41400 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1666464484
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_457
timestamp 1666464484
transform 1 0 43148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_467
timestamp 1666464484
transform 1 0 44068 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_484
timestamp 1666464484
transform 1 0 45632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_494
timestamp 1666464484
transform 1 0 46552 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1666464484
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1666464484
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1666464484
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_609
timestamp 1666464484
transform 1 0 57132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_614
timestamp 1666464484
transform 1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1666464484
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_232
timestamp 1666464484
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1666464484
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1666464484
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_276
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_284
timestamp 1666464484
transform 1 0 27232 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_297
timestamp 1666464484
transform 1 0 28428 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_300
timestamp 1666464484
transform 1 0 28704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1666464484
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_328
timestamp 1666464484
transform 1 0 31280 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_345
timestamp 1666464484
transform 1 0 32844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_352
timestamp 1666464484
transform 1 0 33488 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_358
timestamp 1666464484
transform 1 0 34040 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1666464484
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_370
timestamp 1666464484
transform 1 0 35144 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_381
timestamp 1666464484
transform 1 0 36156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_388
timestamp 1666464484
transform 1 0 36800 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_394
timestamp 1666464484
transform 1 0 37352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_401
timestamp 1666464484
transform 1 0 37996 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1666464484
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_431
timestamp 1666464484
transform 1 0 40756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_435
timestamp 1666464484
transform 1 0 41124 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_439
timestamp 1666464484
transform 1 0 41492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_448
timestamp 1666464484
transform 1 0 42320 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_454
timestamp 1666464484
transform 1 0 42872 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_458
timestamp 1666464484
transform 1 0 43240 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_465
timestamp 1666464484
transform 1 0 43884 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_471
timestamp 1666464484
transform 1 0 44436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666464484
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_485
timestamp 1666464484
transform 1 0 45724 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_491
timestamp 1666464484
transform 1 0 46276 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_503
timestamp 1666464484
transform 1 0 47380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_515
timestamp 1666464484
transform 1 0 48484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_527
timestamp 1666464484
transform 1 0 49588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1666464484
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1666464484
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1666464484
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1666464484
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_9
timestamp 1666464484
transform 1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1666464484
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_266
timestamp 1666464484
transform 1 0 25576 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1666464484
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_289
timestamp 1666464484
transform 1 0 27692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_298
timestamp 1666464484
transform 1 0 28520 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_307
timestamp 1666464484
transform 1 0 29348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_321
timestamp 1666464484
transform 1 0 30636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1666464484
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_358
timestamp 1666464484
transform 1 0 34040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_368
timestamp 1666464484
transform 1 0 34960 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_376
timestamp 1666464484
transform 1 0 35696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_382
timestamp 1666464484
transform 1 0 36248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1666464484
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1666464484
transform 1 0 38088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1666464484
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_413
timestamp 1666464484
transform 1 0 39100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_421
timestamp 1666464484
transform 1 0 39836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_436
timestamp 1666464484
transform 1 0 41216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1666464484
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_461
timestamp 1666464484
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_481
timestamp 1666464484
transform 1 0 45356 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_487
timestamp 1666464484
transform 1 0 45908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_499
timestamp 1666464484
transform 1 0 47012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666464484
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1666464484
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1666464484
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1666464484
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1666464484
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1666464484
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1666464484
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1666464484
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_322
timestamp 1666464484
transform 1 0 30728 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_351
timestamp 1666464484
transform 1 0 33396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_357
timestamp 1666464484
transform 1 0 33948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1666464484
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_371
timestamp 1666464484
transform 1 0 35236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_378
timestamp 1666464484
transform 1 0 35880 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_396
timestamp 1666464484
transform 1 0 37536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_402
timestamp 1666464484
transform 1 0 38088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_412
timestamp 1666464484
transform 1 0 39008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1666464484
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_432
timestamp 1666464484
transform 1 0 40848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_444
timestamp 1666464484
transform 1 0 41952 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_455
timestamp 1666464484
transform 1 0 42964 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_467
timestamp 1666464484
transform 1 0 44068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1666464484
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_485
timestamp 1666464484
transform 1 0 45724 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_495
timestamp 1666464484
transform 1 0 46644 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_507
timestamp 1666464484
transform 1 0 47748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_519
timestamp 1666464484
transform 1 0 48852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1666464484
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1666464484
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1666464484
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1666464484
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_264
timestamp 1666464484
transform 1 0 25392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1666464484
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_296
timestamp 1666464484
transform 1 0 28336 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_308
timestamp 1666464484
transform 1 0 29440 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_320
timestamp 1666464484
transform 1 0 30544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_324
timestamp 1666464484
transform 1 0 30912 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_327
timestamp 1666464484
transform 1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1666464484
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_343
timestamp 1666464484
transform 1 0 32660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_346
timestamp 1666464484
transform 1 0 32936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_352
timestamp 1666464484
transform 1 0 33488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_364
timestamp 1666464484
transform 1 0 34592 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_370
timestamp 1666464484
transform 1 0 35144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_378
timestamp 1666464484
transform 1 0 35880 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1666464484
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_397
timestamp 1666464484
transform 1 0 37628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_415
timestamp 1666464484
transform 1 0 39284 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_425
timestamp 1666464484
transform 1 0 40204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_429
timestamp 1666464484
transform 1 0 40572 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_439
timestamp 1666464484
transform 1 0 41492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1666464484
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_458
timestamp 1666464484
transform 1 0 43240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_462
timestamp 1666464484
transform 1 0 43608 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_469
timestamp 1666464484
transform 1 0 44252 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_483
timestamp 1666464484
transform 1 0 45540 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_489
timestamp 1666464484
transform 1 0 46092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_501
timestamp 1666464484
transform 1 0 47196 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1666464484
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1666464484
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1666464484
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_282
timestamp 1666464484
transform 1 0 27048 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_288
timestamp 1666464484
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1666464484
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_317
timestamp 1666464484
transform 1 0 30268 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1666464484
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_352
timestamp 1666464484
transform 1 0 33488 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1666464484
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_374
timestamp 1666464484
transform 1 0 35512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_398
timestamp 1666464484
transform 1 0 37720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_404
timestamp 1666464484
transform 1 0 38272 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1666464484
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_428
timestamp 1666464484
transform 1 0 40480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_436
timestamp 1666464484
transform 1 0 41216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_442
timestamp 1666464484
transform 1 0 41768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_454
timestamp 1666464484
transform 1 0 42872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_460
timestamp 1666464484
transform 1 0 43424 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_472
timestamp 1666464484
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_485
timestamp 1666464484
transform 1 0 45724 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_497
timestamp 1666464484
transform 1 0 46828 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_509
timestamp 1666464484
transform 1 0 47932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_521
timestamp 1666464484
transform 1 0 49036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_529
timestamp 1666464484
transform 1 0 49772 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1666464484
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1666464484
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1666464484
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_252
timestamp 1666464484
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_264
timestamp 1666464484
transform 1 0 25392 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_270
timestamp 1666464484
transform 1 0 25944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1666464484
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1666464484
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_292
timestamp 1666464484
transform 1 0 27968 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1666464484
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1666464484
transform 1 0 28796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_325
timestamp 1666464484
transform 1 0 31004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1666464484
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_345
timestamp 1666464484
transform 1 0 32844 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_356
timestamp 1666464484
transform 1 0 33856 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_363
timestamp 1666464484
transform 1 0 34500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_369
timestamp 1666464484
transform 1 0 35052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_377
timestamp 1666464484
transform 1 0 35788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_384
timestamp 1666464484
transform 1 0 36432 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1666464484
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_413
timestamp 1666464484
transform 1 0 39100 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_425
timestamp 1666464484
transform 1 0 40204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_429
timestamp 1666464484
transform 1 0 40572 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_439
timestamp 1666464484
transform 1 0 41492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1666464484
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_499
timestamp 1666464484
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1666464484
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1666464484
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_241
timestamp 1666464484
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1666464484
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_278
timestamp 1666464484
transform 1 0 26680 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1666464484
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1666464484
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_320
timestamp 1666464484
transform 1 0 30544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_330
timestamp 1666464484
transform 1 0 31464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_336
timestamp 1666464484
transform 1 0 32016 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_342
timestamp 1666464484
transform 1 0 32568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_353
timestamp 1666464484
transform 1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1666464484
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_372
timestamp 1666464484
transform 1 0 35328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_376
timestamp 1666464484
transform 1 0 35696 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_400
timestamp 1666464484
transform 1 0 37904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_410
timestamp 1666464484
transform 1 0 38824 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1666464484
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_425
timestamp 1666464484
transform 1 0 40204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_431
timestamp 1666464484
transform 1 0 40756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_437
timestamp 1666464484
transform 1 0 41308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_451
timestamp 1666464484
transform 1 0 42596 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_461
timestamp 1666464484
transform 1 0 43516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_473
timestamp 1666464484
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1666464484
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_251
timestamp 1666464484
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_257
timestamp 1666464484
transform 1 0 24748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1666464484
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1666464484
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_303
timestamp 1666464484
transform 1 0 28980 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_311
timestamp 1666464484
transform 1 0 29716 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1666464484
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_348
timestamp 1666464484
transform 1 0 33120 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_359
timestamp 1666464484
transform 1 0 34132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_383
timestamp 1666464484
transform 1 0 36340 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1666464484
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_397
timestamp 1666464484
transform 1 0 37628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_407
timestamp 1666464484
transform 1 0 38548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_413
timestamp 1666464484
transform 1 0 39100 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_419
timestamp 1666464484
transform 1 0 39652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_431
timestamp 1666464484
transform 1 0 40756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1666464484
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_455
timestamp 1666464484
transform 1 0 42964 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_467
timestamp 1666464484
transform 1 0 44068 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_479
timestamp 1666464484
transform 1 0 45172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_491
timestamp 1666464484
transform 1 0 46276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1666464484
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1666464484
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1666464484
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_217
timestamp 1666464484
transform 1 0 21068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1666464484
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1666464484
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_238
timestamp 1666464484
transform 1 0 23000 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1666464484
transform 1 0 23276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1666464484
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_268
timestamp 1666464484
transform 1 0 25760 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_276
timestamp 1666464484
transform 1 0 26496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1666464484
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1666464484
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_298
timestamp 1666464484
transform 1 0 28520 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1666464484
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_317
timestamp 1666464484
transform 1 0 30268 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_324
timestamp 1666464484
transform 1 0 30912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_331
timestamp 1666464484
transform 1 0 31556 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_339
timestamp 1666464484
transform 1 0 32292 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_344
timestamp 1666464484
transform 1 0 32752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_350
timestamp 1666464484
transform 1 0 33304 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_358
timestamp 1666464484
transform 1 0 34040 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1666464484
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_372
timestamp 1666464484
transform 1 0 35328 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_407
timestamp 1666464484
transform 1 0 38548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666464484
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_201
timestamp 1666464484
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1666464484
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1666464484
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_244
timestamp 1666464484
transform 1 0 23552 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_252
timestamp 1666464484
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1666464484
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1666464484
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1666464484
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1666464484
transform 1 0 29256 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1666464484
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_362
timestamp 1666464484
transform 1 0 34408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_374
timestamp 1666464484
transform 1 0 35512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_380
timestamp 1666464484
transform 1 0 36064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1666464484
transform 1 0 36616 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666464484
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1666464484
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1666464484
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1666464484
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_177
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_185
timestamp 1666464484
transform 1 0 18124 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1666464484
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_217
timestamp 1666464484
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_229
timestamp 1666464484
transform 1 0 22172 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1666464484
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_267
timestamp 1666464484
transform 1 0 25668 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_275
timestamp 1666464484
transform 1 0 26404 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_283
timestamp 1666464484
transform 1 0 27140 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_287
timestamp 1666464484
transform 1 0 27508 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1666464484
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_297
timestamp 1666464484
transform 1 0 28428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1666464484
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_326
timestamp 1666464484
transform 1 0 31096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_334
timestamp 1666464484
transform 1 0 31832 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1666464484
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_394
timestamp 1666464484
transform 1 0 37352 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_406
timestamp 1666464484
transform 1 0 38456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1666464484
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666464484
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1666464484
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_9
timestamp 1666464484
transform 1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1666464484
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_189
timestamp 1666464484
transform 1 0 18492 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_195
timestamp 1666464484
transform 1 0 19044 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1666464484
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_208
timestamp 1666464484
transform 1 0 20240 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1666464484
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_243
timestamp 1666464484
transform 1 0 23460 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_247
timestamp 1666464484
transform 1 0 23828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1666464484
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_264
timestamp 1666464484
transform 1 0 25392 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_272
timestamp 1666464484
transform 1 0 26128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_288
timestamp 1666464484
transform 1 0 27600 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_299
timestamp 1666464484
transform 1 0 28612 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_309
timestamp 1666464484
transform 1 0 29532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1666464484
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1666464484
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_346
timestamp 1666464484
transform 1 0 32936 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 33672 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_378
timestamp 1666464484
transform 1 0 35880 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1666464484
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1666464484
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1666464484
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_609
timestamp 1666464484
transform 1 0 57132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_614
timestamp 1666464484
transform 1 0 57592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1666464484
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_206
timestamp 1666464484
transform 1 0 20056 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1666464484
transform 1 0 20884 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_219
timestamp 1666464484
transform 1 0 21252 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_227
timestamp 1666464484
transform 1 0 21988 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_234
timestamp 1666464484
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_246
timestamp 1666464484
transform 1 0 23736 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1666464484
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_262
timestamp 1666464484
transform 1 0 25208 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_273
timestamp 1666464484
transform 1 0 26220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_297
timestamp 1666464484
transform 1 0 28428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_324
timestamp 1666464484
transform 1 0 30912 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_330
timestamp 1666464484
transform 1 0 31464 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_336
timestamp 1666464484
transform 1 0 32016 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_339
timestamp 1666464484
transform 1 0 32292 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_347
timestamp 1666464484
transform 1 0 33028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_355
timestamp 1666464484
transform 1 0 33764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 1666464484
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666464484
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1666464484
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1666464484
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_191
timestamp 1666464484
transform 1 0 18676 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_199
timestamp 1666464484
transform 1 0 19412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1666464484
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_211
timestamp 1666464484
transform 1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1666464484
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_238
timestamp 1666464484
transform 1 0 23000 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_250
timestamp 1666464484
transform 1 0 24104 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1666464484
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1666464484
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1666464484
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1666464484
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_321
timestamp 1666464484
transform 1 0 30636 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1666464484
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_343
timestamp 1666464484
transform 1 0 32660 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_350
timestamp 1666464484
transform 1 0 33304 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_356
timestamp 1666464484
transform 1 0 33856 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_362
timestamp 1666464484
transform 1 0 34408 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_369
timestamp 1666464484
transform 1 0 35052 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_375
timestamp 1666464484
transform 1 0 35604 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_382
timestamp 1666464484
transform 1 0 36248 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1666464484
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666464484
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1666464484
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 1666464484
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_214
timestamp 1666464484
transform 1 0 20792 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_220
timestamp 1666464484
transform 1 0 21344 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_224
timestamp 1666464484
transform 1 0 21712 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_229
timestamp 1666464484
transform 1 0 22172 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_236
timestamp 1666464484
transform 1 0 22816 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_244
timestamp 1666464484
transform 1 0 23552 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1666464484
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_259
timestamp 1666464484
transform 1 0 24932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1666464484
transform 1 0 26036 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_278
timestamp 1666464484
transform 1 0 26680 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1666464484
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_298
timestamp 1666464484
transform 1 0 28520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1666464484
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_317
timestamp 1666464484
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_325
timestamp 1666464484
transform 1 0 31004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_332
timestamp 1666464484
transform 1 0 31648 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_340
timestamp 1666464484
transform 1 0 32384 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_348
timestamp 1666464484
transform 1 0 33120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1666464484
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_370
timestamp 1666464484
transform 1 0 35144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_374
timestamp 1666464484
transform 1 0 35512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_382
timestamp 1666464484
transform 1 0 36248 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_388
timestamp 1666464484
transform 1 0 36800 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_402
timestamp 1666464484
transform 1 0 38088 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_414
timestamp 1666464484
transform 1 0 39192 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_153
timestamp 1666464484
transform 1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1666464484
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_177
timestamp 1666464484
transform 1 0 17388 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_187
timestamp 1666464484
transform 1 0 18308 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_199
timestamp 1666464484
transform 1 0 19412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1666464484
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_233
timestamp 1666464484
transform 1 0 22540 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_245
timestamp 1666464484
transform 1 0 23644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_259
timestamp 1666464484
transform 1 0 24932 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1666464484
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1666464484
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1666464484
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_328
timestamp 1666464484
transform 1 0 31280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_344
timestamp 1666464484
transform 1 0 32752 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_353
timestamp 1666464484
transform 1 0 33580 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_364
timestamp 1666464484
transform 1 0 34592 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_375
timestamp 1666464484
transform 1 0 35604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_383
timestamp 1666464484
transform 1 0 36340 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1666464484
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666464484
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_176
timestamp 1666464484
transform 1 0 17296 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp 1666464484
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_203
timestamp 1666464484
transform 1 0 19780 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_211
timestamp 1666464484
transform 1 0 20516 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1666464484
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_228
timestamp 1666464484
transform 1 0 22080 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_241
timestamp 1666464484
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1666464484
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1666464484
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_268
timestamp 1666464484
transform 1 0 25760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp 1666464484
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_282
timestamp 1666464484
transform 1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_292
timestamp 1666464484
transform 1 0 27968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_298
timestamp 1666464484
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1666464484
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_317
timestamp 1666464484
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_322
timestamp 1666464484
transform 1 0 30728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_344
timestamp 1666464484
transform 1 0 32752 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1666464484
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_369
timestamp 1666464484
transform 1 0 35052 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_376
timestamp 1666464484
transform 1 0 35696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_385
timestamp 1666464484
transform 1 0 36524 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_398
timestamp 1666464484
transform 1 0 37720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_410
timestamp 1666464484
transform 1 0 38824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1666464484
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666464484
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1666464484
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_191
timestamp 1666464484
transform 1 0 18676 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_206
timestamp 1666464484
transform 1 0 20056 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_213
timestamp 1666464484
transform 1 0 20700 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_219
timestamp 1666464484
transform 1 0 21252 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1666464484
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_247
timestamp 1666464484
transform 1 0 23828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_260
timestamp 1666464484
transform 1 0 25024 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_288
timestamp 1666464484
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_294
timestamp 1666464484
transform 1 0 28152 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_300
timestamp 1666464484
transform 1 0 28704 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_304
timestamp 1666464484
transform 1 0 29072 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_310
timestamp 1666464484
transform 1 0 29624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_314
timestamp 1666464484
transform 1 0 29992 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_324
timestamp 1666464484
transform 1 0 30912 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1666464484
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_343
timestamp 1666464484
transform 1 0 32660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_348
timestamp 1666464484
transform 1 0 33120 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_362
timestamp 1666464484
transform 1 0 34408 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_376
timestamp 1666464484
transform 1 0 35696 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_384
timestamp 1666464484
transform 1 0 36432 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_401
timestamp 1666464484
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_412
timestamp 1666464484
transform 1 0 39008 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_419
timestamp 1666464484
transform 1 0 39652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_431
timestamp 1666464484
transform 1 0 40756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_443
timestamp 1666464484
transform 1 0 41860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666464484
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp 1666464484
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_164
timestamp 1666464484
transform 1 0 16192 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1666464484
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_205
timestamp 1666464484
transform 1 0 19964 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1666464484
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_220
timestamp 1666464484
transform 1 0 21344 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_230
timestamp 1666464484
transform 1 0 22264 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_242
timestamp 1666464484
transform 1 0 23368 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1666464484
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_261
timestamp 1666464484
transform 1 0 25116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_269
timestamp 1666464484
transform 1 0 25852 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_278
timestamp 1666464484
transform 1 0 26680 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_291
timestamp 1666464484
transform 1 0 27876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1666464484
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_314
timestamp 1666464484
transform 1 0 29992 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_326
timestamp 1666464484
transform 1 0 31096 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_330
timestamp 1666464484
transform 1 0 31464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_340
timestamp 1666464484
transform 1 0 32384 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_348
timestamp 1666464484
transform 1 0 33120 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1666464484
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1666464484
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_369
timestamp 1666464484
transform 1 0 35052 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_380
timestamp 1666464484
transform 1 0 36064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_384
timestamp 1666464484
transform 1 0 36432 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_391
timestamp 1666464484
transform 1 0 37076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_400
timestamp 1666464484
transform 1 0 37904 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_428
timestamp 1666464484
transform 1 0 40480 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_440
timestamp 1666464484
transform 1 0 41584 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_452
timestamp 1666464484
transform 1 0 42688 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_464
timestamp 1666464484
transform 1 0 43792 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_156
timestamp 1666464484
transform 1 0 15456 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1666464484
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_177
timestamp 1666464484
transform 1 0 17388 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_186
timestamp 1666464484
transform 1 0 18216 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_211
timestamp 1666464484
transform 1 0 20516 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1666464484
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1666464484
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_242
timestamp 1666464484
transform 1 0 23368 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_250
timestamp 1666464484
transform 1 0 24104 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1666464484
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1666464484
transform 1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1666464484
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1666464484
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_287
timestamp 1666464484
transform 1 0 27508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_296
timestamp 1666464484
transform 1 0 28336 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_306
timestamp 1666464484
transform 1 0 29256 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_314
timestamp 1666464484
transform 1 0 29992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_320
timestamp 1666464484
transform 1 0 30544 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_324
timestamp 1666464484
transform 1 0 30912 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_328
timestamp 1666464484
transform 1 0 31280 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1666464484
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_347
timestamp 1666464484
transform 1 0 33028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_356
timestamp 1666464484
transform 1 0 33856 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_362
timestamp 1666464484
transform 1 0 34408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_368
timestamp 1666464484
transform 1 0 34960 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_374
timestamp 1666464484
transform 1 0 35512 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_378
timestamp 1666464484
transform 1 0 35880 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1666464484
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_400
timestamp 1666464484
transform 1 0 37904 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_410
timestamp 1666464484
transform 1 0 38824 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_431
timestamp 1666464484
transform 1 0 40756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_443
timestamp 1666464484
transform 1 0 41860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1666464484
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_149
timestamp 1666464484
transform 1 0 14812 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_159
timestamp 1666464484
transform 1 0 15732 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_171
timestamp 1666464484
transform 1 0 16836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_181
timestamp 1666464484
transform 1 0 17756 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1666464484
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1666464484
transform 1 0 20424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_220
timestamp 1666464484
transform 1 0 21344 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_231
timestamp 1666464484
transform 1 0 22356 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1666464484
transform 1 0 22908 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_241
timestamp 1666464484
transform 1 0 23276 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1666464484
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_263
timestamp 1666464484
transform 1 0 25300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_267
timestamp 1666464484
transform 1 0 25668 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_276
timestamp 1666464484
transform 1 0 26496 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_284
timestamp 1666464484
transform 1 0 27232 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_292
timestamp 1666464484
transform 1 0 27968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_296
timestamp 1666464484
transform 1 0 28336 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1666464484
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_322
timestamp 1666464484
transform 1 0 30728 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_339
timestamp 1666464484
transform 1 0 32292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_344
timestamp 1666464484
transform 1 0 32752 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_356
timestamp 1666464484
transform 1 0 33856 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1666464484
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_374
timestamp 1666464484
transform 1 0 35512 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_383
timestamp 1666464484
transform 1 0 36340 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_395
timestamp 1666464484
transform 1 0 37444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_407
timestamp 1666464484
transform 1 0 38548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_412
timestamp 1666464484
transform 1 0 39008 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1666464484
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1666464484
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_185
timestamp 1666464484
transform 1 0 18124 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1666464484
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1666464484
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_201
timestamp 1666464484
transform 1 0 19596 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_204
timestamp 1666464484
transform 1 0 19872 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_210
timestamp 1666464484
transform 1 0 20424 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1666464484
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 1666464484
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_238
timestamp 1666464484
transform 1 0 23000 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_247
timestamp 1666464484
transform 1 0 23828 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_255
timestamp 1666464484
transform 1 0 24564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_260
timestamp 1666464484
transform 1 0 25024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_264
timestamp 1666464484
transform 1 0 25392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_269
timestamp 1666464484
transform 1 0 25852 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_275
timestamp 1666464484
transform 1 0 26404 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1666464484
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_285
timestamp 1666464484
transform 1 0 27324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_296
timestamp 1666464484
transform 1 0 28336 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_306
timestamp 1666464484
transform 1 0 29256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_315
timestamp 1666464484
transform 1 0 30084 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_328
timestamp 1666464484
transform 1 0 31280 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1666464484
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_342
timestamp 1666464484
transform 1 0 32568 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_348
timestamp 1666464484
transform 1 0 33120 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_359
timestamp 1666464484
transform 1 0 34132 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_365
timestamp 1666464484
transform 1 0 34684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_377
timestamp 1666464484
transform 1 0 35788 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1666464484
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_402
timestamp 1666464484
transform 1 0 38088 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_414
timestamp 1666464484
transform 1 0 39192 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_426
timestamp 1666464484
transform 1 0 40296 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_438
timestamp 1666464484
transform 1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1666464484
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1666464484
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_614
timestamp 1666464484
transform 1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1666464484
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_9
timestamp 1666464484
transform 1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1666464484
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_151
timestamp 1666464484
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_163
timestamp 1666464484
transform 1 0 16100 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_176
timestamp 1666464484
transform 1 0 17296 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1666464484
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_202
timestamp 1666464484
transform 1 0 19688 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_210
timestamp 1666464484
transform 1 0 20424 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_219
timestamp 1666464484
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_225
timestamp 1666464484
transform 1 0 21804 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_231
timestamp 1666464484
transform 1 0 22356 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_239
timestamp 1666464484
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_261
timestamp 1666464484
transform 1 0 25116 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_267
timestamp 1666464484
transform 1 0 25668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_278
timestamp 1666464484
transform 1 0 26680 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_286
timestamp 1666464484
transform 1 0 27416 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_292
timestamp 1666464484
transform 1 0 27968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_302
timestamp 1666464484
transform 1 0 28888 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1666464484
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_324
timestamp 1666464484
transform 1 0 30912 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_328
timestamp 1666464484
transform 1 0 31280 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_338
timestamp 1666464484
transform 1 0 32200 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_353
timestamp 1666464484
transform 1 0 33580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1666464484
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_381
timestamp 1666464484
transform 1 0 36156 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_387
timestamp 1666464484
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_399
timestamp 1666464484
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_411
timestamp 1666464484
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666464484
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_144
timestamp 1666464484
transform 1 0 14352 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_152
timestamp 1666464484
transform 1 0 15088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_156
timestamp 1666464484
transform 1 0 15456 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1666464484
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_178
timestamp 1666464484
transform 1 0 17480 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_186
timestamp 1666464484
transform 1 0 18216 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_191
timestamp 1666464484
transform 1 0 18676 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_202
timestamp 1666464484
transform 1 0 19688 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_206
timestamp 1666464484
transform 1 0 20056 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_213
timestamp 1666464484
transform 1 0 20700 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_219
timestamp 1666464484
transform 1 0 21252 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1666464484
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1666464484
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1666464484
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_256
timestamp 1666464484
transform 1 0 24656 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_267
timestamp 1666464484
transform 1 0 25668 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1666464484
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_288
timestamp 1666464484
transform 1 0 27600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_295
timestamp 1666464484
transform 1 0 28244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_299
timestamp 1666464484
transform 1 0 28612 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_316
timestamp 1666464484
transform 1 0 30176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_327
timestamp 1666464484
transform 1 0 31188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_331
timestamp 1666464484
transform 1 0 31556 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1666464484
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_344
timestamp 1666464484
transform 1 0 32752 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_352
timestamp 1666464484
transform 1 0 33488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_356
timestamp 1666464484
transform 1 0 33856 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1666464484
transform 1 0 34408 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1666464484
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666464484
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1666464484
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1666464484
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1666464484
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_173
timestamp 1666464484
transform 1 0 17020 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_181
timestamp 1666464484
transform 1 0 17756 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1666464484
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_202
timestamp 1666464484
transform 1 0 19688 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_214
timestamp 1666464484
transform 1 0 20792 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_223
timestamp 1666464484
transform 1 0 21620 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_238
timestamp 1666464484
transform 1 0 23000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1666464484
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_262
timestamp 1666464484
transform 1 0 25208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_271
timestamp 1666464484
transform 1 0 26036 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_283
timestamp 1666464484
transform 1 0 27140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_291
timestamp 1666464484
transform 1 0 27876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1666464484
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_318
timestamp 1666464484
transform 1 0 30360 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_324
timestamp 1666464484
transform 1 0 30912 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_329
timestamp 1666464484
transform 1 0 31372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_335
timestamp 1666464484
transform 1 0 31924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_339
timestamp 1666464484
transform 1 0 32292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_347
timestamp 1666464484
transform 1 0 33028 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_355
timestamp 1666464484
transform 1 0 33764 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1666464484
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_375
timestamp 1666464484
transform 1 0 35604 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_381
timestamp 1666464484
transform 1 0 36156 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_387
timestamp 1666464484
transform 1 0 36708 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_399
timestamp 1666464484
transform 1 0 37812 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_411
timestamp 1666464484
transform 1 0 38916 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666464484
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_157
timestamp 1666464484
transform 1 0 15548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1666464484
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_184
timestamp 1666464484
transform 1 0 18032 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_195
timestamp 1666464484
transform 1 0 19044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_202
timestamp 1666464484
transform 1 0 19688 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_208
timestamp 1666464484
transform 1 0 20240 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1666464484
transform 1 0 20976 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_234
timestamp 1666464484
transform 1 0 22632 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_242
timestamp 1666464484
transform 1 0 23368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_252
timestamp 1666464484
transform 1 0 24288 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1666464484
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1666464484
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1666464484
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1666464484
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_292
timestamp 1666464484
transform 1 0 27968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_299
timestamp 1666464484
transform 1 0 28612 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_309
timestamp 1666464484
transform 1 0 29532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1666464484
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_324
timestamp 1666464484
transform 1 0 30912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_333
timestamp 1666464484
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_345
timestamp 1666464484
transform 1 0 32844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_351
timestamp 1666464484
transform 1 0 33396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_359
timestamp 1666464484
transform 1 0 34132 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_363
timestamp 1666464484
transform 1 0 34500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1666464484
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666464484
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666464484
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1666464484
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1666464484
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_160
timestamp 1666464484
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1666464484
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_176
timestamp 1666464484
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_182
timestamp 1666464484
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_188
timestamp 1666464484
transform 1 0 18400 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1666464484
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_201
timestamp 1666464484
transform 1 0 19596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_204
timestamp 1666464484
transform 1 0 19872 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_216
timestamp 1666464484
transform 1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_224
timestamp 1666464484
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_227
timestamp 1666464484
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_239
timestamp 1666464484
transform 1 0 23092 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_264
timestamp 1666464484
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1666464484
transform 1 0 26036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_275
timestamp 1666464484
transform 1 0 26404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_279
timestamp 1666464484
transform 1 0 26772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_287
timestamp 1666464484
transform 1 0 27508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1666464484
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1666464484
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666464484
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_324
timestamp 1666464484
transform 1 0 30912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_328
timestamp 1666464484
transform 1 0 31280 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1666464484
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_346
timestamp 1666464484
transform 1 0 32936 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_354
timestamp 1666464484
transform 1 0 33672 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1666464484
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1666464484
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_376
timestamp 1666464484
transform 1 0 35696 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_382
timestamp 1666464484
transform 1 0 36248 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_394
timestamp 1666464484
transform 1 0 37352 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_406
timestamp 1666464484
transform 1 0 38456 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1666464484
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666464484
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666464484
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1666464484
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666464484
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666464484
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666464484
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666464484
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_155
timestamp 1666464484
transform 1 0 15364 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_159
timestamp 1666464484
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_173
timestamp 1666464484
transform 1 0 17020 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_176
timestamp 1666464484
transform 1 0 17296 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_184
timestamp 1666464484
transform 1 0 18032 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_206
timestamp 1666464484
transform 1 0 20056 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_216
timestamp 1666464484
transform 1 0 20976 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1666464484
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_234
timestamp 1666464484
transform 1 0 22632 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_243
timestamp 1666464484
transform 1 0 23460 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_251
timestamp 1666464484
transform 1 0 24196 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_258
timestamp 1666464484
transform 1 0 24840 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666464484
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_290
timestamp 1666464484
transform 1 0 27784 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_303
timestamp 1666464484
transform 1 0 28980 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_314
timestamp 1666464484
transform 1 0 29992 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_320
timestamp 1666464484
transform 1 0 30544 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_326
timestamp 1666464484
transform 1 0 31096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1666464484
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_345
timestamp 1666464484
transform 1 0 32844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_351
timestamp 1666464484
transform 1 0 33396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_355
timestamp 1666464484
transform 1 0 33764 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_379
timestamp 1666464484
transform 1 0 35972 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666464484
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666464484
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666464484
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1666464484
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1666464484
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1666464484
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_161
timestamp 1666464484
transform 1 0 15916 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_170
timestamp 1666464484
transform 1 0 16744 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_183
timestamp 1666464484
transform 1 0 17940 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_192
timestamp 1666464484
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_231
timestamp 1666464484
transform 1 0 22356 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_238
timestamp 1666464484
transform 1 0 23000 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_244
timestamp 1666464484
transform 1 0 23552 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1666464484
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_261
timestamp 1666464484
transform 1 0 25116 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_267
timestamp 1666464484
transform 1 0 25668 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_292
timestamp 1666464484
transform 1 0 27968 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_298
timestamp 1666464484
transform 1 0 28520 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1666464484
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_313
timestamp 1666464484
transform 1 0 29900 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_324
timestamp 1666464484
transform 1 0 30912 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_330
timestamp 1666464484
transform 1 0 31464 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_338
timestamp 1666464484
transform 1 0 32200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1666464484
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_369
timestamp 1666464484
transform 1 0 35052 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_393
timestamp 1666464484
transform 1 0 37260 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_405
timestamp 1666464484
transform 1 0 38364 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_417
timestamp 1666464484
transform 1 0 39468 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1666464484
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666464484
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666464484
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666464484
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1666464484
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_177
timestamp 1666464484
transform 1 0 17388 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_186
timestamp 1666464484
transform 1 0 18216 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1666464484
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_198
timestamp 1666464484
transform 1 0 19320 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_204
timestamp 1666464484
transform 1 0 19872 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_215
timestamp 1666464484
transform 1 0 20884 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_219
timestamp 1666464484
transform 1 0 21252 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1666464484
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_235
timestamp 1666464484
transform 1 0 22724 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_251
timestamp 1666464484
transform 1 0 24196 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_265
timestamp 1666464484
transform 1 0 25484 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1666464484
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_290
timestamp 1666464484
transform 1 0 27784 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_298
timestamp 1666464484
transform 1 0 28520 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_304
timestamp 1666464484
transform 1 0 29072 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_310
timestamp 1666464484
transform 1 0 29624 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_322
timestamp 1666464484
transform 1 0 30728 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1666464484
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_347
timestamp 1666464484
transform 1 0 33028 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_355
timestamp 1666464484
transform 1 0 33764 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_363
timestamp 1666464484
transform 1 0 34500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_372
timestamp 1666464484
transform 1 0 35328 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_378
timestamp 1666464484
transform 1 0 35880 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_384
timestamp 1666464484
transform 1 0 36432 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1666464484
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1666464484
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1666464484
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666464484
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666464484
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_168
timestamp 1666464484
transform 1 0 16560 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_174
timestamp 1666464484
transform 1 0 17112 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_177
timestamp 1666464484
transform 1 0 17388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_183
timestamp 1666464484
transform 1 0 17940 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1666464484
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_203
timestamp 1666464484
transform 1 0 19780 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_225
timestamp 1666464484
transform 1 0 21804 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_238
timestamp 1666464484
transform 1 0 23000 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1666464484
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_257
timestamp 1666464484
transform 1 0 24748 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_262
timestamp 1666464484
transform 1 0 25208 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_268
timestamp 1666464484
transform 1 0 25760 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_273
timestamp 1666464484
transform 1 0 26220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_280
timestamp 1666464484
transform 1 0 26864 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_286
timestamp 1666464484
transform 1 0 27416 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_294
timestamp 1666464484
transform 1 0 28152 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1666464484
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1666464484
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_323
timestamp 1666464484
transform 1 0 30820 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_329
timestamp 1666464484
transform 1 0 31372 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_335
timestamp 1666464484
transform 1 0 31924 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_338
timestamp 1666464484
transform 1 0 32200 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_349
timestamp 1666464484
transform 1 0 33212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_355
timestamp 1666464484
transform 1 0 33764 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1666464484
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_369
timestamp 1666464484
transform 1 0 35052 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_375
timestamp 1666464484
transform 1 0 35604 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_400
timestamp 1666464484
transform 1 0 37904 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_412
timestamp 1666464484
transform 1 0 39008 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666464484
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1666464484
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666464484
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666464484
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666464484
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_177
timestamp 1666464484
transform 1 0 17388 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_184
timestamp 1666464484
transform 1 0 18032 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_201
timestamp 1666464484
transform 1 0 19596 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_206
timestamp 1666464484
transform 1 0 20056 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_216
timestamp 1666464484
transform 1 0 20976 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1666464484
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_235
timestamp 1666464484
transform 1 0 22724 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_244
timestamp 1666464484
transform 1 0 23552 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_254
timestamp 1666464484
transform 1 0 24472 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_265
timestamp 1666464484
transform 1 0 25484 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_271
timestamp 1666464484
transform 1 0 26036 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1666464484
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_290
timestamp 1666464484
transform 1 0 27784 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_298
timestamp 1666464484
transform 1 0 28520 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_307
timestamp 1666464484
transform 1 0 29348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_311
timestamp 1666464484
transform 1 0 29716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_317
timestamp 1666464484
transform 1 0 30268 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_347
timestamp 1666464484
transform 1 0 33028 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_384
timestamp 1666464484
transform 1 0 36432 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666464484
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666464484
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1666464484
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1666464484
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1666464484
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_9
timestamp 1666464484
transform 1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666464484
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666464484
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_177
timestamp 1666464484
transform 1 0 17388 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_182
timestamp 1666464484
transform 1 0 17848 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1666464484
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_215
timestamp 1666464484
transform 1 0 20884 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_218
timestamp 1666464484
transform 1 0 21160 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_229
timestamp 1666464484
transform 1 0 22172 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_242
timestamp 1666464484
transform 1 0 23368 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_70_249
timestamp 1666464484
transform 1 0 24012 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_258
timestamp 1666464484
transform 1 0 24840 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_264
timestamp 1666464484
transform 1 0 25392 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_268
timestamp 1666464484
transform 1 0 25760 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_271
timestamp 1666464484
transform 1 0 26036 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_288
timestamp 1666464484
transform 1 0 27600 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666464484
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_313
timestamp 1666464484
transform 1 0 29900 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_326
timestamp 1666464484
transform 1 0 31096 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_330
timestamp 1666464484
transform 1 0 31464 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_338
timestamp 1666464484
transform 1 0 32200 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_345
timestamp 1666464484
transform 1 0 32844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_352
timestamp 1666464484
transform 1 0 33488 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_359
timestamp 1666464484
transform 1 0 34132 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_369
timestamp 1666464484
transform 1 0 35052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_373
timestamp 1666464484
transform 1 0 35420 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_376
timestamp 1666464484
transform 1 0 35696 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_382
timestamp 1666464484
transform 1 0 36248 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_394
timestamp 1666464484
transform 1 0 37352 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_406
timestamp 1666464484
transform 1 0 38456 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_418
timestamp 1666464484
transform 1 0 39560 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666464484
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_615
timestamp 1666464484
transform 1 0 57684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1666464484
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666464484
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666464484
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_189
timestamp 1666464484
transform 1 0 18492 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_199
timestamp 1666464484
transform 1 0 19412 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_211
timestamp 1666464484
transform 1 0 20516 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1666464484
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_234
timestamp 1666464484
transform 1 0 22632 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_243
timestamp 1666464484
transform 1 0 23460 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_247
timestamp 1666464484
transform 1 0 23828 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_255
timestamp 1666464484
transform 1 0 24564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_269
timestamp 1666464484
transform 1 0 25852 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1666464484
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_288
timestamp 1666464484
transform 1 0 27600 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_294
timestamp 1666464484
transform 1 0 28152 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_297
timestamp 1666464484
transform 1 0 28428 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_303
timestamp 1666464484
transform 1 0 28980 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_312
timestamp 1666464484
transform 1 0 29808 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_318
timestamp 1666464484
transform 1 0 30360 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_324
timestamp 1666464484
transform 1 0 30912 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_328
timestamp 1666464484
transform 1 0 31280 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_331
timestamp 1666464484
transform 1 0 31556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666464484
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_344
timestamp 1666464484
transform 1 0 32752 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_358
timestamp 1666464484
transform 1 0 34040 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_364
timestamp 1666464484
transform 1 0 34592 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_376
timestamp 1666464484
transform 1 0 35696 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_388
timestamp 1666464484
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666464484
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666464484
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1666464484
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1666464484
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666464484
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666464484
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666464484
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_207
timestamp 1666464484
transform 1 0 20148 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_213
timestamp 1666464484
transform 1 0 20700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1666464484
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_227
timestamp 1666464484
transform 1 0 21988 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_235
timestamp 1666464484
transform 1 0 22724 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1666464484
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_257
timestamp 1666464484
transform 1 0 24748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_268
timestamp 1666464484
transform 1 0 25760 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_272
timestamp 1666464484
transform 1 0 26128 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_275
timestamp 1666464484
transform 1 0 26404 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_287
timestamp 1666464484
transform 1 0 27508 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_293
timestamp 1666464484
transform 1 0 28060 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_297
timestamp 1666464484
transform 1 0 28428 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_306
timestamp 1666464484
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_314
timestamp 1666464484
transform 1 0 29992 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_324
timestamp 1666464484
transform 1 0 30912 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_330
timestamp 1666464484
transform 1 0 31464 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_347
timestamp 1666464484
transform 1 0 33028 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_356
timestamp 1666464484
transform 1 0 33856 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_371
timestamp 1666464484
transform 1 0 35236 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_378
timestamp 1666464484
transform 1 0 35880 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_384
timestamp 1666464484
transform 1 0 36432 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_396
timestamp 1666464484
transform 1 0 37536 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_408
timestamp 1666464484
transform 1 0 38640 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666464484
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666464484
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666464484
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666464484
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666464484
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_215
timestamp 1666464484
transform 1 0 20884 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_219
timestamp 1666464484
transform 1 0 21252 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1666464484
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_235
timestamp 1666464484
transform 1 0 22724 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_241
timestamp 1666464484
transform 1 0 23276 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_249
timestamp 1666464484
transform 1 0 24012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_256
timestamp 1666464484
transform 1 0 24656 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_263
timestamp 1666464484
transform 1 0 25300 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_272
timestamp 1666464484
transform 1 0 26128 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1666464484
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_295
timestamp 1666464484
transform 1 0 28244 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_307
timestamp 1666464484
transform 1 0 29348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_323
timestamp 1666464484
transform 1 0 30820 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1666464484
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_345
timestamp 1666464484
transform 1 0 32844 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_367
timestamp 1666464484
transform 1 0 34868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_379
timestamp 1666464484
transform 1 0 35972 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666464484
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666464484
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666464484
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666464484
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1666464484
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1666464484
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666464484
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_201
timestamp 1666464484
transform 1 0 19596 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_204
timestamp 1666464484
transform 1 0 19872 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_215
timestamp 1666464484
transform 1 0 20884 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_219
timestamp 1666464484
transform 1 0 21252 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_225
timestamp 1666464484
transform 1 0 21804 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_235
timestamp 1666464484
transform 1 0 22724 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_239
timestamp 1666464484
transform 1 0 23092 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_242
timestamp 1666464484
transform 1 0 23368 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1666464484
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_261
timestamp 1666464484
transform 1 0 25116 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_272
timestamp 1666464484
transform 1 0 26128 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_280
timestamp 1666464484
transform 1 0 26864 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_288
timestamp 1666464484
transform 1 0 27600 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_296
timestamp 1666464484
transform 1 0 28336 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1666464484
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_318
timestamp 1666464484
transform 1 0 30360 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_326
timestamp 1666464484
transform 1 0 31096 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_332
timestamp 1666464484
transform 1 0 31648 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_340
timestamp 1666464484
transform 1 0 32384 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_344
timestamp 1666464484
transform 1 0 32752 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_348
timestamp 1666464484
transform 1 0 33120 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 1666464484
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_372
timestamp 1666464484
transform 1 0 35328 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_378
timestamp 1666464484
transform 1 0 35880 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_390
timestamp 1666464484
transform 1 0 36984 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_402
timestamp 1666464484
transform 1 0 38088 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_414
timestamp 1666464484
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666464484
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666464484
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666464484
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666464484
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_199
timestamp 1666464484
transform 1 0 19412 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_211
timestamp 1666464484
transform 1 0 20516 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_219
timestamp 1666464484
transform 1 0 21252 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_229
timestamp 1666464484
transform 1 0 22172 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_241
timestamp 1666464484
transform 1 0 23276 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_250
timestamp 1666464484
transform 1 0 24104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_257
timestamp 1666464484
transform 1 0 24748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_263
timestamp 1666464484
transform 1 0 25300 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_271
timestamp 1666464484
transform 1 0 26036 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_277
timestamp 1666464484
transform 1 0 26588 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_288
timestamp 1666464484
transform 1 0 27600 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_315
timestamp 1666464484
transform 1 0 30084 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_322
timestamp 1666464484
transform 1 0 30728 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_332
timestamp 1666464484
transform 1 0 31648 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_345
timestamp 1666464484
transform 1 0 32844 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_353
timestamp 1666464484
transform 1 0 33580 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_360
timestamp 1666464484
transform 1 0 34224 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_366
timestamp 1666464484
transform 1 0 34776 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_372
timestamp 1666464484
transform 1 0 35328 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_384
timestamp 1666464484
transform 1 0 36432 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666464484
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666464484
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666464484
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666464484
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1666464484
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1666464484
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666464484
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666464484
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_185
timestamp 1666464484
transform 1 0 18124 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1666464484
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_212
timestamp 1666464484
transform 1 0 20608 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_222
timestamp 1666464484
transform 1 0 21528 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_234
timestamp 1666464484
transform 1 0 22632 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_242
timestamp 1666464484
transform 1 0 23368 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1666464484
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_258
timestamp 1666464484
transform 1 0 24840 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_279
timestamp 1666464484
transform 1 0 26772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_290
timestamp 1666464484
transform 1 0 27784 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_297
timestamp 1666464484
transform 1 0 28428 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1666464484
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_318
timestamp 1666464484
transform 1 0 30360 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_328
timestamp 1666464484
transform 1 0 31280 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_336
timestamp 1666464484
transform 1 0 32016 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_340
timestamp 1666464484
transform 1 0 32384 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_347
timestamp 1666464484
transform 1 0 33028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_370
timestamp 1666464484
transform 1 0 35144 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_376
timestamp 1666464484
transform 1 0 35696 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_388
timestamp 1666464484
transform 1 0 36800 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_400
timestamp 1666464484
transform 1 0 37904 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_412
timestamp 1666464484
transform 1 0 39008 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666464484
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1666464484
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666464484
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666464484
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666464484
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666464484
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_200
timestamp 1666464484
transform 1 0 19504 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_208
timestamp 1666464484
transform 1 0 20240 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_211
timestamp 1666464484
transform 1 0 20516 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_219
timestamp 1666464484
transform 1 0 21252 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_230
timestamp 1666464484
transform 1 0 22264 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_234
timestamp 1666464484
transform 1 0 22632 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_238
timestamp 1666464484
transform 1 0 23000 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_246
timestamp 1666464484
transform 1 0 23736 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_255
timestamp 1666464484
transform 1 0 24564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_265
timestamp 1666464484
transform 1 0 25484 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_277
timestamp 1666464484
transform 1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_287
timestamp 1666464484
transform 1 0 27508 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_294
timestamp 1666464484
transform 1 0 28152 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_312
timestamp 1666464484
transform 1 0 29808 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_316
timestamp 1666464484
transform 1 0 30176 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_320
timestamp 1666464484
transform 1 0 30544 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_330
timestamp 1666464484
transform 1 0 31464 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_342
timestamp 1666464484
transform 1 0 32568 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_346
timestamp 1666464484
transform 1 0 32936 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_360
timestamp 1666464484
transform 1 0 34224 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_369
timestamp 1666464484
transform 1 0 35052 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_381
timestamp 1666464484
transform 1 0 36156 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_389
timestamp 1666464484
transform 1 0 36892 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1666464484
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1666464484
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666464484
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666464484
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1666464484
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1666464484
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666464484
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_201
timestamp 1666464484
transform 1 0 19596 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_207
timestamp 1666464484
transform 1 0 20148 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_213
timestamp 1666464484
transform 1 0 20700 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_222
timestamp 1666464484
transform 1 0 21528 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_237
timestamp 1666464484
transform 1 0 22908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1666464484
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_259
timestamp 1666464484
transform 1 0 24932 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_271
timestamp 1666464484
transform 1 0 26036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_280
timestamp 1666464484
transform 1 0 26864 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_289
timestamp 1666464484
transform 1 0 27692 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_297
timestamp 1666464484
transform 1 0 28428 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1666464484
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_316
timestamp 1666464484
transform 1 0 30176 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_330
timestamp 1666464484
transform 1 0 31464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_339
timestamp 1666464484
transform 1 0 32292 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_354
timestamp 1666464484
transform 1 0 33672 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_360
timestamp 1666464484
transform 1 0 34224 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_369
timestamp 1666464484
transform 1 0 35052 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_381
timestamp 1666464484
transform 1 0 36156 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_393
timestamp 1666464484
transform 1 0 37260 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_405
timestamp 1666464484
transform 1 0 38364 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1666464484
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1666464484
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666464484
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666464484
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_213
timestamp 1666464484
transform 1 0 20700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1666464484
transform 1 0 21528 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_235
timestamp 1666464484
transform 1 0 22724 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_245
timestamp 1666464484
transform 1 0 23644 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_269
timestamp 1666464484
transform 1 0 25852 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1666464484
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_290
timestamp 1666464484
transform 1 0 27784 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_304
timestamp 1666464484
transform 1 0 29072 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_310
timestamp 1666464484
transform 1 0 29624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_317
timestamp 1666464484
transform 1 0 30268 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_328
timestamp 1666464484
transform 1 0 31280 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1666464484
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_348
timestamp 1666464484
transform 1 0 33120 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_374
timestamp 1666464484
transform 1 0 35512 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_380
timestamp 1666464484
transform 1 0 36064 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1666464484
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1666464484
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666464484
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1666464484
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1666464484
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_211
timestamp 1666464484
transform 1 0 20516 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_217
timestamp 1666464484
transform 1 0 21068 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_227
timestamp 1666464484
transform 1 0 21988 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_237
timestamp 1666464484
transform 1 0 22908 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_249
timestamp 1666464484
transform 1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_261
timestamp 1666464484
transform 1 0 25116 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_271
timestamp 1666464484
transform 1 0 26036 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_282
timestamp 1666464484
transform 1 0 27048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_293
timestamp 1666464484
transform 1 0 28060 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1666464484
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_327
timestamp 1666464484
transform 1 0 31188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_347
timestamp 1666464484
transform 1 0 33028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1666464484
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_369
timestamp 1666464484
transform 1 0 35052 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_381
timestamp 1666464484
transform 1 0 36156 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_393
timestamp 1666464484
transform 1 0 37260 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_405
timestamp 1666464484
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1666464484
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1666464484
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666464484
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1666464484
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_615
timestamp 1666464484
transform 1 0 57684 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1666464484
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_9
timestamp 1666464484
transform 1 0 1932 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1666464484
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_229
timestamp 1666464484
transform 1 0 22172 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_234
timestamp 1666464484
transform 1 0 22632 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_242
timestamp 1666464484
transform 1 0 23368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_246
timestamp 1666464484
transform 1 0 23736 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_253
timestamp 1666464484
transform 1 0 24380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_257
timestamp 1666464484
transform 1 0 24748 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_265
timestamp 1666464484
transform 1 0 25484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1666464484
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_289
timestamp 1666464484
transform 1 0 27692 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_300
timestamp 1666464484
transform 1 0 28704 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_304
timestamp 1666464484
transform 1 0 29072 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_307
timestamp 1666464484
transform 1 0 29348 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_317
timestamp 1666464484
transform 1 0 30268 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_327
timestamp 1666464484
transform 1 0 31188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_333
timestamp 1666464484
transform 1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_345
timestamp 1666464484
transform 1 0 32844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_355
timestamp 1666464484
transform 1 0 33764 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_367
timestamp 1666464484
transform 1 0 34868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_379
timestamp 1666464484
transform 1 0 35972 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1666464484
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1666464484
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_230
timestamp 1666464484
transform 1 0 22264 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_244
timestamp 1666464484
transform 1 0 23552 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1666464484
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_257
timestamp 1666464484
transform 1 0 24748 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_264
timestamp 1666464484
transform 1 0 25392 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_270
timestamp 1666464484
transform 1 0 25944 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_280
timestamp 1666464484
transform 1 0 26864 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_286
timestamp 1666464484
transform 1 0 27416 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_294
timestamp 1666464484
transform 1 0 28152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1666464484
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_315
timestamp 1666464484
transform 1 0 30084 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_318
timestamp 1666464484
transform 1 0 30360 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_335
timestamp 1666464484
transform 1 0 31924 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_343
timestamp 1666464484
transform 1 0 32660 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_353
timestamp 1666464484
transform 1 0 33580 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_359
timestamp 1666464484
transform 1 0 34132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1666464484
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1666464484
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1666464484
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_233
timestamp 1666464484
transform 1 0 22540 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_239
timestamp 1666464484
transform 1 0 23092 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_83_247
timestamp 1666464484
transform 1 0 23828 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_255
timestamp 1666464484
transform 1 0 24564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_262
timestamp 1666464484
transform 1 0 25208 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_268
timestamp 1666464484
transform 1 0 25760 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_301
timestamp 1666464484
transform 1 0 28796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_308
timestamp 1666464484
transform 1 0 29440 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_316
timestamp 1666464484
transform 1 0 30176 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_319
timestamp 1666464484
transform 1 0 30452 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_345
timestamp 1666464484
transform 1 0 32844 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_352
timestamp 1666464484
transform 1 0 33488 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_358
timestamp 1666464484
transform 1 0 34040 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_370
timestamp 1666464484
transform 1 0 35144 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_382
timestamp 1666464484
transform 1 0 36248 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_390
timestamp 1666464484
transform 1 0 36984 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1666464484
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1666464484
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_313
timestamp 1666464484
transform 1 0 29900 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_325
timestamp 1666464484
transform 1 0 31004 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_337
timestamp 1666464484
transform 1 0 32108 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_349
timestamp 1666464484
transform 1 0 33212 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_361
timestamp 1666464484
transform 1 0 34316 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1666464484
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1666464484
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1666464484
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1666464484
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1666464484
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1666464484
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1666464484
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1666464484
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1666464484
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1666464484
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1666464484
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1666464484
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1666464484
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1666464484
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1666464484
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_9
timestamp 1666464484
transform 1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1666464484
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1666464484
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1666464484
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_614
timestamp 1666464484
transform 1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1666464484
transform 1 0 58420 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1666464484
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1666464484
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1666464484
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1666464484
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1666464484
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1666464484
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1666464484
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1666464484
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1666464484
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1666464484
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1666464484
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1666464484
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1666464484
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1666464484
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1666464484
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1666464484
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1666464484
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1666464484
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1666464484
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1666464484
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1666464484
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1666464484
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1666464484
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1666464484
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1666464484
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1666464484
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1666464484
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1666464484
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1666464484
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1666464484
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1666464484
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1666464484
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1666464484
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1666464484
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1666464484
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1666464484
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1666464484
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1666464484
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1666464484
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1666464484
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1666464484
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1666464484
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1666464484
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1666464484
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1666464484
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1666464484
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1666464484
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1666464484
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1666464484
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1666464484
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1666464484
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1666464484
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1666464484
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1666464484
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1666464484
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1666464484
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1666464484
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1666464484
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1666464484
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1666464484
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1666464484
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1666464484
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1666464484
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1666464484
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1666464484
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1666464484
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1666464484
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1666464484
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1666464484
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1666464484
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1666464484
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1666464484
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1666464484
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1666464484
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1666464484
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1666464484
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1666464484
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1666464484
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1666464484
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1666464484
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1666464484
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1666464484
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1666464484
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1666464484
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1666464484
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1666464484
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1666464484
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1666464484
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1666464484
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1666464484
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1666464484
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1666464484
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1666464484
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1666464484
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1666464484
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1666464484
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1666464484
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1666464484
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1666464484
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1666464484
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1666464484
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1666464484
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1666464484
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1666464484
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1666464484
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1666464484
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1666464484
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1666464484
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1666464484
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1666464484
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1666464484
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1666464484
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1666464484
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1666464484
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1666464484
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1666464484
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1666464484
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1666464484
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1666464484
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1666464484
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1666464484
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1666464484
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1666464484
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1666464484
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1666464484
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1666464484
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1666464484
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1666464484
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1666464484
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1666464484
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1666464484
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1666464484
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1666464484
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1666464484
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1666464484
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1666464484
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1666464484
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1666464484
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1666464484
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1666464484
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1666464484
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1666464484
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1666464484
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1666464484
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1666464484
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1666464484
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1666464484
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1666464484
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1666464484
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1666464484
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1666464484
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1666464484
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1666464484
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1666464484
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1666464484
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1666464484
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1666464484
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1666464484
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1666464484
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1666464484
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1666464484
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1666464484
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1666464484
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1666464484
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1666464484
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1666464484
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1666464484
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1666464484
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1666464484
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1666464484
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1666464484
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1666464484
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1666464484
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1666464484
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1666464484
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1666464484
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1666464484
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_11
timestamp 1666464484
transform 1 0 2116 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_17
timestamp 1666464484
transform 1 0 2668 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_25
timestamp 1666464484
transform 1 0 3404 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1666464484
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1666464484
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1666464484
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1666464484
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1666464484
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1666464484
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1666464484
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1666464484
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1666464484
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1666464484
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1666464484
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1666464484
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1666464484
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1666464484
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1666464484
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1666464484
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1666464484
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1666464484
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1666464484
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1666464484
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1666464484
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1666464484
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1666464484
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1666464484
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_372
timestamp 1666464484
transform 1 0 35328 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_378
timestamp 1666464484
transform 1 0 35880 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_390
timestamp 1666464484
transform 1 0 36984 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_402
timestamp 1666464484
transform 1 0 38088 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_414
timestamp 1666464484
transform 1 0 39192 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1666464484
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1666464484
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1666464484
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1666464484
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1666464484
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1666464484
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1666464484
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1666464484
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1666464484
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1666464484
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1666464484
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1666464484
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_615
timestamp 1666464484
transform 1 0 57684 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1666464484
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_9
timestamp 1666464484
transform 1 0 1932 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_21
timestamp 1666464484
transform 1 0 3036 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1666464484
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_41
timestamp 1666464484
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1666464484
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1666464484
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1666464484
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_91
timestamp 1666464484
transform 1 0 9476 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1666464484
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1666464484
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_125
timestamp 1666464484
transform 1 0 12604 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_133
timestamp 1666464484
transform 1 0 13340 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1666464484
transform 1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_141
timestamp 1666464484
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_147
timestamp 1666464484
transform 1 0 14628 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_159
timestamp 1666464484
transform 1 0 15732 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1666464484
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_197
timestamp 1666464484
transform 1 0 19228 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_203
timestamp 1666464484
transform 1 0 19780 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1666464484
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1666464484
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1666464484
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1666464484
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_259
timestamp 1666464484
transform 1 0 24932 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_265
timestamp 1666464484
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1666464484
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1666464484
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1666464484
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_101_309
timestamp 1666464484
transform 1 0 29532 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_314
timestamp 1666464484
transform 1 0 29992 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_322
timestamp 1666464484
transform 1 0 30728 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_334
timestamp 1666464484
transform 1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1666464484
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1666464484
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_365
timestamp 1666464484
transform 1 0 34684 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_373
timestamp 1666464484
transform 1 0 35420 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_378
timestamp 1666464484
transform 1 0 35880 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_390
timestamp 1666464484
transform 1 0 36984 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1666464484
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1666464484
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_429
timestamp 1666464484
transform 1 0 40572 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_433
timestamp 1666464484
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1666464484
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1666464484
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1666464484
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1666464484
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_477
timestamp 1666464484
transform 1 0 44988 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_485
timestamp 1666464484
transform 1 0 45724 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_489
timestamp 1666464484
transform 1 0 46092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1666464484
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1666464484
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1666464484
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1666464484
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_553
timestamp 1666464484
transform 1 0 51980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_558
timestamp 1666464484
transform 1 0 52440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_567
timestamp 1666464484
transform 1 0 53268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_579
timestamp 1666464484
transform 1 0 54372 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_587
timestamp 1666464484
transform 1 0 55108 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_601
timestamp 1666464484
transform 1 0 56396 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_609
timestamp 1666464484
transform 1 0 57132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1666464484
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1666464484
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0990_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 45724 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0991_
timestamp 1666464484
transform 1 0 43700 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0992_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36800 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0993_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 38548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0994_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37444 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _0995_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 40204 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_1  _0996_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _0997_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 42320 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0998_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36432 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _0999_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 39284 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_4  _1000_
timestamp 1666464484
transform 1 0 38548 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1001_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36616 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1002_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31004 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1003_
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1004_
timestamp 1666464484
transform 1 0 46000 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1005_
timestamp 1666464484
transform 1 0 42964 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _1006_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44620 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1666464484
transform -1 0 31464 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1008_
timestamp 1666464484
transform -1 0 30912 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1009_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1010_
timestamp 1666464484
transform 1 0 28612 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1011_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22264 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1012_
timestamp 1666464484
transform -1 0 23368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1013_
timestamp 1666464484
transform 1 0 32476 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1014_
timestamp 1666464484
transform -1 0 25208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1015_
timestamp 1666464484
transform -1 0 25208 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1016_
timestamp 1666464484
transform -1 0 33488 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1017_
timestamp 1666464484
transform -1 0 31188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1018_
timestamp 1666464484
transform -1 0 31464 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1019_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30636 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 1666464484
transform -1 0 28612 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30452 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1022_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1666464484
transform -1 0 29808 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1666464484
transform 1 0 35604 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1666464484
transform -1 0 30176 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1026_
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1027_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31280 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29348 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_4  _1029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30176 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_2  _1030_
timestamp 1666464484
transform -1 0 33764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30360 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1032_
timestamp 1666464484
transform 1 0 27876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1033_
timestamp 1666464484
transform -1 0 30544 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1034_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1666464484
transform 1 0 33304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1036_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1037_
timestamp 1666464484
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1666464484
transform 1 0 26128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1039_
timestamp 1666464484
transform -1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1040_
timestamp 1666464484
transform 1 0 19412 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 1666464484
transform 1 0 27140 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1666464484
transform -1 0 26680 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1666464484
transform -1 0 26680 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1044_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1047_
timestamp 1666464484
transform 1 0 25024 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1666464484
transform -1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1049_
timestamp 1666464484
transform -1 0 27600 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1666464484
transform -1 0 26220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1666464484
transform -1 0 32568 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1052_
timestamp 1666464484
transform 1 0 32292 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1053_
timestamp 1666464484
transform -1 0 33580 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1054_
timestamp 1666464484
transform 1 0 32292 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1055_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34224 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1666464484
transform 1 0 22356 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1057_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1058_
timestamp 1666464484
transform 1 0 23368 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32384 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32568 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1061_
timestamp 1666464484
transform 1 0 33212 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1062_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27416 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1063_
timestamp 1666464484
transform -1 0 26680 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1064_
timestamp 1666464484
transform -1 0 26864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1065_
timestamp 1666464484
transform 1 0 30912 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1066_
timestamp 1666464484
transform -1 0 25484 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1067_
timestamp 1666464484
transform -1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1068_
timestamp 1666464484
transform -1 0 34224 0 1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__a31o_1  _1069_
timestamp 1666464484
transform 1 0 27140 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _1071_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1666464484
transform 1 0 17020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1073_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34224 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1074_
timestamp 1666464484
transform 1 0 34868 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1075_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34592 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32476 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1077_
timestamp 1666464484
transform -1 0 33672 0 1 44608
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1078_
timestamp 1666464484
transform 1 0 23736 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1079_
timestamp 1666464484
transform 1 0 21528 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1080_
timestamp 1666464484
transform -1 0 22632 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1081_
timestamp 1666464484
transform -1 0 27968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1082_
timestamp 1666464484
transform -1 0 20056 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1666464484
transform 1 0 28060 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1084_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22172 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1666464484
transform -1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1086_
timestamp 1666464484
transform -1 0 23460 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1087_
timestamp 1666464484
transform 1 0 31096 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1088_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28152 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1089_
timestamp 1666464484
transform 1 0 30268 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 1666464484
transform 1 0 26312 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1666464484
transform -1 0 27600 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1092_
timestamp 1666464484
transform 1 0 20240 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _1093_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_2  _1094_
timestamp 1666464484
transform 1 0 26404 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1095_
timestamp 1666464484
transform -1 0 24380 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1096_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23644 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1097_
timestamp 1666464484
transform -1 0 24840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1098_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1666464484
transform 1 0 23644 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1100_
timestamp 1666464484
transform 1 0 23736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _1101_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23552 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1102_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23000 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1103_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30728 0 1 46784
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1666464484
transform -1 0 22264 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1105_
timestamp 1666464484
transform -1 0 25392 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1106_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1107_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25300 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1108_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1109_
timestamp 1666464484
transform -1 0 21620 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1110_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28612 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1666464484
transform 1 0 19412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1112_
timestamp 1666464484
transform -1 0 19044 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1113_
timestamp 1666464484
transform -1 0 18032 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1114_
timestamp 1666464484
transform 1 0 20424 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1115_
timestamp 1666464484
transform 1 0 20424 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1116_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29164 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _1117_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33488 0 -1 45696
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _1118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33028 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1119_
timestamp 1666464484
transform 1 0 23092 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_2  _1121_
timestamp 1666464484
transform 1 0 28152 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1122_
timestamp 1666464484
transform 1 0 21988 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1123_
timestamp 1666464484
transform -1 0 30268 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1124_
timestamp 1666464484
transform 1 0 23368 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1126_
timestamp 1666464484
transform -1 0 24656 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1127_
timestamp 1666464484
transform -1 0 35144 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1666464484
transform -1 0 20056 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1129_
timestamp 1666464484
transform 1 0 20884 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1130_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19780 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 1666464484
transform 1 0 19412 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1666464484
transform 1 0 19412 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1133_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19688 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1134_
timestamp 1666464484
transform -1 0 25484 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1135_
timestamp 1666464484
transform 1 0 27232 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1136_
timestamp 1666464484
transform -1 0 21528 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1137_
timestamp 1666464484
transform -1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1138_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21528 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1139_
timestamp 1666464484
transform 1 0 20884 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1140_
timestamp 1666464484
transform -1 0 22264 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1141_
timestamp 1666464484
transform -1 0 28888 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1142_
timestamp 1666464484
transform 1 0 20976 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _1143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19780 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1666464484
transform -1 0 18676 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1145_
timestamp 1666464484
transform -1 0 18308 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1666464484
transform -1 0 17296 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1147_
timestamp 1666464484
transform -1 0 17480 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1666464484
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1149_
timestamp 1666464484
transform 1 0 23828 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1150_
timestamp 1666464484
transform -1 0 27692 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1666464484
transform 1 0 26496 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1152_
timestamp 1666464484
transform 1 0 27140 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 1666464484
transform 1 0 29716 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1154_
timestamp 1666464484
transform -1 0 29256 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _1155_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30176 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1156_
timestamp 1666464484
transform -1 0 29164 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1157_
timestamp 1666464484
transform -1 0 31648 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1158_
timestamp 1666464484
transform 1 0 29716 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1159_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25392 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1160_
timestamp 1666464484
transform 1 0 16836 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1161_
timestamp 1666464484
transform 1 0 16100 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1162_
timestamp 1666464484
transform 1 0 16100 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1666464484
transform -1 0 16376 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1164_
timestamp 1666464484
transform 1 0 28704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1165_
timestamp 1666464484
transform 1 0 28796 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1166_
timestamp 1666464484
transform 1 0 28612 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1167_
timestamp 1666464484
transform -1 0 29256 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_4  _1168_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31188 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_1  _1169_
timestamp 1666464484
transform -1 0 28980 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 1666464484
transform -1 0 21528 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1171_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22356 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1172_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1173_
timestamp 1666464484
transform -1 0 20976 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1174_
timestamp 1666464484
transform 1 0 27232 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1175_
timestamp 1666464484
transform -1 0 27692 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1176_
timestamp 1666464484
transform 1 0 27416 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1177_
timestamp 1666464484
transform -1 0 27968 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1178_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1179_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1180_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29900 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 1666464484
transform -1 0 20884 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1182_
timestamp 1666464484
transform 1 0 24564 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1183_
timestamp 1666464484
transform -1 0 23000 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1184_
timestamp 1666464484
transform -1 0 21804 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1185_
timestamp 1666464484
transform 1 0 22264 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1186_
timestamp 1666464484
transform -1 0 23000 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1187_
timestamp 1666464484
transform 1 0 22264 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1188_
timestamp 1666464484
transform -1 0 22632 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1189_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22356 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1190_
timestamp 1666464484
transform 1 0 22724 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1191_
timestamp 1666464484
transform 1 0 22356 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1192_
timestamp 1666464484
transform -1 0 32292 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1193_
timestamp 1666464484
transform 1 0 23276 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1194_
timestamp 1666464484
transform -1 0 22724 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27600 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1196_
timestamp 1666464484
transform 1 0 26128 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1197_
timestamp 1666464484
transform 1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1198_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22632 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1199_
timestamp 1666464484
transform 1 0 20608 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1200_
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1666464484
transform -1 0 28152 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1202_
timestamp 1666464484
transform -1 0 29164 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1204_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23000 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1666464484
transform -1 0 23828 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1206_
timestamp 1666464484
transform 1 0 20240 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_4  _1207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19872 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1208_
timestamp 1666464484
transform -1 0 17388 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1210_
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1211_
timestamp 1666464484
transform 1 0 31648 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1212_
timestamp 1666464484
transform 1 0 25392 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_1  _1213_
timestamp 1666464484
transform 1 0 24104 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1666464484
transform 1 0 27232 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1215_
timestamp 1666464484
transform -1 0 27784 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1216_
timestamp 1666464484
transform -1 0 29808 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1217_
timestamp 1666464484
transform 1 0 28152 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1218_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__o211ai_4  _1219_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25208 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__a21oi_1  _1220_
timestamp 1666464484
transform 1 0 17664 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1221_
timestamp 1666464484
transform -1 0 18768 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1222_
timestamp 1666464484
transform -1 0 17940 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1223_
timestamp 1666464484
transform 1 0 15088 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1224_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16100 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1225_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16100 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1226_
timestamp 1666464484
transform 1 0 17204 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1227_
timestamp 1666464484
transform -1 0 18860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1228_
timestamp 1666464484
transform 1 0 14904 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1666464484
transform -1 0 15824 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1230_
timestamp 1666464484
transform -1 0 14996 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1231_
timestamp 1666464484
transform 1 0 14720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp 1666464484
transform -1 0 14352 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1233_
timestamp 1666464484
transform 1 0 15640 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1234_
timestamp 1666464484
transform -1 0 16100 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23092 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1666464484
transform -1 0 21252 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1666464484
transform 1 0 20792 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1238_
timestamp 1666464484
transform -1 0 28152 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1239_
timestamp 1666464484
transform -1 0 26680 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1240_
timestamp 1666464484
transform -1 0 26680 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1666464484
transform -1 0 25024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1242_
timestamp 1666464484
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1666464484
transform 1 0 28520 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1244_
timestamp 1666464484
transform 1 0 24380 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1245_
timestamp 1666464484
transform -1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1246_
timestamp 1666464484
transform 1 0 18124 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1247_
timestamp 1666464484
transform 1 0 30544 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1248_
timestamp 1666464484
transform -1 0 29256 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1249_
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1250_
timestamp 1666464484
transform 1 0 28152 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1251_
timestamp 1666464484
transform 1 0 33396 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1666464484
transform 1 0 29716 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1253_
timestamp 1666464484
transform 1 0 30268 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1254_
timestamp 1666464484
transform -1 0 30268 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1255_
timestamp 1666464484
transform 1 0 28612 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1256_
timestamp 1666464484
transform -1 0 18216 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1257_
timestamp 1666464484
transform -1 0 18308 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1258_
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1259_
timestamp 1666464484
transform -1 0 21252 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1260_
timestamp 1666464484
transform -1 0 19504 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1261_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18400 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1262_
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1263_
timestamp 1666464484
transform 1 0 25484 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1264_
timestamp 1666464484
transform -1 0 24104 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1265_
timestamp 1666464484
transform 1 0 23460 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1266_
timestamp 1666464484
transform -1 0 24104 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1666464484
transform 1 0 19780 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1268_
timestamp 1666464484
transform 1 0 18216 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1269_
timestamp 1666464484
transform 1 0 18400 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1270_
timestamp 1666464484
transform -1 0 18768 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1271_
timestamp 1666464484
transform -1 0 17296 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1272_
timestamp 1666464484
transform 1 0 15548 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1666464484
transform -1 0 16284 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1274_
timestamp 1666464484
transform -1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1275_
timestamp 1666464484
transform -1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1276_
timestamp 1666464484
transform -1 0 16284 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_1  _1277_
timestamp 1666464484
transform -1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1278_
timestamp 1666464484
transform 1 0 26772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_2  _1279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19412 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__o41ai_4  _1280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 38080
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1281_
timestamp 1666464484
transform 1 0 33396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1666464484
transform 1 0 33580 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1283_
timestamp 1666464484
transform 1 0 31188 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1285_
timestamp 1666464484
transform -1 0 29256 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1286_
timestamp 1666464484
transform 1 0 30544 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _1287_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30084 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1288_
timestamp 1666464484
transform 1 0 19780 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1289_
timestamp 1666464484
transform -1 0 20700 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1290_
timestamp 1666464484
transform -1 0 23828 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1291_
timestamp 1666464484
transform 1 0 23460 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1292_
timestamp 1666464484
transform 1 0 24564 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1666464484
transform -1 0 26036 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1666464484
transform 1 0 28612 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1295_
timestamp 1666464484
transform 1 0 24564 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1666464484
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1297_
timestamp 1666464484
transform -1 0 23828 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 1666464484
transform -1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1299_
timestamp 1666464484
transform 1 0 24564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1300_
timestamp 1666464484
transform 1 0 23184 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19320 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1302_
timestamp 1666464484
transform 1 0 20424 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1303_
timestamp 1666464484
transform -1 0 27600 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1304_
timestamp 1666464484
transform 1 0 25852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1305_
timestamp 1666464484
transform 1 0 28152 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1307_
timestamp 1666464484
transform 1 0 27508 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1308_
timestamp 1666464484
transform 1 0 27140 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1309_
timestamp 1666464484
transform 1 0 19412 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1310_
timestamp 1666464484
transform 1 0 19872 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1311_
timestamp 1666464484
transform 1 0 20148 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1666464484
transform -1 0 20792 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1666464484
transform -1 0 19964 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1314_
timestamp 1666464484
transform 1 0 18216 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1315_
timestamp 1666464484
transform 1 0 18032 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1316_
timestamp 1666464484
transform -1 0 18492 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1317_
timestamp 1666464484
transform 1 0 16928 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1318_
timestamp 1666464484
transform 1 0 17572 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1319_
timestamp 1666464484
transform -1 0 18952 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1320_
timestamp 1666464484
transform -1 0 21344 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1321_
timestamp 1666464484
transform -1 0 23460 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1322_
timestamp 1666464484
transform -1 0 23000 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1323_
timestamp 1666464484
transform -1 0 22540 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1324_
timestamp 1666464484
transform 1 0 22816 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1325_
timestamp 1666464484
transform -1 0 21988 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1666464484
transform 1 0 25760 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1327_
timestamp 1666464484
transform 1 0 31280 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1328_
timestamp 1666464484
transform 1 0 32292 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1329_
timestamp 1666464484
transform 1 0 32292 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1330_
timestamp 1666464484
transform 1 0 25116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1331_
timestamp 1666464484
transform -1 0 23276 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1332_
timestamp 1666464484
transform -1 0 23000 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1333_
timestamp 1666464484
transform 1 0 24380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1666464484
transform 1 0 24196 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1666464484
transform 1 0 27968 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1336_
timestamp 1666464484
transform -1 0 25668 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1337_
timestamp 1666464484
transform 1 0 22356 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1338_
timestamp 1666464484
transform -1 0 21344 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1339_
timestamp 1666464484
transform 1 0 20792 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1340_
timestamp 1666464484
transform 1 0 21712 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1341_
timestamp 1666464484
transform -1 0 21988 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1342_
timestamp 1666464484
transform 1 0 20884 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1666464484
transform -1 0 20884 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1344_
timestamp 1666464484
transform -1 0 20240 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1345_
timestamp 1666464484
transform 1 0 17940 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1346_
timestamp 1666464484
transform 1 0 17756 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1347_
timestamp 1666464484
transform 1 0 24748 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1348_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1666464484
transform 1 0 32476 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1350_
timestamp 1666464484
transform 1 0 33856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1351_
timestamp 1666464484
transform 1 0 32292 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1352_
timestamp 1666464484
transform 1 0 31556 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1353_
timestamp 1666464484
transform 1 0 32292 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_1  _1354_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30268 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30728 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1356_
timestamp 1666464484
transform -1 0 31740 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1357_
timestamp 1666464484
transform -1 0 28704 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1358_
timestamp 1666464484
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1359_
timestamp 1666464484
transform 1 0 24932 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1360_
timestamp 1666464484
transform 1 0 24840 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1361_
timestamp 1666464484
transform -1 0 22724 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1362_
timestamp 1666464484
transform 1 0 23920 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1363_
timestamp 1666464484
transform 1 0 25576 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1364_
timestamp 1666464484
transform -1 0 24104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1365_
timestamp 1666464484
transform 1 0 24564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1366_
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1367_
timestamp 1666464484
transform 1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1368_
timestamp 1666464484
transform 1 0 32292 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1369_
timestamp 1666464484
transform -1 0 33028 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1370_
timestamp 1666464484
transform 1 0 27048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1371_
timestamp 1666464484
transform 1 0 31004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1372_
timestamp 1666464484
transform -1 0 32200 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _1373_
timestamp 1666464484
transform -1 0 22356 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1374_
timestamp 1666464484
transform -1 0 31832 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1375_
timestamp 1666464484
transform -1 0 23828 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1376_
timestamp 1666464484
transform -1 0 23736 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1666464484
transform -1 0 22816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1378_
timestamp 1666464484
transform -1 0 22632 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1379_
timestamp 1666464484
transform -1 0 22172 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1380_
timestamp 1666464484
transform -1 0 22632 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1381_
timestamp 1666464484
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1382_
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1383_
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1384_
timestamp 1666464484
transform -1 0 21252 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1385_
timestamp 1666464484
transform 1 0 25024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1666464484
transform 1 0 26772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1387_
timestamp 1666464484
transform 1 0 27968 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1388_
timestamp 1666464484
transform 1 0 29716 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1389_
timestamp 1666464484
transform -1 0 30912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1390_
timestamp 1666464484
transform -1 0 31188 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1391_
timestamp 1666464484
transform -1 0 27600 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1392_
timestamp 1666464484
transform -1 0 27968 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1393_
timestamp 1666464484
transform -1 0 28520 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1394_
timestamp 1666464484
transform -1 0 28980 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1395_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30084 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1396_
timestamp 1666464484
transform 1 0 29624 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29072 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1398_
timestamp 1666464484
transform 1 0 29716 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1399_
timestamp 1666464484
transform -1 0 32936 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1666464484
transform -1 0 25392 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1401_
timestamp 1666464484
transform 1 0 31372 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1666464484
transform -1 0 31280 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1403_
timestamp 1666464484
transform 1 0 30360 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1404_
timestamp 1666464484
transform -1 0 30912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1405_
timestamp 1666464484
transform -1 0 31096 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1406_
timestamp 1666464484
transform 1 0 24656 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1407_
timestamp 1666464484
transform 1 0 24748 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1408_
timestamp 1666464484
transform -1 0 25760 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1409_
timestamp 1666464484
transform 1 0 22264 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1410_
timestamp 1666464484
transform 1 0 23092 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1411_
timestamp 1666464484
transform -1 0 22724 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1412_
timestamp 1666464484
transform -1 0 21528 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1413_
timestamp 1666464484
transform -1 0 27140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1414_
timestamp 1666464484
transform 1 0 27140 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1415_
timestamp 1666464484
transform -1 0 26496 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1666464484
transform 1 0 30268 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1417_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29624 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1418_
timestamp 1666464484
transform -1 0 29256 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1419_
timestamp 1666464484
transform -1 0 26680 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1420_
timestamp 1666464484
transform -1 0 26128 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1421_
timestamp 1666464484
transform 1 0 25116 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 1666464484
transform -1 0 24840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1423_
timestamp 1666464484
transform -1 0 24564 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _1424_
timestamp 1666464484
transform 1 0 24932 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1425_
timestamp 1666464484
transform 1 0 25576 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1426_
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1427_
timestamp 1666464484
transform -1 0 26312 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1666464484
transform 1 0 30820 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1429_
timestamp 1666464484
transform 1 0 31372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1430_
timestamp 1666464484
transform 1 0 32292 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _1431_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1432_
timestamp 1666464484
transform -1 0 33856 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1433_
timestamp 1666464484
transform 1 0 32292 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1434_
timestamp 1666464484
transform 1 0 31832 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1435_
timestamp 1666464484
transform -1 0 33028 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1666464484
transform 1 0 33120 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1437_
timestamp 1666464484
transform 1 0 32476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1438_
timestamp 1666464484
transform 1 0 32660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1439_
timestamp 1666464484
transform -1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1440_
timestamp 1666464484
transform 1 0 29624 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _1441_
timestamp 1666464484
transform 1 0 32016 0 1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _1442_
timestamp 1666464484
transform 1 0 25116 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1443_
timestamp 1666464484
transform 1 0 24380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1444_
timestamp 1666464484
transform -1 0 25852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1445_
timestamp 1666464484
transform -1 0 21068 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1666464484
transform 1 0 20608 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1447_
timestamp 1666464484
transform 1 0 19136 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1448_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1449_
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _1450_
timestamp 1666464484
transform 1 0 32384 0 -1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1451_
timestamp 1666464484
transform -1 0 35144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1452_
timestamp 1666464484
transform -1 0 33488 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1453_
timestamp 1666464484
transform 1 0 32568 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1454_
timestamp 1666464484
transform -1 0 33028 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1455_
timestamp 1666464484
transform -1 0 27508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1456_
timestamp 1666464484
transform -1 0 26680 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1666464484
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1458_
timestamp 1666464484
transform -1 0 26680 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1459_
timestamp 1666464484
transform 1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1460_
timestamp 1666464484
transform -1 0 30360 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1461_
timestamp 1666464484
transform 1 0 30636 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 1666464484
transform -1 0 30912 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1463_
timestamp 1666464484
transform 1 0 31096 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1464_
timestamp 1666464484
transform 1 0 34868 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1465_
timestamp 1666464484
transform 1 0 33304 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1466_
timestamp 1666464484
transform 1 0 32936 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1467_
timestamp 1666464484
transform -1 0 33120 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1468_
timestamp 1666464484
transform 1 0 33212 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _1469_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33488 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1470_
timestamp 1666464484
transform -1 0 34132 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1471_
timestamp 1666464484
transform 1 0 34132 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1472_
timestamp 1666464484
transform 1 0 34776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1473_
timestamp 1666464484
transform 1 0 33948 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1474_
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1475_
timestamp 1666464484
transform 1 0 32752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1476_
timestamp 1666464484
transform -1 0 32936 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1477_
timestamp 1666464484
transform 1 0 36616 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1478_
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _1479_
timestamp 1666464484
transform 1 0 33856 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1480_
timestamp 1666464484
transform 1 0 35144 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1481_
timestamp 1666464484
transform 1 0 31280 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1482_
timestamp 1666464484
transform 1 0 27232 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1483_
timestamp 1666464484
transform 1 0 27508 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1484_
timestamp 1666464484
transform 1 0 27692 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1485_
timestamp 1666464484
transform 1 0 28428 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp 1666464484
transform 1 0 29716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1487_
timestamp 1666464484
transform 1 0 31096 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1488_
timestamp 1666464484
transform -1 0 30728 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1489_
timestamp 1666464484
transform 1 0 34868 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1490_
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1491_
timestamp 1666464484
transform -1 0 32752 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1492_
timestamp 1666464484
transform -1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1493_
timestamp 1666464484
transform 1 0 35512 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1494_
timestamp 1666464484
transform -1 0 36340 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1495_
timestamp 1666464484
transform -1 0 35880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1496_
timestamp 1666464484
transform -1 0 35696 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1497_
timestamp 1666464484
transform -1 0 36432 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1498_
timestamp 1666464484
transform -1 0 36064 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1499_
timestamp 1666464484
transform -1 0 36248 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1500_
timestamp 1666464484
transform 1 0 35696 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1501_
timestamp 1666464484
transform 1 0 35420 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1502_
timestamp 1666464484
transform -1 0 36524 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 1666464484
transform -1 0 35328 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1504_
timestamp 1666464484
transform 1 0 37444 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1505_
timestamp 1666464484
transform -1 0 25116 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1506_
timestamp 1666464484
transform 1 0 36340 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1507_
timestamp 1666464484
transform 1 0 37444 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1508_
timestamp 1666464484
transform -1 0 39008 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1509_
timestamp 1666464484
transform 1 0 38640 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1666464484
transform 1 0 40020 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1666464484
transform 1 0 39376 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1512_
timestamp 1666464484
transform 1 0 39560 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1513_
timestamp 1666464484
transform 1 0 28796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1514_
timestamp 1666464484
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1515_
timestamp 1666464484
transform -1 0 37076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1516_
timestamp 1666464484
transform 1 0 37444 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1517_
timestamp 1666464484
transform -1 0 38824 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1518_
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1519_
timestamp 1666464484
transform 1 0 37260 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1666464484
transform 1 0 37444 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1521_
timestamp 1666464484
transform 1 0 15456 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1522_
timestamp 1666464484
transform 1 0 16192 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1523_
timestamp 1666464484
transform -1 0 34960 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1524_
timestamp 1666464484
transform -1 0 42596 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1525_
timestamp 1666464484
transform 1 0 42596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1526_
timestamp 1666464484
transform 1 0 43976 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _1527_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 43424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1528_
timestamp 1666464484
transform 1 0 45172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1529_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 44620 0 -1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_4  _1530_
timestamp 1666464484
transform 1 0 45172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1531_
timestamp 1666464484
transform -1 0 44528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1532_
timestamp 1666464484
transform -1 0 43884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1533_
timestamp 1666464484
transform -1 0 45632 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _1534_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 45816 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1535_
timestamp 1666464484
transform -1 0 44068 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1536_
timestamp 1666464484
transform 1 0 43700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1537_
timestamp 1666464484
transform -1 0 41032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1538_
timestamp 1666464484
transform 1 0 43516 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1539_
timestamp 1666464484
transform -1 0 44344 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1540_
timestamp 1666464484
transform -1 0 39468 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1541_
timestamp 1666464484
transform -1 0 40480 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1542_
timestamp 1666464484
transform -1 0 42136 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1543_
timestamp 1666464484
transform 1 0 40020 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1544_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 44528 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1545_
timestamp 1666464484
transform 1 0 41952 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1546_
timestamp 1666464484
transform 1 0 37812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1547_
timestamp 1666464484
transform 1 0 39192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _1548_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38824 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1666464484
transform 1 0 39836 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1666464484
transform 1 0 40204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1551_
timestamp 1666464484
transform 1 0 38732 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1552_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 41216 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1553_
timestamp 1666464484
transform 1 0 37444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1666464484
transform 1 0 39008 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1555_
timestamp 1666464484
transform 1 0 39100 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 1666464484
transform 1 0 29624 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1557_
timestamp 1666464484
transform -1 0 30084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1558_
timestamp 1666464484
transform 1 0 39284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _1559_
timestamp 1666464484
transform -1 0 47012 0 -1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__a21bo_1  _1560_
timestamp 1666464484
transform -1 0 42872 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1561_
timestamp 1666464484
transform 1 0 41216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _1562_
timestamp 1666464484
transform -1 0 45540 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1563_
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1564_
timestamp 1666464484
transform 1 0 36432 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1565_
timestamp 1666464484
transform -1 0 45632 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _1566_
timestamp 1666464484
transform 1 0 42596 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1567_
timestamp 1666464484
transform 1 0 37628 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1568_
timestamp 1666464484
transform -1 0 45540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1569_
timestamp 1666464484
transform -1 0 43976 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1570_
timestamp 1666464484
transform -1 0 43884 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1571_
timestamp 1666464484
transform -1 0 43976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_2  _1572_
timestamp 1666464484
transform -1 0 45816 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1573_
timestamp 1666464484
transform 1 0 44712 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1574_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43608 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1575_
timestamp 1666464484
transform 1 0 36156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1576_
timestamp 1666464484
transform -1 0 39008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1577_
timestamp 1666464484
transform -1 0 37260 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1578_
timestamp 1666464484
transform 1 0 37444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1579_
timestamp 1666464484
transform -1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1580_
timestamp 1666464484
transform 1 0 35696 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1581_
timestamp 1666464484
transform 1 0 39468 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_4  _1582_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 45356 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1666464484
transform 1 0 34684 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1584_
timestamp 1666464484
transform -1 0 43792 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1585_
timestamp 1666464484
transform -1 0 36156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1586_
timestamp 1666464484
transform 1 0 35420 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _1587_
timestamp 1666464484
transform -1 0 35788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1588_
timestamp 1666464484
transform 1 0 38364 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1589_
timestamp 1666464484
transform 1 0 40020 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1590_
timestamp 1666464484
transform 1 0 31096 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1591_
timestamp 1666464484
transform 1 0 45724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1592_
timestamp 1666464484
transform -1 0 44804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37168 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1594_
timestamp 1666464484
transform 1 0 41032 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1595_
timestamp 1666464484
transform 1 0 46460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_2  _1596_
timestamp 1666464484
transform 1 0 45172 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _1597_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 39560 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1598_
timestamp 1666464484
transform -1 0 39008 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1599_
timestamp 1666464484
transform -1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1600_
timestamp 1666464484
transform 1 0 37904 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1601_
timestamp 1666464484
transform 1 0 35328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1602_
timestamp 1666464484
transform -1 0 35696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1603_
timestamp 1666464484
transform 1 0 41676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1604_
timestamp 1666464484
transform 1 0 42320 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1605_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 42964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1606_
timestamp 1666464484
transform 1 0 40112 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1607_
timestamp 1666464484
transform -1 0 43240 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1608_
timestamp 1666464484
transform 1 0 42412 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1609_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 41584 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1610_
timestamp 1666464484
transform 1 0 42872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1611_
timestamp 1666464484
transform -1 0 46092 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1612_
timestamp 1666464484
transform -1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1613_
timestamp 1666464484
transform -1 0 44528 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1614_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 43516 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1615_
timestamp 1666464484
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1616_
timestamp 1666464484
transform -1 0 34132 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1617_
timestamp 1666464484
transform 1 0 44344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _1618_
timestamp 1666464484
transform 1 0 44988 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1619_
timestamp 1666464484
transform 1 0 43884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1620_
timestamp 1666464484
transform 1 0 36432 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1621_
timestamp 1666464484
transform -1 0 36156 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1622_
timestamp 1666464484
transform 1 0 37444 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1623_
timestamp 1666464484
transform -1 0 36800 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1624_
timestamp 1666464484
transform -1 0 43056 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1625_
timestamp 1666464484
transform 1 0 43976 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1626_
timestamp 1666464484
transform 1 0 42964 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1627_
timestamp 1666464484
transform 1 0 41952 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1628_
timestamp 1666464484
transform -1 0 37812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1629_
timestamp 1666464484
transform -1 0 43976 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1630_
timestamp 1666464484
transform 1 0 45172 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1631_
timestamp 1666464484
transform 1 0 45172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1632_
timestamp 1666464484
transform -1 0 41492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1633_
timestamp 1666464484
transform -1 0 43148 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _1634_
timestamp 1666464484
transform 1 0 42320 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _1635_
timestamp 1666464484
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1636_
timestamp 1666464484
transform -1 0 37444 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1637_
timestamp 1666464484
transform 1 0 33672 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _1638_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33580 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1639_
timestamp 1666464484
transform 1 0 35512 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1640_
timestamp 1666464484
transform 1 0 41124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1641_
timestamp 1666464484
transform -1 0 36248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1642_
timestamp 1666464484
transform 1 0 38456 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1643_
timestamp 1666464484
transform -1 0 34408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1666464484
transform 1 0 43056 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1645_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34040 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1646_
timestamp 1666464484
transform 1 0 42872 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1647_
timestamp 1666464484
transform 1 0 34960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1648_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33856 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1649_
timestamp 1666464484
transform 1 0 37904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1650_
timestamp 1666464484
transform -1 0 38824 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1651_
timestamp 1666464484
transform 1 0 37720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1652_
timestamp 1666464484
transform -1 0 38272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1653_
timestamp 1666464484
transform -1 0 41124 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1654_
timestamp 1666464484
transform -1 0 41584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1655_
timestamp 1666464484
transform 1 0 40020 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1656_
timestamp 1666464484
transform 1 0 39192 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1657_
timestamp 1666464484
transform 1 0 37628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1658_
timestamp 1666464484
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1659_
timestamp 1666464484
transform 1 0 31556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1660_
timestamp 1666464484
transform 1 0 27784 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1661_
timestamp 1666464484
transform 1 0 27232 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1662_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29256 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1663_
timestamp 1666464484
transform 1 0 31096 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1664_
timestamp 1666464484
transform 1 0 39652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1665_
timestamp 1666464484
transform 1 0 42412 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1666_
timestamp 1666464484
transform 1 0 41308 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1667_
timestamp 1666464484
transform 1 0 45172 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1668_
timestamp 1666464484
transform -1 0 41032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 1666464484
transform -1 0 41952 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1670_
timestamp 1666464484
transform 1 0 40848 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _1671_
timestamp 1666464484
transform 1 0 40572 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__a311o_1  _1672_
timestamp 1666464484
transform 1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1673_
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1674_
timestamp 1666464484
transform -1 0 43976 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1675_
timestamp 1666464484
transform -1 0 35696 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1666464484
transform 1 0 44988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1677_
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1678_
timestamp 1666464484
transform 1 0 34776 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1679_
timestamp 1666464484
transform -1 0 31556 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1680_
timestamp 1666464484
transform -1 0 30728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1681_
timestamp 1666464484
transform -1 0 31648 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1682_
timestamp 1666464484
transform 1 0 32476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1683_
timestamp 1666464484
transform 1 0 32568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1684_
timestamp 1666464484
transform 1 0 33672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1685_
timestamp 1666464484
transform -1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp 1666464484
transform -1 0 35144 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1687_
timestamp 1666464484
transform -1 0 34408 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1688_
timestamp 1666464484
transform 1 0 34408 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1689_
timestamp 1666464484
transform -1 0 36524 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1690_
timestamp 1666464484
transform -1 0 36248 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1691_
timestamp 1666464484
transform -1 0 35788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1692_
timestamp 1666464484
transform 1 0 36248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1693_
timestamp 1666464484
transform 1 0 35420 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1694_
timestamp 1666464484
transform 1 0 35512 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1695_
timestamp 1666464484
transform -1 0 35144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1696_
timestamp 1666464484
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1697_
timestamp 1666464484
transform -1 0 34224 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1698_
timestamp 1666464484
transform 1 0 33396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1699_
timestamp 1666464484
transform 1 0 33212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1700_
timestamp 1666464484
transform -1 0 39560 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1701_
timestamp 1666464484
transform 1 0 38088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1702_
timestamp 1666464484
transform 1 0 35328 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1703_
timestamp 1666464484
transform 1 0 35788 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1704_
timestamp 1666464484
transform -1 0 38088 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1705_
timestamp 1666464484
transform -1 0 33948 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1706_
timestamp 1666464484
transform 1 0 31372 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _1707_
timestamp 1666464484
transform 1 0 34408 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1708_
timestamp 1666464484
transform 1 0 42964 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1709_
timestamp 1666464484
transform -1 0 42320 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1710_
timestamp 1666464484
transform -1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1711_
timestamp 1666464484
transform -1 0 42136 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1712_
timestamp 1666464484
transform 1 0 40572 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1713_
timestamp 1666464484
transform 1 0 40020 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1714_
timestamp 1666464484
transform 1 0 40664 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1715_
timestamp 1666464484
transform -1 0 41216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1716_
timestamp 1666464484
transform 1 0 40664 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1717_
timestamp 1666464484
transform 1 0 40112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1718_
timestamp 1666464484
transform 1 0 40020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1719_
timestamp 1666464484
transform 1 0 32108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1720_
timestamp 1666464484
transform -1 0 33580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1721_
timestamp 1666464484
transform -1 0 32752 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1722_
timestamp 1666464484
transform 1 0 36800 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _1723_
timestamp 1666464484
transform -1 0 44712 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1724_
timestamp 1666464484
transform 1 0 41768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1725_
timestamp 1666464484
transform 1 0 41308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1726_
timestamp 1666464484
transform -1 0 41216 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1727_
timestamp 1666464484
transform 1 0 39100 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1728_
timestamp 1666464484
transform -1 0 40204 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1729_
timestamp 1666464484
transform 1 0 45172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1730_
timestamp 1666464484
transform -1 0 41584 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1731_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 41308 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1732_
timestamp 1666464484
transform -1 0 36984 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1733_
timestamp 1666464484
transform 1 0 28428 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1734_
timestamp 1666464484
transform 1 0 28520 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1735_
timestamp 1666464484
transform 1 0 32568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1736_
timestamp 1666464484
transform -1 0 32936 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1737_
timestamp 1666464484
transform -1 0 30360 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1738_
timestamp 1666464484
transform -1 0 30360 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1739_
timestamp 1666464484
transform 1 0 29716 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1740_
timestamp 1666464484
transform 1 0 30452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1741_
timestamp 1666464484
transform 1 0 31004 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1742_
timestamp 1666464484
transform 1 0 31004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1743_
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1744_
timestamp 1666464484
transform 1 0 31188 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1745_
timestamp 1666464484
transform -1 0 29256 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1746_
timestamp 1666464484
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1747_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1748_
timestamp 1666464484
transform -1 0 38456 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1749_
timestamp 1666464484
transform -1 0 39652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1750_
timestamp 1666464484
transform 1 0 38180 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1751_
timestamp 1666464484
transform -1 0 40296 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1752_
timestamp 1666464484
transform -1 0 39560 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1753_
timestamp 1666464484
transform 1 0 37720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1754_
timestamp 1666464484
transform 1 0 37260 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1755_
timestamp 1666464484
transform -1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1756_
timestamp 1666464484
transform 1 0 32752 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1757_
timestamp 1666464484
transform -1 0 33028 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_2  _1758_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 38916 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _1759_
timestamp 1666464484
transform -1 0 27692 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1760_
timestamp 1666464484
transform -1 0 35328 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 1666464484
transform 1 0 34684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1762_
timestamp 1666464484
transform -1 0 34960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 1666464484
transform -1 0 39744 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1764_
timestamp 1666464484
transform 1 0 35144 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1765_
timestamp 1666464484
transform -1 0 44068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1766_
timestamp 1666464484
transform 1 0 38824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1767_
timestamp 1666464484
transform 1 0 34868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1768_
timestamp 1666464484
transform -1 0 27784 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1769_
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1770_
timestamp 1666464484
transform 1 0 31004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1771_
timestamp 1666464484
transform 1 0 31372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1772_
timestamp 1666464484
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1773_
timestamp 1666464484
transform -1 0 36616 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1774_
timestamp 1666464484
transform -1 0 36892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1775_
timestamp 1666464484
transform -1 0 32844 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1776_
timestamp 1666464484
transform -1 0 38456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1777_
timestamp 1666464484
transform 1 0 38824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1778_
timestamp 1666464484
transform 1 0 36800 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1779_
timestamp 1666464484
transform 1 0 30912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1780_
timestamp 1666464484
transform 1 0 31096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1781_
timestamp 1666464484
transform 1 0 30176 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1782_
timestamp 1666464484
transform 1 0 29256 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1783_
timestamp 1666464484
transform 1 0 27232 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1784_
timestamp 1666464484
transform 1 0 28336 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1785_
timestamp 1666464484
transform -1 0 29164 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _1786_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1787_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1788_
timestamp 1666464484
transform 1 0 28704 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _1789_
timestamp 1666464484
transform -1 0 27692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1790_
timestamp 1666464484
transform -1 0 28060 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1791_
timestamp 1666464484
transform -1 0 33856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1792_
timestamp 1666464484
transform -1 0 33948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1793_
timestamp 1666464484
transform 1 0 43148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1794_
timestamp 1666464484
transform 1 0 40572 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1795_
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp 1666464484
transform -1 0 31832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1797_
timestamp 1666464484
transform 1 0 32384 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1798_
timestamp 1666464484
transform -1 0 32752 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1799_
timestamp 1666464484
transform -1 0 32016 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1800_
timestamp 1666464484
transform -1 0 28152 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1801_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1802_
timestamp 1666464484
transform -1 0 39008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1803_
timestamp 1666464484
transform -1 0 40664 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1804_
timestamp 1666464484
transform -1 0 40296 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1805_
timestamp 1666464484
transform 1 0 38548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1806_
timestamp 1666464484
transform -1 0 26864 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1807_
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1666464484
transform 1 0 30176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1809_
timestamp 1666464484
transform -1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1810_
timestamp 1666464484
transform -1 0 25944 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1811_
timestamp 1666464484
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1812_
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1666464484
transform 1 0 26404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1814_
timestamp 1666464484
transform -1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1815_
timestamp 1666464484
transform -1 0 26404 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1816_
timestamp 1666464484
transform 1 0 25300 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1817_
timestamp 1666464484
transform -1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1818_
timestamp 1666464484
transform 1 0 37536 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1819_
timestamp 1666464484
transform 1 0 36340 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1820_
timestamp 1666464484
transform -1 0 35972 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1821_
timestamp 1666464484
transform -1 0 37812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1822_
timestamp 1666464484
transform 1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1823_
timestamp 1666464484
transform 1 0 36340 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1824_
timestamp 1666464484
transform 1 0 35604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1825_
timestamp 1666464484
transform 1 0 32476 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1826_
timestamp 1666464484
transform -1 0 33212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1827_
timestamp 1666464484
transform -1 0 31832 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1828_
timestamp 1666464484
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1829_
timestamp 1666464484
transform 1 0 28244 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1830_
timestamp 1666464484
transform 1 0 35328 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1831_
timestamp 1666464484
transform -1 0 35144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1832_
timestamp 1666464484
transform -1 0 34132 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1833_
timestamp 1666464484
transform 1 0 33304 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1834_
timestamp 1666464484
transform 1 0 32660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1835_
timestamp 1666464484
transform 1 0 27784 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1836_
timestamp 1666464484
transform -1 0 28060 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1837_
timestamp 1666464484
transform 1 0 39376 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1838_
timestamp 1666464484
transform 1 0 39928 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1839_
timestamp 1666464484
transform -1 0 37536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1840_
timestamp 1666464484
transform 1 0 41216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1841_
timestamp 1666464484
transform -1 0 40664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1842_
timestamp 1666464484
transform 1 0 40112 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1843_
timestamp 1666464484
transform 1 0 40020 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1844_
timestamp 1666464484
transform 1 0 38824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1845_
timestamp 1666464484
transform -1 0 30360 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1846_
timestamp 1666464484
transform -1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1847_
timestamp 1666464484
transform -1 0 27140 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1848_
timestamp 1666464484
transform 1 0 25484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1849_
timestamp 1666464484
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1850_
timestamp 1666464484
transform 1 0 25576 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1851_
timestamp 1666464484
transform -1 0 25208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1852_
timestamp 1666464484
transform 1 0 25024 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1853_
timestamp 1666464484
transform 1 0 26036 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1854_
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1666464484
transform -1 0 28520 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1856_
timestamp 1666464484
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1857_
timestamp 1666464484
transform 1 0 33212 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1858_
timestamp 1666464484
transform 1 0 33764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1859_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1860_
timestamp 1666464484
transform 1 0 32384 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1861_
timestamp 1666464484
transform -1 0 32844 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1862_
timestamp 1666464484
transform -1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1863_
timestamp 1666464484
transform 1 0 35788 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1864_
timestamp 1666464484
transform 1 0 35696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1865_
timestamp 1666464484
transform 1 0 35696 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1866_
timestamp 1666464484
transform -1 0 30176 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1867_
timestamp 1666464484
transform 1 0 28612 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1868_
timestamp 1666464484
transform -1 0 35604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1869_
timestamp 1666464484
transform -1 0 35512 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1870_
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1871_
timestamp 1666464484
transform -1 0 34684 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1872_
timestamp 1666464484
transform 1 0 33396 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1873_
timestamp 1666464484
transform 1 0 31556 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1874_
timestamp 1666464484
transform 1 0 32292 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1875_
timestamp 1666464484
transform 1 0 31096 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1876_
timestamp 1666464484
transform -1 0 30452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1877_
timestamp 1666464484
transform -1 0 30820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1878_
timestamp 1666464484
transform -1 0 30728 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1879_
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1880_
timestamp 1666464484
transform -1 0 26680 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1881_
timestamp 1666464484
transform -1 0 24564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1882_
timestamp 1666464484
transform 1 0 24932 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1883_
timestamp 1666464484
transform -1 0 25392 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1884_
timestamp 1666464484
transform -1 0 39284 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1885_
timestamp 1666464484
transform 1 0 35880 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1886_
timestamp 1666464484
transform -1 0 27876 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1887_
timestamp 1666464484
transform 1 0 27508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1888_
timestamp 1666464484
transform 1 0 26956 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _1889_
timestamp 1666464484
transform 1 0 37168 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1890_
timestamp 1666464484
transform 1 0 34132 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1891_
timestamp 1666464484
transform -1 0 34408 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1892_
timestamp 1666464484
transform -1 0 31464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1893_
timestamp 1666464484
transform -1 0 32292 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1894_
timestamp 1666464484
transform 1 0 30728 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1895_
timestamp 1666464484
transform -1 0 25852 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1896_
timestamp 1666464484
transform -1 0 32660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1897_
timestamp 1666464484
transform 1 0 44160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1898_
timestamp 1666464484
transform 1 0 42136 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1899_
timestamp 1666464484
transform 1 0 36432 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1900_
timestamp 1666464484
transform -1 0 43332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1901_
timestamp 1666464484
transform 1 0 31832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1902_
timestamp 1666464484
transform -1 0 30636 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1903_
timestamp 1666464484
transform 1 0 29716 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1904_
timestamp 1666464484
transform 1 0 22540 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1905_
timestamp 1666464484
transform 1 0 30084 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _1906_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1907_
timestamp 1666464484
transform -1 0 24012 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ba_1  _1908_
timestamp 1666464484
transform 1 0 24932 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1909_
timestamp 1666464484
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1910_
timestamp 1666464484
transform -1 0 23184 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1911_
timestamp 1666464484
transform -1 0 25392 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1912_
timestamp 1666464484
transform 1 0 22816 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1913_
timestamp 1666464484
transform 1 0 32292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1914_
timestamp 1666464484
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1915_
timestamp 1666464484
transform 1 0 33028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_2  _1916_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _1917_
timestamp 1666464484
transform 1 0 31280 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1918_
timestamp 1666464484
transform 1 0 29808 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1919_
timestamp 1666464484
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1920_
timestamp 1666464484
transform -1 0 25024 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1921_
timestamp 1666464484
transform 1 0 24196 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1922_
timestamp 1666464484
transform 1 0 37444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1923_
timestamp 1666464484
transform -1 0 33488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1924_
timestamp 1666464484
transform 1 0 32384 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1925_
timestamp 1666464484
transform 1 0 30268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1926_
timestamp 1666464484
transform 1 0 29256 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1927_
timestamp 1666464484
transform -1 0 28888 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1928_
timestamp 1666464484
transform 1 0 23092 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1929_
timestamp 1666464484
transform -1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1930_
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1931_
timestamp 1666464484
transform -1 0 23920 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1932_
timestamp 1666464484
transform 1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1933_
timestamp 1666464484
transform -1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1934_
timestamp 1666464484
transform -1 0 22356 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1666464484
transform 1 0 33580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1936_
timestamp 1666464484
transform -1 0 30728 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1937_
timestamp 1666464484
transform -1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1938_
timestamp 1666464484
transform 1 0 28612 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_2  _1939_
timestamp 1666464484
transform -1 0 29072 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1940_
timestamp 1666464484
transform 1 0 27968 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1941_
timestamp 1666464484
transform -1 0 27600 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1942_
timestamp 1666464484
transform 1 0 33672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1943_
timestamp 1666464484
transform 1 0 33120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1944_
timestamp 1666464484
transform -1 0 31188 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1945_
timestamp 1666464484
transform -1 0 30544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1946_
timestamp 1666464484
transform -1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1947_
timestamp 1666464484
transform 1 0 25852 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _1948_
timestamp 1666464484
transform -1 0 26588 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _1949_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24656 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _1950_
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_1  _1951_
timestamp 1666464484
transform -1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1952_
timestamp 1666464484
transform 1 0 23184 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1953_
timestamp 1666464484
transform -1 0 24840 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__or2b_1  _1954_
timestamp 1666464484
transform 1 0 25024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1955_
timestamp 1666464484
transform -1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1956_
timestamp 1666464484
transform 1 0 33856 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1957_
timestamp 1666464484
transform 1 0 29256 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1958_
timestamp 1666464484
transform -1 0 29072 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1959_
timestamp 1666464484
transform 1 0 28336 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1960_
timestamp 1666464484
transform -1 0 27416 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1961_
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1962_
timestamp 1666464484
transform -1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1963_
timestamp 1666464484
transform -1 0 24748 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 1666464484
transform -1 0 23920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1965_
timestamp 1666464484
transform -1 0 23644 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1966_
timestamp 1666464484
transform -1 0 23920 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1967_
timestamp 1666464484
transform 1 0 23368 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__nand4_1  _1968_
timestamp 1666464484
transform 1 0 23368 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1969_
timestamp 1666464484
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1970_
timestamp 1666464484
transform -1 0 27876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1971_
timestamp 1666464484
transform 1 0 25852 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1972_
timestamp 1666464484
transform -1 0 26312 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1973_
timestamp 1666464484
transform -1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _1974_
timestamp 1666464484
transform 1 0 37536 0 1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1975_
timestamp 1666464484
transform 1 0 28152 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1976_
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1977_
timestamp 1666464484
transform 1 0 32660 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1978_
timestamp 1666464484
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1979_
timestamp 1666464484
transform 1 0 34224 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1980_
timestamp 1666464484
transform -1 0 34316 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1981_
timestamp 1666464484
transform 1 0 33580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1982_
timestamp 1666464484
transform 1 0 33672 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1983_
timestamp 1666464484
transform 1 0 36156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1984_
timestamp 1666464484
transform 1 0 35144 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1985_
timestamp 1666464484
transform 1 0 35052 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1986_
timestamp 1666464484
transform -1 0 35880 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1987_
timestamp 1666464484
transform -1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1988_
timestamp 1666464484
transform 1 0 33856 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1989_
timestamp 1666464484
transform 1 0 34868 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1990_
timestamp 1666464484
transform -1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1991_
timestamp 1666464484
transform -1 0 35512 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1992_
timestamp 1666464484
transform -1 0 34408 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1993_
timestamp 1666464484
transform -1 0 35328 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1994_
timestamp 1666464484
transform -1 0 35420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1995_
timestamp 1666464484
transform 1 0 35788 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1996_
timestamp 1666464484
transform 1 0 33856 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1997_
timestamp 1666464484
transform 1 0 33856 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1998_
timestamp 1666464484
transform -1 0 35328 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1999_
timestamp 1666464484
transform 1 0 34684 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2000_
timestamp 1666464484
transform 1 0 33764 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2001_
timestamp 1666464484
transform -1 0 34132 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2002_
timestamp 1666464484
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2003_
timestamp 1666464484
transform -1 0 34408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2004_
timestamp 1666464484
transform 1 0 33948 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2005_
timestamp 1666464484
transform -1 0 35604 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2006_
timestamp 1666464484
transform -1 0 34132 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2007_
timestamp 1666464484
transform -1 0 33028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2008_
timestamp 1666464484
transform -1 0 28152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2009_
timestamp 1666464484
transform -1 0 27324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2010_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31464 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2011_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29256 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2012_
timestamp 1666464484
transform 1 0 27416 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2013_
timestamp 1666464484
transform 1 0 29164 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2014_
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2015_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31832 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2016_
timestamp 1666464484
transform 1 0 29716 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dlxtn_1  _2017_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _2018_
timestamp 1666464484
transform -1 0 33488 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2019_
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2020_
timestamp 1666464484
transform 1 0 35880 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2021_
timestamp 1666464484
transform -1 0 33396 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2022_
timestamp 1666464484
transform 1 0 35880 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2023_
timestamp 1666464484
transform 1 0 35236 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2024_
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2025_
timestamp 1666464484
transform 1 0 24564 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dlxtn_1  _2026_
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_4  _2027_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35696 0 1 39168
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_1  _2028_
timestamp 1666464484
transform 1 0 33580 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2029_
timestamp 1666464484
transform 1 0 35144 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_4  _2030_
timestamp 1666464484
transform 1 0 34592 0 -1 36992
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_4  _2031_
timestamp 1666464484
transform 1 0 34776 0 -1 35904
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _2032_
timestamp 1666464484
transform 1 0 33764 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2033_
timestamp 1666464484
transform -1 0 24196 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2034_
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2035_
timestamp 1666464484
transform 1 0 28428 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout44
timestamp 1666464484
transform 1 0 33672 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1666464484
transform -1 0 38824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1666464484
transform -1 0 24104 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1666464484
transform 1 0 30912 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1666464484
transform 1 0 27876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1666464484
transform -1 0 36340 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36156 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 30360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1666464484
transform 1 0 2668 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1666464484
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 58420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1666464484
transform -1 0 6072 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 58052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform -1 0 1932 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform 1 0 58052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform 1 0 46460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform 1 0 58052 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1666464484
transform -1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1666464484
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1666464484
transform -1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1666464484
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1666464484
transform 1 0 35512 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1666464484
transform 1 0 52900 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform 1 0 58052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform 1 0 58052 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform 1 0 14260 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform -1 0 9476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform 1 0 49036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform 1 0 41308 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform -1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform 1 0 58052 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1666464484
transform 1 0 58052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1666464484
transform -1 0 19780 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1666464484
transform -1 0 24932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1666464484
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1666464484
transform -1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1666464484
transform -1 0 1932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1666464484
transform 1 0 58052 0 -1 29376
box -38 -48 406 592
<< labels >>
flabel metal2 s 30286 59200 30342 59800 0 FreeSans 224 90 0 0 ACK
port 0 nsew signal input
flabel metal2 s 2594 59200 2650 59800 0 FreeSans 224 90 0 0 Bit_In
port 1 nsew signal input
flabel metal2 s 43810 200 43866 800 0 FreeSans 224 90 0 0 EN
port 2 nsew signal input
flabel metal3 s 59200 5448 59800 5568 0 FreeSans 480 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal3 s 200 46248 800 46368 0 FreeSans 480 0 0 0 I[10]
port 4 nsew signal tristate
flabel metal2 s 59910 200 59966 800 0 FreeSans 224 90 0 0 I[11]
port 5 nsew signal tristate
flabel metal2 s 54758 200 54814 800 0 FreeSans 224 90 0 0 I[12]
port 6 nsew signal tristate
flabel metal3 s 59200 40128 59800 40248 0 FreeSans 480 0 0 0 I[1]
port 7 nsew signal tristate
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 I[2]
port 8 nsew signal tristate
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 I[3]
port 9 nsew signal tristate
flabel metal2 s 46386 59200 46442 59800 0 FreeSans 224 90 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 45568 59800 45688 0 FreeSans 480 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 I[7]
port 13 nsew signal tristate
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 I[8]
port 14 nsew signal tristate
flabel metal3 s 200 40128 800 40248 0 FreeSans 480 0 0 0 I[9]
port 15 nsew signal tristate
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 Q[0]
port 16 nsew signal tristate
flabel metal2 s 35438 59200 35494 59800 0 FreeSans 224 90 0 0 Q[10]
port 17 nsew signal tristate
flabel metal2 s 52182 59200 52238 59800 0 FreeSans 224 90 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 17008 59800 17128 0 FreeSans 480 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal3 s 59200 51688 59800 51808 0 FreeSans 480 0 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 13542 59200 13598 59800 0 FreeSans 224 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal3 s 59200 34008 59800 34128 0 FreeSans 480 0 0 0 Q[5]
port 24 nsew signal tristate
flabel metal2 s 8390 59200 8446 59800 0 FreeSans 224 90 0 0 Q[6]
port 25 nsew signal tristate
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 Q[7]
port 26 nsew signal tristate
flabel metal2 s 48962 200 49018 800 0 FreeSans 224 90 0 0 Q[8]
port 27 nsew signal tristate
flabel metal2 s 41234 59200 41290 59800 0 FreeSans 224 90 0 0 Q[9]
port 28 nsew signal tristate
flabel metal3 s 59200 10888 59800 11008 0 FreeSans 480 0 0 0 REQ_SAMPLE
port 29 nsew signal input
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 RST
port 30 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 addI[0]
port 31 nsew signal tristate
flabel metal3 s 200 51688 800 51808 0 FreeSans 480 0 0 0 addI[1]
port 32 nsew signal tristate
flabel metal3 s 59200 22448 59800 22568 0 FreeSans 480 0 0 0 addI[2]
port 33 nsew signal tristate
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 addI[3]
port 34 nsew signal tristate
flabel metal3 s 59200 57128 59800 57248 0 FreeSans 480 0 0 0 addI[4]
port 35 nsew signal tristate
flabel metal2 s 57334 59200 57390 59800 0 FreeSans 224 90 0 0 addI[5]
port 36 nsew signal tristate
flabel metal2 s 19338 59200 19394 59800 0 FreeSans 224 90 0 0 addQ[0]
port 37 nsew signal tristate
flabel metal2 s 24490 59200 24546 59800 0 FreeSans 224 90 0 0 addQ[1]
port 38 nsew signal tristate
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 addQ[2]
port 39 nsew signal tristate
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 addQ[3]
port 40 nsew signal tristate
flabel metal3 s 200 57808 800 57928 0 FreeSans 480 0 0 0 addQ[4]
port 41 nsew signal tristate
flabel metal3 s 59200 28568 59800 28688 0 FreeSans 480 0 0 0 addQ[5]
port 42 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 30406 57494 30406 57494 0 ACK
rlabel metal1 2714 57494 2714 57494 0 Bit_In
rlabel metal1 43884 2414 43884 2414 0 EN
rlabel via2 58282 5525 58282 5525 0 I[0]
rlabel metal3 1188 46308 1188 46308 0 I[10]
rlabel metal2 59938 1520 59938 1520 0 I[11]
rlabel metal2 54786 823 54786 823 0 I[12]
rlabel metal2 58282 40273 58282 40273 0 I[1]
rlabel metal2 21942 1520 21942 1520 0 I[2]
rlabel metal2 32890 1520 32890 1520 0 I[3]
rlabel metal1 46552 57562 46552 57562 0 I[4]
rlabel metal3 1188 23188 1188 23188 0 I[5]
rlabel metal2 58282 45713 58282 45713 0 I[6]
rlabel metal3 1188 34748 1188 34748 0 I[7]
rlabel metal2 10994 1520 10994 1520 0 I[8]
rlabel metal3 1188 40188 1188 40188 0 I[9]
rlabel metal3 1188 17068 1188 17068 0 Q[0]
rlabel metal1 35604 57562 35604 57562 0 Q[10]
rlabel metal1 52670 57562 52670 57562 0 Q[11]
rlabel via2 58282 17051 58282 17051 0 Q[12]
rlabel via2 58282 51765 58282 51765 0 Q[1]
rlabel metal1 14030 57562 14030 57562 0 Q[2]
rlabel metal2 46 1520 46 1520 0 Q[3]
rlabel metal3 1188 11628 1188 11628 0 Q[4]
rlabel metal1 58098 34714 58098 34714 0 Q[5]
rlabel metal1 8832 57562 8832 57562 0 Q[6]
rlabel metal3 1188 5508 1188 5508 0 Q[7]
rlabel metal2 48990 1520 48990 1520 0 Q[8]
rlabel metal1 41492 57562 41492 57562 0 Q[9]
rlabel metal2 58282 10999 58282 10999 0 REQ_SAMPLE
rlabel metal1 5796 2414 5796 2414 0 RST
rlabel metal2 26174 12036 26174 12036 0 _0000_
rlabel metal2 25714 12036 25714 12036 0 _0001_
rlabel metal2 26910 30090 26910 30090 0 _0002_
rlabel metal1 26634 29716 26634 29716 0 _0003_
rlabel metal1 27140 10642 27140 10642 0 _0004_
rlabel metal1 33166 29478 33166 29478 0 _0005_
rlabel metal2 31142 28254 31142 28254 0 _0006_
rlabel metal1 29532 32946 29532 32946 0 _0007_
rlabel metal2 33166 25500 33166 25500 0 _0008_
rlabel metal1 35926 26010 35926 26010 0 _0009_
rlabel via1 35650 24667 35650 24667 0 _0010_
rlabel metal1 33488 24242 33488 24242 0 _0011_
rlabel metal1 35824 27642 35824 27642 0 _0012_
rlabel metal1 35466 27098 35466 27098 0 _0013_
rlabel metal2 36110 39644 36110 39644 0 _0014_
rlabel metal2 33902 39508 33902 39508 0 _0015_
rlabel metal2 35374 38114 35374 38114 0 _0016_
rlabel metal2 35006 36924 35006 36924 0 _0017_
rlabel metal2 35190 35836 35190 35836 0 _0018_
rlabel metal1 33534 29750 33534 29750 0 _0019_
rlabel metal1 27324 9146 27324 9146 0 _0020_
rlabel metal1 30958 12240 30958 12240 0 _0021_
rlabel metal1 23598 21964 23598 21964 0 _0022_
rlabel metal2 24794 22780 24794 22780 0 _0023_
rlabel metal1 21942 23052 21942 23052 0 _0024_
rlabel metal1 24426 19822 24426 19822 0 _0025_
rlabel metal1 23460 20026 23460 20026 0 _0026_
rlabel metal2 32430 18666 32430 18666 0 _0027_
rlabel metal2 33350 16014 33350 16014 0 _0028_
rlabel metal1 31970 16490 31970 16490 0 _0029_
rlabel metal2 24610 17170 24610 17170 0 _0030_
rlabel metal2 31050 21828 31050 21828 0 _0031_
rlabel metal2 30498 21658 30498 21658 0 _0032_
rlabel metal1 25024 18734 25024 18734 0 _0033_
rlabel metal1 24518 18258 24518 18258 0 _0034_
rlabel via1 24242 18598 24242 18598 0 _0035_
rlabel metal1 23828 18734 23828 18734 0 _0036_
rlabel metal1 32614 19414 32614 19414 0 _0037_
rlabel metal2 33258 18904 33258 18904 0 _0038_
rlabel metal1 30360 19346 30360 19346 0 _0039_
rlabel metal1 29762 19312 29762 19312 0 _0040_
rlabel metal1 28980 19346 28980 19346 0 _0041_
rlabel metal2 25254 11934 25254 11934 0 _0042_
rlabel metal1 25944 18802 25944 18802 0 _0043_
rlabel metal2 23506 19108 23506 19108 0 _0044_
rlabel metal2 23874 20196 23874 20196 0 _0045_
rlabel metal1 23736 20910 23736 20910 0 _0046_
rlabel metal1 22816 21930 22816 21930 0 _0047_
rlabel metal1 23046 22950 23046 22950 0 _0048_
rlabel metal2 21758 22474 21758 22474 0 _0049_
rlabel metal1 32683 15402 32683 15402 0 _0050_
rlabel metal1 28566 15028 28566 15028 0 _0051_
rlabel metal1 28842 14926 28842 14926 0 _0052_
rlabel metal2 28934 18156 28934 18156 0 _0053_
rlabel metal1 27370 14960 27370 14960 0 _0054_
rlabel metal2 28014 14790 28014 14790 0 _0055_
rlabel metal2 27186 14110 27186 14110 0 _0056_
rlabel metal1 33764 16082 33764 16082 0 _0057_
rlabel metal1 27278 15504 27278 15504 0 _0058_
rlabel metal2 30774 13056 30774 13056 0 _0059_
rlabel metal1 26680 13294 26680 13294 0 _0060_
rlabel metal1 26726 14994 26726 14994 0 _0061_
rlabel metal2 21942 37128 21942 37128 0 _0062_
rlabel metal2 25622 14926 25622 14926 0 _0063_
rlabel metal2 23966 15198 23966 15198 0 _0064_
rlabel metal2 24334 16558 24334 16558 0 _0065_
rlabel metal2 24242 16014 24242 16014 0 _0066_
rlabel metal2 23782 21794 23782 21794 0 _0067_
rlabel metal1 23828 17170 23828 17170 0 _0068_
rlabel viali 25620 13906 25620 13906 0 _0069_
rlabel metal2 29670 14416 29670 14416 0 _0070_
rlabel metal2 33902 13974 33902 13974 0 _0071_
rlabel metal1 22908 46546 22908 46546 0 _0072_
rlabel metal1 29072 13906 29072 13906 0 _0073_
rlabel metal1 28750 13498 28750 13498 0 _0074_
rlabel metal1 27876 13906 27876 13906 0 _0075_
rlabel metal1 25346 13872 25346 13872 0 _0076_
rlabel metal2 24426 13600 24426 13600 0 _0077_
rlabel metal1 24702 13906 24702 13906 0 _0078_
rlabel metal2 24334 13328 24334 13328 0 _0079_
rlabel metal1 23644 14042 23644 14042 0 _0080_
rlabel metal1 23598 13906 23598 13906 0 _0081_
rlabel metal2 23874 13260 23874 13260 0 _0082_
rlabel metal1 21390 44812 21390 44812 0 _0083_
rlabel metal1 24978 13192 24978 13192 0 _0084_
rlabel metal1 24794 13158 24794 13158 0 _0085_
rlabel metal1 26174 13294 26174 13294 0 _0086_
rlabel metal1 24978 13294 24978 13294 0 _0087_
rlabel metal2 25898 13124 25898 13124 0 _0088_
rlabel metal1 28842 28560 28842 28560 0 _0089_
rlabel metal2 33626 41684 33626 41684 0 _0090_
rlabel metal2 33258 26554 33258 26554 0 _0091_
rlabel metal2 33810 35071 33810 35071 0 _0092_
rlabel metal1 33810 25908 33810 25908 0 _0093_
rlabel metal1 33764 25466 33764 25466 0 _0094_
rlabel metal1 35190 36176 35190 36176 0 _0095_
rlabel metal1 35834 25942 35834 25942 0 _0096_
rlabel metal2 35558 24922 35558 24922 0 _0097_
rlabel metal1 28290 36754 28290 36754 0 _0098_
rlabel metal2 34362 24582 34362 24582 0 _0099_
rlabel metal1 35328 27370 35328 27370 0 _0100_
rlabel metal2 34822 27302 34822 27302 0 _0101_
rlabel metal1 34914 26996 34914 26996 0 _0102_
rlabel metal2 34730 27132 34730 27132 0 _0103_
rlabel metal1 34316 37978 34316 37978 0 _0104_
rlabel metal1 24978 47464 24978 47464 0 _0105_
rlabel metal2 34730 38352 34730 38352 0 _0106_
rlabel metal1 34178 37128 34178 37128 0 _0107_
rlabel metal2 34086 36924 34086 36924 0 _0108_
rlabel metal1 34086 36006 34086 36006 0 _0109_
rlabel metal1 34638 35802 34638 35802 0 _0110_
rlabel metal1 33304 34442 33304 34442 0 _0111_
rlabel metal1 33258 44234 33258 44234 0 _0112_
rlabel metal1 27600 8942 27600 8942 0 _0113_
rlabel metal1 30774 45458 30774 45458 0 _0114_
rlabel metal1 31004 40562 31004 40562 0 _0115_
rlabel metal1 31004 36346 31004 36346 0 _0116_
rlabel metal1 28750 35666 28750 35666 0 _0117_
rlabel metal1 29762 41174 29762 41174 0 _0118_
rlabel metal1 29624 41106 29624 41106 0 _0119_
rlabel metal1 29348 41106 29348 41106 0 _0120_
rlabel metal1 32798 40426 32798 40426 0 _0121_
rlabel metal1 28934 40018 28934 40018 0 _0122_
rlabel metal1 28520 37230 28520 37230 0 _0123_
rlabel metal1 30567 37842 30567 37842 0 _0124_
rlabel metal1 29992 35734 29992 35734 0 _0125_
rlabel metal2 35282 35904 35282 35904 0 _0126_
rlabel metal2 27462 11730 27462 11730 0 _0127_
rlabel metal1 30682 26554 30682 26554 0 _0128_
rlabel metal1 29256 12070 29256 12070 0 _0129_
rlabel metal1 27508 11866 27508 11866 0 _0130_
rlabel metal1 26772 11730 26772 11730 0 _0131_
rlabel via2 26266 30379 26266 30379 0 _0132_
rlabel metal1 20240 32742 20240 32742 0 _0133_
rlabel metal1 27186 30124 27186 30124 0 _0134_
rlabel metal1 26542 30362 26542 30362 0 _0135_
rlabel metal1 27600 27438 27600 27438 0 _0136_
rlabel metal2 25530 11900 25530 11900 0 _0137_
rlabel metal1 26588 29274 26588 29274 0 _0138_
rlabel metal2 32430 43554 32430 43554 0 _0139_
rlabel metal2 27462 42160 27462 42160 0 _0140_
rlabel metal2 33350 46784 33350 46784 0 _0141_
rlabel metal1 34546 42670 34546 42670 0 _0142_
rlabel via2 33718 41123 33718 41123 0 _0143_
rlabel metal1 26772 37230 26772 37230 0 _0144_
rlabel metal1 26266 35088 26266 35088 0 _0145_
rlabel via2 29026 40035 29026 40035 0 _0146_
rlabel metal1 32568 40494 32568 40494 0 _0147_
rlabel metal1 31878 40460 31878 40460 0 _0148_
rlabel metal1 32936 46614 32936 46614 0 _0149_
rlabel metal2 26634 45662 26634 45662 0 _0150_
rlabel metal1 26588 38726 26588 38726 0 _0151_
rlabel metal1 25070 38964 25070 38964 0 _0152_
rlabel metal1 32522 36584 32522 36584 0 _0153_
rlabel metal1 25852 38930 25852 38930 0 _0154_
rlabel metal1 33902 37740 33902 37740 0 _0155_
rlabel metal1 32890 39508 32890 39508 0 _0156_
rlabel metal1 27278 38726 27278 38726 0 _0157_
rlabel metal2 26082 38522 26082 38522 0 _0158_
rlabel metal1 21436 38318 21436 38318 0 _0159_
rlabel metal2 17526 36924 17526 36924 0 _0160_
rlabel metal2 28934 36856 28934 36856 0 _0161_
rlabel metal1 33442 41480 33442 41480 0 _0162_
rlabel metal1 34730 40494 34730 40494 0 _0163_
rlabel via2 21758 40477 21758 40477 0 _0164_
rlabel metal2 32706 41004 32706 41004 0 _0165_
rlabel metal1 22034 40528 22034 40528 0 _0166_
rlabel metal1 20009 40494 20009 40494 0 _0167_
rlabel metal1 19872 40086 19872 40086 0 _0168_
rlabel metal1 20470 37876 20470 37876 0 _0169_
rlabel via1 19914 40154 19914 40154 0 _0170_
rlabel metal1 27462 37876 27462 37876 0 _0171_
rlabel metal1 23046 40086 23046 40086 0 _0172_
rlabel metal2 24794 40868 24794 40868 0 _0173_
rlabel metal2 21206 40902 21206 40902 0 _0174_
rlabel metal1 25898 41718 25898 41718 0 _0175_
rlabel metal1 28750 43758 28750 43758 0 _0176_
rlabel metal1 27462 44336 27462 44336 0 _0177_
rlabel metal1 26848 43350 26848 43350 0 _0178_
rlabel metal2 20746 42789 20746 42789 0 _0179_
rlabel metal1 20240 40698 20240 40698 0 _0180_
rlabel metal2 18814 38556 18814 38556 0 _0181_
rlabel viali 23690 43755 23690 43755 0 _0182_
rlabel metal1 24748 37842 24748 37842 0 _0183_
rlabel metal2 24150 36992 24150 36992 0 _0184_
rlabel metal2 24242 37196 24242 37196 0 _0185_
rlabel metal1 23230 40460 23230 40460 0 _0186_
rlabel metal1 24012 36754 24012 36754 0 _0187_
rlabel metal2 21574 36652 21574 36652 0 _0188_
rlabel metal1 22402 38930 22402 38930 0 _0189_
rlabel metal2 21298 46818 21298 46818 0 _0190_
rlabel metal2 31786 47396 31786 47396 0 _0191_
rlabel via3 22195 39916 22195 39916 0 _0192_
rlabel metal2 25208 39950 25208 39950 0 _0193_
rlabel metal2 25806 44302 25806 44302 0 _0194_
rlabel metal3 24127 39780 24127 39780 0 _0195_
rlabel metal1 21482 37230 21482 37230 0 _0196_
rlabel metal2 19642 36550 19642 36550 0 _0197_
rlabel metal1 19366 35564 19366 35564 0 _0198_
rlabel metal1 19228 36686 19228 36686 0 _0199_
rlabel metal1 17802 36652 17802 36652 0 _0200_
rlabel metal2 20562 36618 20562 36618 0 _0201_
rlabel metal2 18722 39984 18722 39984 0 _0202_
rlabel metal1 28106 41582 28106 41582 0 _0203_
rlabel metal1 25116 42194 25116 42194 0 _0204_
rlabel metal1 32338 38930 32338 38930 0 _0205_
rlabel metal1 22402 40970 22402 40970 0 _0206_
rlabel metal1 20746 40970 20746 40970 0 _0207_
rlabel metal2 28474 46988 28474 46988 0 _0208_
rlabel metal1 20838 42058 20838 42058 0 _0209_
rlabel via1 23965 43282 23965 43282 0 _0210_
rlabel metal1 20378 42160 20378 42160 0 _0211_
rlabel metal1 19780 41990 19780 41990 0 _0212_
rlabel metal1 21528 41038 21528 41038 0 _0213_
rlabel metal1 21344 40970 21344 40970 0 _0214_
rlabel metal2 20746 39066 20746 39066 0 _0215_
rlabel metal1 20562 41106 20562 41106 0 _0216_
rlabel via1 20746 36771 20746 36771 0 _0217_
rlabel metal2 19458 35734 19458 35734 0 _0218_
rlabel metal2 19550 35462 19550 35462 0 _0219_
rlabel metal1 18170 35666 18170 35666 0 _0220_
rlabel metal1 20194 43656 20194 43656 0 _0221_
rlabel metal1 22310 44846 22310 44846 0 _0222_
rlabel metal1 20102 43792 20102 43792 0 _0223_
rlabel metal1 23690 45798 23690 45798 0 _0224_
rlabel metal2 21206 44268 21206 44268 0 _0225_
rlabel metal1 20654 43146 20654 43146 0 _0226_
rlabel metal2 22218 44064 22218 44064 0 _0227_
rlabel metal1 23690 41106 23690 41106 0 _0228_
rlabel metal1 20792 43758 20792 43758 0 _0229_
rlabel metal1 18354 35054 18354 35054 0 _0230_
rlabel metal2 18262 34918 18262 34918 0 _0231_
rlabel metal1 17204 35054 17204 35054 0 _0232_
rlabel metal1 16284 35122 16284 35122 0 _0233_
rlabel metal2 16146 36278 16146 36278 0 _0234_
rlabel metal2 17250 38624 17250 38624 0 _0235_
rlabel metal1 21252 37978 21252 37978 0 _0236_
rlabel metal1 32177 38522 32177 38522 0 _0237_
rlabel metal1 27646 37162 27646 37162 0 _0238_
rlabel metal1 26496 37842 26496 37842 0 _0239_
rlabel metal1 29854 45934 29854 45934 0 _0240_
rlabel metal2 30498 40715 30498 40715 0 _0241_
rlabel metal1 26266 44404 26266 44404 0 _0242_
rlabel metal1 29624 43894 29624 43894 0 _0243_
rlabel metal1 30958 42874 30958 42874 0 _0244_
rlabel metal2 26174 37961 26174 37961 0 _0245_
rlabel metal1 16330 38284 16330 38284 0 _0246_
rlabel metal1 16146 38964 16146 38964 0 _0247_
rlabel metal2 16606 38556 16606 38556 0 _0248_
rlabel metal2 16330 37502 16330 37502 0 _0249_
rlabel via1 15594 35802 15594 35802 0 _0250_
rlabel metal1 30958 39066 30958 39066 0 _0251_
rlabel metal1 29210 38386 29210 38386 0 _0252_
rlabel via1 22864 37230 22864 37230 0 _0253_
rlabel metal1 29716 46002 29716 46002 0 _0254_
rlabel metal2 31786 37468 31786 37468 0 _0255_
rlabel metal1 23092 37162 23092 37162 0 _0256_
rlabel metal1 20470 38964 20470 38964 0 _0257_
rlabel via1 22494 37230 22494 37230 0 _0258_
rlabel metal1 20470 36720 20470 36720 0 _0259_
rlabel metal2 21022 35020 21022 35020 0 _0260_
rlabel metal1 27094 31926 27094 31926 0 _0261_
rlabel metal1 27140 31450 27140 31450 0 _0262_
rlabel metal2 27830 31144 27830 31144 0 _0263_
rlabel metal1 21758 31722 21758 31722 0 _0264_
rlabel metal1 20792 33490 20792 33490 0 _0265_
rlabel metal2 27002 32980 27002 32980 0 _0266_
rlabel metal1 29992 42874 29992 42874 0 _0267_
rlabel metal1 21068 41990 21068 41990 0 _0268_
rlabel metal1 23276 38318 23276 38318 0 _0269_
rlabel metal1 23230 37672 23230 37672 0 _0270_
rlabel metal1 30406 38760 30406 38760 0 _0271_
rlabel metal2 22494 43996 22494 43996 0 _0272_
rlabel metal1 24104 43282 24104 43282 0 _0273_
rlabel metal1 22448 43078 22448 43078 0 _0274_
rlabel metal1 22770 34714 22770 34714 0 _0275_
rlabel metal2 23690 35836 23690 35836 0 _0276_
rlabel via1 23048 35666 23048 35666 0 _0277_
rlabel metal1 22356 45594 22356 45594 0 _0278_
rlabel metal1 24196 43758 24196 43758 0 _0279_
rlabel metal1 22770 45050 22770 45050 0 _0280_
rlabel metal2 22862 35785 22862 35785 0 _0281_
rlabel metal2 27094 40732 27094 40732 0 _0282_
rlabel metal1 25576 39814 25576 39814 0 _0283_
rlabel metal1 23598 34612 23598 34612 0 _0284_
rlabel metal1 21896 33422 21896 33422 0 _0285_
rlabel metal2 15686 33150 15686 33150 0 _0286_
rlabel metal2 17434 33490 17434 33490 0 _0287_
rlabel metal1 27920 42194 27920 42194 0 _0288_
rlabel metal1 29118 42738 29118 42738 0 _0289_
rlabel metal2 21390 39457 21390 39457 0 _0290_
rlabel metal1 20746 39372 20746 39372 0 _0291_
rlabel via2 23414 39253 23414 39253 0 _0292_
rlabel metal1 20240 39066 20240 39066 0 _0293_
rlabel metal1 19964 33490 19964 33490 0 _0294_
rlabel metal1 15594 33014 15594 33014 0 _0295_
rlabel metal1 15364 33422 15364 33422 0 _0296_
rlabel metal1 18078 39066 18078 39066 0 _0297_
rlabel metal2 32522 38080 32522 38080 0 _0298_
rlabel metal1 25530 43418 25530 43418 0 _0299_
rlabel metal1 25806 37196 25806 37196 0 _0300_
rlabel metal2 27186 43962 27186 43962 0 _0301_
rlabel metal1 26956 43826 26956 43826 0 _0302_
rlabel metal1 29716 35190 29716 35190 0 _0303_
rlabel metal2 28290 43452 28290 43452 0 _0304_
rlabel metal1 26496 43758 26496 43758 0 _0305_
rlabel metal1 19542 38182 19542 38182 0 _0306_
rlabel metal2 17710 38012 17710 38012 0 _0307_
rlabel metal1 18078 38522 18078 38522 0 _0308_
rlabel metal1 16146 33490 16146 33490 0 _0309_
rlabel metal1 15870 34918 15870 34918 0 _0310_
rlabel metal2 14950 35326 14950 35326 0 _0311_
rlabel metal1 15318 35666 15318 35666 0 _0312_
rlabel metal1 18032 36142 18032 36142 0 _0313_
rlabel metal1 16698 37298 16698 37298 0 _0314_
rlabel metal2 15594 36958 15594 36958 0 _0315_
rlabel metal1 15824 37162 15824 37162 0 _0316_
rlabel metal1 14352 35258 14352 35258 0 _0317_
rlabel metal1 14306 35632 14306 35632 0 _0318_
rlabel metal1 16100 31314 16100 31314 0 _0319_
rlabel metal1 16008 30906 16008 30906 0 _0320_
rlabel metal2 21758 34748 21758 34748 0 _0321_
rlabel metal2 21114 34714 21114 34714 0 _0322_
rlabel metal2 21758 33116 21758 33116 0 _0323_
rlabel metal1 28244 37434 28244 37434 0 _0324_
rlabel metal1 27278 35598 27278 35598 0 _0325_
rlabel metal1 24978 34612 24978 34612 0 _0326_
rlabel metal1 24886 34034 24886 34034 0 _0327_
rlabel metal1 24656 32878 24656 32878 0 _0328_
rlabel metal1 25530 32878 25530 32878 0 _0329_
rlabel metal1 18170 31314 18170 31314 0 _0330_
rlabel metal2 17986 33660 17986 33660 0 _0331_
rlabel metal1 29808 39474 29808 39474 0 _0332_
rlabel metal1 28704 39610 28704 39610 0 _0333_
rlabel metal2 28566 43384 28566 43384 0 _0334_
rlabel metal2 29210 40188 29210 40188 0 _0335_
rlabel metal2 32246 40630 32246 40630 0 _0336_
rlabel metal1 29762 36754 29762 36754 0 _0337_
rlabel metal1 30168 40154 30168 40154 0 _0338_
rlabel metal1 29578 40018 29578 40018 0 _0339_
rlabel metal1 20424 33626 20424 33626 0 _0340_
rlabel metal1 18308 31246 18308 31246 0 _0341_
rlabel metal1 18262 31824 18262 31824 0 _0342_
rlabel metal1 18400 40018 18400 40018 0 _0343_
rlabel metal1 19872 44370 19872 44370 0 _0344_
rlabel metal1 18538 43248 18538 43248 0 _0345_
rlabel metal1 18906 43316 18906 43316 0 _0346_
rlabel metal1 26220 42738 26220 42738 0 _0347_
rlabel metal2 20286 43078 20286 43078 0 _0348_
rlabel via1 23529 43282 23529 43282 0 _0349_
rlabel metal2 23782 42976 23782 42976 0 _0350_
rlabel metal1 20470 43350 20470 43350 0 _0351_
rlabel metal1 18998 40562 18998 40562 0 _0352_
rlabel metal2 18538 39984 18538 39984 0 _0353_
rlabel metal1 18576 39338 18576 39338 0 _0354_
rlabel metal2 18078 35530 18078 35530 0 _0355_
rlabel metal2 16698 31042 16698 31042 0 _0356_
rlabel metal1 15732 31450 15732 31450 0 _0357_
rlabel metal1 15088 31314 15088 31314 0 _0358_
rlabel metal2 15410 31994 15410 31994 0 _0359_
rlabel metal1 14858 31280 14858 31280 0 _0360_
rlabel metal2 16974 30158 16974 30158 0 _0361_
rlabel metal1 33810 34646 33810 34646 0 _0362_
rlabel metal1 19596 38386 19596 38386 0 _0363_
rlabel metal2 20010 36176 20010 36176 0 _0364_
rlabel metal1 27048 36074 27048 36074 0 _0365_
rlabel metal1 30958 42058 30958 42058 0 _0366_
rlabel metal2 30774 41786 30774 41786 0 _0367_
rlabel metal1 32568 38998 32568 38998 0 _0368_
rlabel metal1 29900 41514 29900 41514 0 _0369_
rlabel metal2 30682 41990 30682 41990 0 _0370_
rlabel metal1 28290 40086 28290 40086 0 _0371_
rlabel via1 20554 30634 20554 30634 0 _0372_
rlabel metal2 23782 34850 23782 34850 0 _0373_
rlabel metal1 22954 34578 22954 34578 0 _0374_
rlabel metal1 24518 38454 24518 38454 0 _0375_
rlabel metal1 32039 34578 32039 34578 0 _0376_
rlabel metal1 25208 36210 25208 36210 0 _0377_
rlabel metal3 26381 37060 26381 37060 0 _0378_
rlabel metal2 24794 35530 24794 35530 0 _0379_
rlabel metal1 24334 33558 24334 33558 0 _0380_
rlabel metal2 23506 33252 23506 33252 0 _0381_
rlabel metal2 23598 32810 23598 32810 0 _0382_
rlabel metal1 24150 31994 24150 31994 0 _0383_
rlabel metal1 20976 31722 20976 31722 0 _0384_
rlabel metal2 25990 33252 25990 33252 0 _0385_
rlabel metal1 19642 32436 19642 32436 0 _0386_
rlabel metal2 27462 40154 27462 40154 0 _0387_
rlabel metal1 26772 39610 26772 39610 0 _0388_
rlabel metal1 28060 38794 28060 38794 0 _0389_
rlabel metal1 27876 39542 27876 39542 0 _0390_
rlabel metal1 27600 39610 27600 39610 0 _0391_
rlabel metal2 27508 39542 27508 39542 0 _0392_
rlabel metal2 20010 32028 20010 32028 0 _0393_
rlabel metal1 20516 30906 20516 30906 0 _0394_
rlabel metal2 20194 30396 20194 30396 0 _0395_
rlabel metal1 20378 30600 20378 30600 0 _0396_
rlabel metal1 19550 29614 19550 29614 0 _0397_
rlabel metal2 18630 32028 18630 32028 0 _0398_
rlabel metal1 18492 30226 18492 30226 0 _0399_
rlabel metal1 18584 28458 18584 28458 0 _0400_
rlabel metal1 19090 28526 19090 28526 0 _0401_
rlabel metal1 18630 28560 18630 28560 0 _0402_
rlabel metal1 20838 29682 20838 29682 0 _0403_
rlabel metal1 22632 34510 22632 34510 0 _0404_
rlabel metal2 22034 32912 22034 32912 0 _0405_
rlabel metal2 22586 30906 22586 30906 0 _0406_
rlabel metal2 23046 32266 23046 32266 0 _0407_
rlabel metal2 21896 39100 21896 39100 0 _0408_
rlabel metal1 25530 36788 25530 36788 0 _0409_
rlabel metal1 32798 36788 32798 36788 0 _0410_
rlabel metal2 32706 38828 32706 38828 0 _0411_
rlabel metal1 25622 36652 25622 36652 0 _0412_
rlabel metal2 25806 32164 25806 32164 0 _0413_
rlabel metal2 22770 31178 22770 31178 0 _0414_
rlabel metal2 21758 29818 21758 29818 0 _0415_
rlabel metal2 24242 35785 24242 35785 0 _0416_
rlabel metal1 24932 35666 24932 35666 0 _0417_
rlabel metal1 26772 35802 26772 35802 0 _0418_
rlabel metal1 24794 35802 24794 35802 0 _0419_
rlabel metal1 21643 32810 21643 32810 0 _0420_
rlabel metal2 21298 33354 21298 33354 0 _0421_
rlabel metal1 21942 32912 21942 32912 0 _0422_
rlabel metal2 21850 30192 21850 30192 0 _0423_
rlabel metal2 20838 29376 20838 29376 0 _0424_
rlabel metal1 20010 29614 20010 29614 0 _0425_
rlabel metal2 20010 29308 20010 29308 0 _0426_
rlabel metal1 20056 29002 20056 29002 0 _0427_
rlabel metal2 17986 30566 17986 30566 0 _0428_
rlabel metal1 25392 33626 25392 33626 0 _0429_
rlabel metal2 26450 34034 26450 34034 0 _0430_
rlabel metal1 33672 40494 33672 40494 0 _0431_
rlabel viali 31782 40494 31782 40494 0 _0432_
rlabel metal1 32200 41990 32200 41990 0 _0433_
rlabel metal2 31326 39644 31326 39644 0 _0434_
rlabel metal1 31510 39032 31510 39032 0 _0435_
rlabel metal2 30222 38692 30222 38692 0 _0436_
rlabel metal1 31694 38896 31694 38896 0 _0437_
rlabel via3 31165 38692 31165 38692 0 _0438_
rlabel metal1 24886 31348 24886 31348 0 _0439_
rlabel metal1 24656 30226 24656 30226 0 _0440_
rlabel metal2 24886 40052 24886 40052 0 _0441_
rlabel metal1 24610 39814 24610 39814 0 _0442_
rlabel metal1 23414 42602 23414 42602 0 _0443_
rlabel metal3 24357 38692 24357 38692 0 _0444_
rlabel metal1 30498 31824 30498 31824 0 _0445_
rlabel metal1 24288 30634 24288 30634 0 _0446_
rlabel metal1 24840 30226 24840 30226 0 _0447_
rlabel metal1 24288 28526 24288 28526 0 _0448_
rlabel metal1 33304 39406 33304 39406 0 _0449_
rlabel metal2 32706 36006 32706 36006 0 _0450_
rlabel metal2 31970 35530 31970 35530 0 _0451_
rlabel metal2 27278 34748 27278 34748 0 _0452_
rlabel metal2 32154 35564 32154 35564 0 _0453_
rlabel metal1 31510 34918 31510 34918 0 _0454_
rlabel metal1 24702 34102 24702 34102 0 _0455_
rlabel metal2 23782 29614 23782 29614 0 _0456_
rlabel metal2 23598 28764 23598 28764 0 _0457_
rlabel metal2 22494 27982 22494 27982 0 _0458_
rlabel metal1 22264 30566 22264 30566 0 _0459_
rlabel metal1 22356 29818 22356 29818 0 _0460_
rlabel metal2 22310 29682 22310 29682 0 _0461_
rlabel metal2 20930 27676 20930 27676 0 _0462_
rlabel metal1 19826 29580 19826 29580 0 _0463_
rlabel metal1 19136 28118 19136 28118 0 _0464_
rlabel metal1 20286 27982 20286 27982 0 _0465_
rlabel metal1 27324 41582 27324 41582 0 _0466_
rlabel metal1 26910 41786 26910 41786 0 _0467_
rlabel metal3 27991 34340 27991 34340 0 _0468_
rlabel metal1 30544 35666 30544 35666 0 _0469_
rlabel via1 30958 36550 30958 36550 0 _0470_
rlabel metal1 28382 33966 28382 33966 0 _0471_
rlabel metal3 27623 34476 27623 34476 0 _0472_
rlabel metal1 28198 33830 28198 33830 0 _0473_
rlabel metal2 28474 30396 28474 30396 0 _0474_
rlabel metal1 29394 29614 29394 29614 0 _0475_
rlabel metal2 30130 36890 30130 36890 0 _0476_
rlabel metal2 29670 33932 29670 33932 0 _0477_
rlabel metal2 30130 30430 30130 30430 0 _0478_
rlabel metal1 30820 29206 30820 29206 0 _0479_
rlabel metal1 32292 37230 32292 37230 0 _0480_
rlabel metal1 27922 37332 27922 37332 0 _0481_
rlabel metal2 31234 35292 31234 35292 0 _0482_
rlabel metal1 30774 30770 30774 30770 0 _0483_
rlabel metal2 30958 29886 30958 29886 0 _0484_
rlabel metal2 30774 28050 30774 28050 0 _0485_
rlabel metal1 27738 28662 27738 28662 0 _0486_
rlabel metal1 25300 29138 25300 29138 0 _0487_
rlabel metal2 25162 27948 25162 27948 0 _0488_
rlabel metal1 21206 26996 21206 26996 0 _0489_
rlabel metal2 22310 28220 22310 28220 0 _0490_
rlabel metal1 24426 27982 24426 27982 0 _0491_
rlabel metal2 21390 27404 21390 27404 0 _0492_
rlabel metal1 27140 35734 27140 35734 0 _0493_
rlabel metal2 27186 34476 27186 34476 0 _0494_
rlabel metal1 27646 33898 27646 33898 0 _0495_
rlabel metal1 29578 33626 29578 33626 0 _0496_
rlabel metal1 28842 34034 28842 34034 0 _0497_
rlabel metal1 30130 34102 30130 34102 0 _0498_
rlabel metal2 25622 41412 25622 41412 0 _0499_
rlabel metal2 25714 41548 25714 41548 0 _0500_
rlabel metal2 25162 41276 25162 41276 0 _0501_
rlabel metal1 24518 40698 24518 40698 0 _0502_
rlabel metal1 24978 41072 24978 41072 0 _0503_
rlabel metal1 25438 31790 25438 31790 0 _0504_
rlabel metal2 25990 31076 25990 31076 0 _0505_
rlabel metal2 26082 31484 26082 31484 0 _0506_
rlabel metal1 29624 31382 29624 31382 0 _0507_
rlabel metal2 33994 30770 33994 30770 0 _0508_
rlabel metal2 31510 31110 31510 31110 0 _0509_
rlabel metal1 33350 31416 33350 31416 0 _0510_
rlabel metal1 33994 33558 33994 33558 0 _0511_
rlabel metal1 32614 33456 32614 33456 0 _0512_
rlabel metal2 31970 33796 31970 33796 0 _0513_
rlabel metal2 32522 33286 32522 33286 0 _0514_
rlabel metal1 32522 31824 32522 31824 0 _0515_
rlabel metal2 32982 30906 32982 30906 0 _0516_
rlabel metal1 32660 30702 32660 30702 0 _0517_
rlabel metal1 32706 30022 32706 30022 0 _0518_
rlabel metal1 30222 29240 30222 29240 0 _0519_
rlabel metal2 32798 29376 32798 29376 0 _0520_
rlabel metal2 33626 28254 33626 28254 0 _0521_
rlabel metal2 25438 28220 25438 28220 0 _0522_
rlabel metal1 25622 28084 25622 28084 0 _0523_
rlabel metal1 27830 27846 27830 27846 0 _0524_
rlabel metal1 20286 28594 20286 28594 0 _0525_
rlabel metal2 30406 28254 30406 28254 0 _0526_
rlabel metal1 19458 29002 19458 29002 0 _0527_
rlabel metal1 32706 29172 32706 29172 0 _0528_
rlabel metal2 33166 28662 33166 28662 0 _0529_
rlabel metal1 33902 30736 33902 30736 0 _0530_
rlabel metal1 32706 40052 32706 40052 0 _0531_
rlabel metal1 32384 39610 32384 39610 0 _0532_
rlabel metal1 32614 39814 32614 39814 0 _0533_
rlabel metal1 26634 33456 26634 33456 0 _0534_
rlabel via1 26357 32878 26357 32878 0 _0535_
rlabel metal1 26592 32946 26592 32946 0 _0536_
rlabel metal1 31280 32198 31280 32198 0 _0537_
rlabel metal2 30406 32164 30406 32164 0 _0538_
rlabel metal2 31142 34748 31142 34748 0 _0539_
rlabel metal1 30222 32368 30222 32368 0 _0540_
rlabel metal1 31096 32402 31096 32402 0 _0541_
rlabel metal1 33396 31790 33396 31790 0 _0542_
rlabel metal1 34500 41038 34500 41038 0 _0543_
rlabel metal2 33258 36992 33258 36992 0 _0544_
rlabel metal2 32706 34442 32706 34442 0 _0545_
rlabel metal1 33718 32436 33718 32436 0 _0546_
rlabel metal2 33626 32572 33626 32572 0 _0547_
rlabel metal1 35190 32334 35190 32334 0 _0548_
rlabel metal2 34086 30940 34086 30940 0 _0549_
rlabel metal1 36754 31416 36754 31416 0 _0550_
rlabel metal1 34562 30294 34562 30294 0 _0551_
rlabel metal1 35926 30158 35926 30158 0 _0552_
rlabel metal2 37214 30906 37214 30906 0 _0553_
rlabel metal1 35006 31246 35006 31246 0 _0554_
rlabel metal2 36110 29682 36110 29682 0 _0555_
rlabel metal1 37030 30294 37030 30294 0 _0556_
rlabel metal1 34868 30906 34868 30906 0 _0557_
rlabel metal2 36018 30906 36018 30906 0 _0558_
rlabel metal1 33534 32538 33534 32538 0 _0559_
rlabel metal1 28244 32878 28244 32878 0 _0560_
rlabel metal2 27922 35326 27922 35326 0 _0561_
rlabel metal1 28428 32946 28428 32946 0 _0562_
rlabel metal1 29394 32878 29394 32878 0 _0563_
rlabel metal1 34776 33966 34776 33966 0 _0564_
rlabel metal1 30728 33898 30728 33898 0 _0565_
rlabel metal1 34362 34034 34362 34034 0 _0566_
rlabel metal1 35466 34000 35466 34000 0 _0567_
rlabel metal2 33442 34510 33442 34510 0 _0568_
rlabel metal1 33350 33932 33350 33932 0 _0569_
rlabel metal2 35558 34374 35558 34374 0 _0570_
rlabel metal2 35650 33932 35650 33932 0 _0571_
rlabel metal2 35834 33660 35834 33660 0 _0572_
rlabel metal1 35604 32402 35604 32402 0 _0573_
rlabel metal1 38962 32334 38962 32334 0 _0574_
rlabel metal2 36018 32708 36018 32708 0 _0575_
rlabel metal2 35650 32266 35650 32266 0 _0576_
rlabel viali 38686 32330 38686 32330 0 _0577_
rlabel metal1 35604 30294 35604 30294 0 _0578_
rlabel metal1 36294 31824 36294 31824 0 _0579_
rlabel metal1 35696 56678 35696 56678 0 _0580_
rlabel metal1 38594 33626 38594 33626 0 _0581_
rlabel metal1 36662 32844 36662 32844 0 _0582_
rlabel metal1 37260 34510 37260 34510 0 _0583_
rlabel metal2 38962 34204 38962 34204 0 _0584_
rlabel metal2 40250 33490 40250 33490 0 _0585_
rlabel metal1 39054 32776 39054 32776 0 _0586_
rlabel metal1 40250 33082 40250 33082 0 _0587_
rlabel metal1 39652 32538 39652 32538 0 _0588_
rlabel metal1 37490 31858 37490 31858 0 _0589_
rlabel metal2 36846 33082 36846 33082 0 _0590_
rlabel metal1 37674 32912 37674 32912 0 _0591_
rlabel metal2 37950 32572 37950 32572 0 _0592_
rlabel metal1 38594 32436 38594 32436 0 _0593_
rlabel metal1 38134 32198 38134 32198 0 _0594_
rlabel metal2 37674 32198 37674 32198 0 _0595_
rlabel metal2 16422 37434 16422 37434 0 _0596_
rlabel metal2 41170 21063 41170 21063 0 _0597_
rlabel metal2 41078 26146 41078 26146 0 _0598_
rlabel metal2 42918 20876 42918 20876 0 _0599_
rlabel metal1 43976 18190 43976 18190 0 _0600_
rlabel metal2 37858 16354 37858 16354 0 _0601_
rlabel metal1 42826 24854 42826 24854 0 _0602_
rlabel metal1 36386 25908 36386 25908 0 _0603_
rlabel metal1 36570 19686 36570 19686 0 _0604_
rlabel metal1 44022 19822 44022 19822 0 _0605_
rlabel metal1 40526 20434 40526 20434 0 _0606_
rlabel metal1 44712 19482 44712 19482 0 _0607_
rlabel metal1 36616 18666 36616 18666 0 _0608_
rlabel metal1 37628 16082 37628 16082 0 _0609_
rlabel metal1 41124 18734 41124 18734 0 _0610_
rlabel metal1 40204 15946 40204 15946 0 _0611_
rlabel metal2 41354 17068 41354 17068 0 _0612_
rlabel via1 43554 17578 43554 17578 0 _0613_
rlabel metal1 40204 16558 40204 16558 0 _0614_
rlabel metal1 40342 16524 40342 16524 0 _0615_
rlabel metal2 35742 21607 35742 21607 0 _0616_
rlabel metal2 39514 16354 39514 16354 0 _0617_
rlabel metal1 40894 14042 40894 14042 0 _0618_
rlabel metal1 39652 17102 39652 17102 0 _0619_
rlabel metal1 38778 26010 38778 26010 0 _0620_
rlabel metal1 40020 16966 40020 16966 0 _0621_
rlabel metal1 39698 25466 39698 25466 0 _0622_
rlabel metal2 40434 16524 40434 16524 0 _0623_
rlabel metal1 40020 16082 40020 16082 0 _0624_
rlabel metal1 41078 12852 41078 12852 0 _0625_
rlabel metal2 40526 20332 40526 20332 0 _0626_
rlabel metal2 32614 17612 32614 17612 0 _0627_
rlabel metal1 39698 14994 39698 14994 0 _0628_
rlabel metal1 39284 11526 39284 11526 0 _0629_
rlabel metal2 30038 9146 30038 9146 0 _0630_
rlabel metal1 39652 10710 39652 10710 0 _0631_
rlabel metal1 35926 18326 35926 18326 0 _0632_
rlabel metal1 41676 24922 41676 24922 0 _0633_
rlabel metal1 36616 19346 36616 19346 0 _0634_
rlabel metal1 41216 13906 41216 13906 0 _0635_
rlabel metal1 36570 13430 36570 13430 0 _0636_
rlabel metal2 36478 13770 36478 13770 0 _0637_
rlabel metal1 40894 21352 40894 21352 0 _0638_
rlabel metal1 42458 14926 42458 14926 0 _0639_
rlabel metal1 35512 13838 35512 13838 0 _0640_
rlabel metal1 37950 15538 37950 15538 0 _0641_
rlabel metal1 43792 20434 43792 20434 0 _0642_
rlabel metal2 43378 21216 43378 21216 0 _0643_
rlabel via2 41262 16541 41262 16541 0 _0644_
rlabel metal2 45126 15708 45126 15708 0 _0645_
rlabel metal1 44528 16014 44528 16014 0 _0646_
rlabel metal2 43654 14824 43654 14824 0 _0647_
rlabel metal1 36340 13702 36340 13702 0 _0648_
rlabel metal1 33948 20910 33948 20910 0 _0649_
rlabel metal2 33994 15028 33994 15028 0 _0650_
rlabel metal1 36938 17578 36938 17578 0 _0651_
rlabel metal1 36432 18258 36432 18258 0 _0652_
rlabel metal2 35926 17782 35926 17782 0 _0653_
rlabel metal1 34914 18224 34914 18224 0 _0654_
rlabel metal1 34730 18190 34730 18190 0 _0655_
rlabel metal1 34868 18054 34868 18054 0 _0656_
rlabel metal1 36202 17782 36202 17782 0 _0657_
rlabel metal1 35880 16558 35880 16558 0 _0658_
rlabel metal2 34500 12818 34500 12818 0 _0659_
rlabel metal2 38594 10540 38594 10540 0 _0660_
rlabel metal2 39146 9996 39146 9996 0 _0661_
rlabel metal1 30820 10234 30820 10234 0 _0662_
rlabel metal1 41354 16490 41354 16490 0 _0663_
rlabel metal1 37720 21658 37720 21658 0 _0664_
rlabel via1 34638 19316 34638 19316 0 _0665_
rlabel metal1 38456 16558 38456 16558 0 _0666_
rlabel metal1 38318 19822 38318 19822 0 _0667_
rlabel metal1 39054 19346 39054 19346 0 _0668_
rlabel metal1 36754 21522 36754 21522 0 _0669_
rlabel metal1 39100 16762 39100 16762 0 _0670_
rlabel metal1 38594 16524 38594 16524 0 _0671_
rlabel metal1 35144 12818 35144 12818 0 _0672_
rlabel metal1 33810 10234 33810 10234 0 _0673_
rlabel metal1 42274 13328 42274 13328 0 _0674_
rlabel metal1 33672 22406 33672 22406 0 _0675_
rlabel metal1 42136 18938 42136 18938 0 _0676_
rlabel metal2 42734 16235 42734 16235 0 _0677_
rlabel via2 40526 20757 40526 20757 0 _0678_
rlabel metal2 36018 24208 36018 24208 0 _0679_
rlabel metal1 42044 14994 42044 14994 0 _0680_
rlabel metal1 43194 15028 43194 15028 0 _0681_
rlabel metal1 43976 14790 43976 14790 0 _0682_
rlabel metal1 45126 17510 45126 17510 0 _0683_
rlabel metal1 44252 16422 44252 16422 0 _0684_
rlabel metal1 43470 14892 43470 14892 0 _0685_
rlabel metal2 43378 14688 43378 14688 0 _0686_
rlabel metal2 33902 10302 33902 10302 0 _0687_
rlabel metal2 33718 9724 33718 9724 0 _0688_
rlabel metal2 44298 14076 44298 14076 0 _0689_
rlabel metal1 38410 17612 38410 17612 0 _0690_
rlabel metal2 42182 13498 42182 13498 0 _0691_
rlabel metal1 32752 19754 32752 19754 0 _0692_
rlabel metal1 35650 16966 35650 16966 0 _0693_
rlabel metal1 38962 22610 38962 22610 0 _0694_
rlabel metal2 42458 14212 42458 14212 0 _0695_
rlabel metal2 40342 20604 40342 20604 0 _0696_
rlabel metal1 43700 13430 43700 13430 0 _0697_
rlabel metal1 42780 13294 42780 13294 0 _0698_
rlabel metal1 39054 11730 39054 11730 0 _0699_
rlabel metal1 37260 11186 37260 11186 0 _0700_
rlabel metal2 43930 15980 43930 15980 0 _0701_
rlabel metal1 43286 15436 43286 15436 0 _0702_
rlabel metal2 41170 22304 41170 22304 0 _0703_
rlabel metal2 41814 22814 41814 22814 0 _0704_
rlabel metal2 42550 15521 42550 15521 0 _0705_
rlabel metal2 38226 12886 38226 12886 0 _0706_
rlabel metal2 37490 9758 37490 9758 0 _0707_
rlabel metal1 34500 9554 34500 9554 0 _0708_
rlabel metal1 31602 8942 31602 8942 0 _0709_
rlabel metal2 32982 9282 32982 9282 0 _0710_
rlabel metal1 36064 22066 36064 22066 0 _0711_
rlabel via2 39330 22661 39330 22661 0 _0712_
rlabel metal2 35742 22236 35742 22236 0 _0713_
rlabel metal2 38870 14348 38870 14348 0 _0714_
rlabel metal1 34040 23290 34040 23290 0 _0715_
rlabel metal2 33810 20332 33810 20332 0 _0716_
rlabel metal2 34454 23052 34454 23052 0 _0717_
rlabel via1 39514 22474 39514 22474 0 _0718_
rlabel metal1 34546 22576 34546 22576 0 _0719_
rlabel metal1 31464 11866 31464 11866 0 _0720_
rlabel metal1 37766 19686 37766 19686 0 _0721_
rlabel metal1 36386 20400 36386 20400 0 _0722_
rlabel metal1 37812 13430 37812 13430 0 _0723_
rlabel metal2 37858 12988 37858 12988 0 _0724_
rlabel metal1 41262 12750 41262 12750 0 _0725_
rlabel metal1 39422 12852 39422 12852 0 _0726_
rlabel metal2 39698 12988 39698 12988 0 _0727_
rlabel metal1 37674 12784 37674 12784 0 _0728_
rlabel metal1 37168 12614 37168 12614 0 _0729_
rlabel metal1 31602 11662 31602 11662 0 _0730_
rlabel metal1 31464 12614 31464 12614 0 _0731_
rlabel metal1 28520 12750 28520 12750 0 _0732_
rlabel metal1 28474 12206 28474 12206 0 _0733_
rlabel metal1 31326 11696 31326 11696 0 _0734_
rlabel metal1 31188 11866 31188 11866 0 _0735_
rlabel metal1 41538 16116 41538 16116 0 _0736_
rlabel metal1 42182 16524 42182 16524 0 _0737_
rlabel metal2 41538 15640 41538 15640 0 _0738_
rlabel metal2 33810 19873 33810 19873 0 _0739_
rlabel metal2 41078 14586 41078 14586 0 _0740_
rlabel metal2 41538 13260 41538 13260 0 _0741_
rlabel metal2 40894 13634 40894 13634 0 _0742_
rlabel metal2 40710 14263 40710 14263 0 _0743_
rlabel metal2 35006 14212 35006 14212 0 _0744_
rlabel metal1 36524 16150 36524 16150 0 _0745_
rlabel metal2 40894 21063 40894 21063 0 _0746_
rlabel metal2 35282 14110 35282 14110 0 _0747_
rlabel metal1 37122 12682 37122 12682 0 _0748_
rlabel metal1 35420 12954 35420 12954 0 _0749_
rlabel metal1 32706 12852 32706 12852 0 _0750_
rlabel metal1 30912 11730 30912 11730 0 _0751_
rlabel metal1 30452 11866 30452 11866 0 _0752_
rlabel metal2 31510 10472 31510 10472 0 _0753_
rlabel metal1 33258 8602 33258 8602 0 _0754_
rlabel metal2 33902 8636 33902 8636 0 _0755_
rlabel metal1 32578 14960 32578 14960 0 _0756_
rlabel metal1 34684 11798 34684 11798 0 _0757_
rlabel metal2 33258 14790 33258 14790 0 _0758_
rlabel metal2 34454 11934 34454 11934 0 _0759_
rlabel metal1 34868 9554 34868 9554 0 _0760_
rlabel metal2 36110 10268 36110 10268 0 _0761_
rlabel metal2 35742 9724 35742 9724 0 _0762_
rlabel metal1 35374 8602 35374 8602 0 _0763_
rlabel metal1 35742 11560 35742 11560 0 _0764_
rlabel metal1 35804 11798 35804 11798 0 _0765_
rlabel metal2 35926 9996 35926 9996 0 _0766_
rlabel metal1 34868 8466 34868 8466 0 _0767_
rlabel metal1 33626 8432 33626 8432 0 _0768_
rlabel metal1 33074 7820 33074 7820 0 _0769_
rlabel metal2 33258 8058 33258 8058 0 _0770_
rlabel metal2 33718 7174 33718 7174 0 _0771_
rlabel metal2 38318 10234 38318 10234 0 _0772_
rlabel metal2 37674 9418 37674 9418 0 _0773_
rlabel metal2 36110 8636 36110 8636 0 _0774_
rlabel metal1 37812 8330 37812 8330 0 _0775_
rlabel metal1 35466 7854 35466 7854 0 _0776_
rlabel via1 31142 9146 31142 9146 0 _0777_
rlabel metal2 33534 10880 33534 10880 0 _0778_
rlabel metal1 42090 23120 42090 23120 0 _0779_
rlabel metal1 41124 23154 41124 23154 0 _0780_
rlabel metal1 41538 22746 41538 22746 0 _0781_
rlabel metal1 41124 20434 41124 20434 0 _0782_
rlabel metal1 40526 21522 40526 21522 0 _0783_
rlabel metal2 40342 24582 40342 24582 0 _0784_
rlabel metal2 41078 25568 41078 25568 0 _0785_
rlabel metal1 40848 24242 40848 24242 0 _0786_
rlabel metal2 40710 24480 40710 24480 0 _0787_
rlabel metal1 40802 23086 40802 23086 0 _0788_
rlabel metal1 34408 14042 34408 14042 0 _0789_
rlabel metal2 32522 10710 32522 10710 0 _0790_
rlabel metal1 32836 10778 32836 10778 0 _0791_
rlabel metal1 28658 11152 28658 11152 0 _0792_
rlabel metal1 36800 11322 36800 11322 0 _0793_
rlabel metal1 42320 19890 42320 19890 0 _0794_
rlabel metal2 41722 20094 41722 20094 0 _0795_
rlabel metal1 41124 18258 41124 18258 0 _0796_
rlabel metal1 40342 19856 40342 19856 0 _0797_
rlabel metal1 39422 18938 39422 18938 0 _0798_
rlabel metal1 40434 18054 40434 18054 0 _0799_
rlabel metal1 44482 17680 44482 17680 0 _0800_
rlabel metal2 41538 18020 41538 18020 0 _0801_
rlabel metal1 40848 18394 40848 18394 0 _0802_
rlabel metal1 28566 11220 28566 11220 0 _0803_
rlabel metal1 29394 11118 29394 11118 0 _0804_
rlabel metal1 28980 12410 28980 12410 0 _0805_
rlabel metal2 32614 12580 32614 12580 0 _0806_
rlabel metal1 29854 12376 29854 12376 0 _0807_
rlabel metal1 30268 12750 30268 12750 0 _0808_
rlabel metal1 29900 10098 29900 10098 0 _0809_
rlabel metal2 31050 9826 31050 9826 0 _0810_
rlabel metal1 30728 8466 30728 8466 0 _0811_
rlabel metal1 31280 8602 31280 8602 0 _0812_
rlabel metal2 31418 7548 31418 7548 0 _0813_
rlabel metal1 31280 7310 31280 7310 0 _0814_
rlabel metal1 28888 15470 28888 15470 0 _0815_
rlabel metal1 29624 11322 29624 11322 0 _0816_
rlabel metal1 36478 18326 36478 18326 0 _0817_
rlabel metal1 33258 14994 33258 14994 0 _0818_
rlabel metal1 38226 21114 38226 21114 0 _0819_
rlabel metal1 39376 20570 39376 20570 0 _0820_
rlabel metal1 38134 22202 38134 22202 0 _0821_
rlabel metal1 39560 21862 39560 21862 0 _0822_
rlabel metal1 38640 22542 38640 22542 0 _0823_
rlabel metal1 38042 15470 38042 15470 0 _0824_
rlabel metal1 33810 15028 33810 15028 0 _0825_
rlabel metal2 32798 13906 32798 13906 0 _0826_
rlabel metal1 32890 14042 32890 14042 0 _0827_
rlabel metal1 43470 21522 43470 21522 0 _0828_
rlabel metal2 27646 15810 27646 15810 0 _0829_
rlabel metal1 34638 11594 34638 11594 0 _0830_
rlabel metal1 27370 17850 27370 17850 0 _0831_
rlabel metal1 34868 15674 34868 15674 0 _0832_
rlabel metal1 34592 20230 34592 20230 0 _0833_
rlabel metal2 34638 17476 34638 17476 0 _0834_
rlabel metal2 39330 14144 39330 14144 0 _0835_
rlabel metal1 35236 18598 35236 18598 0 _0836_
rlabel metal1 39238 19312 39238 19312 0 _0837_
rlabel metal2 38870 18972 38870 18972 0 _0838_
rlabel metal1 33902 22032 33902 22032 0 _0839_
rlabel metal1 33327 18870 33327 18870 0 _0840_
rlabel metal2 27278 17544 27278 17544 0 _0841_
rlabel metal2 27462 16252 27462 16252 0 _0842_
rlabel metal1 30866 14246 30866 14246 0 _0843_
rlabel metal1 31372 16082 31372 16082 0 _0844_
rlabel metal1 35558 22202 35558 22202 0 _0845_
rlabel metal1 36156 18938 36156 18938 0 _0846_
rlabel metal1 32798 18292 32798 18292 0 _0847_
rlabel metal2 31418 17850 31418 17850 0 _0848_
rlabel metal1 37651 17646 37651 17646 0 _0849_
rlabel metal1 37858 23596 37858 23596 0 _0850_
rlabel metal1 37168 17646 37168 17646 0 _0851_
rlabel metal1 31970 17612 31970 17612 0 _0852_
rlabel metal2 31142 16796 31142 16796 0 _0853_
rlabel metal1 30498 16014 30498 16014 0 _0854_
rlabel metal1 29946 15878 29946 15878 0 _0855_
rlabel metal1 27554 15980 27554 15980 0 _0856_
rlabel metal1 28842 16082 28842 16082 0 _0857_
rlabel via1 28382 16490 28382 16490 0 _0858_
rlabel metal2 28566 16116 28566 16116 0 _0859_
rlabel metal1 29118 16762 29118 16762 0 _0860_
rlabel metal1 32338 20876 32338 20876 0 _0861_
rlabel metal1 30452 8398 30452 8398 0 _0862_
rlabel metal2 25990 16898 25990 16898 0 _0863_
rlabel metal1 25760 16082 25760 16082 0 _0864_
rlabel metal1 33258 15538 33258 15538 0 _0865_
rlabel metal1 33396 18734 33396 18734 0 _0866_
rlabel metal1 41101 18598 41101 18598 0 _0867_
rlabel metal1 34914 18666 34914 18666 0 _0868_
rlabel metal2 32706 16796 32706 16796 0 _0869_
rlabel metal2 32614 15300 32614 15300 0 _0870_
rlabel metal1 34270 18938 34270 18938 0 _0871_
rlabel metal1 32062 15538 32062 15538 0 _0872_
rlabel metal2 31970 15674 31970 15674 0 _0873_
rlabel metal1 25530 19346 25530 19346 0 _0874_
rlabel metal1 27968 19754 27968 19754 0 _0875_
rlabel metal1 26956 19482 26956 19482 0 _0876_
rlabel metal1 38962 13498 38962 13498 0 _0877_
rlabel metal2 40066 15164 40066 15164 0 _0878_
rlabel metal1 39284 14994 39284 14994 0 _0879_
rlabel via2 38594 14875 38594 14875 0 _0880_
rlabel metal1 25990 19958 25990 19958 0 _0881_
rlabel metal1 32476 21386 32476 21386 0 _0882_
rlabel metal2 25806 18938 25806 18938 0 _0883_
rlabel metal1 30130 14586 30130 14586 0 _0884_
rlabel metal1 25622 18156 25622 18156 0 _0885_
rlabel metal1 25622 17646 25622 17646 0 _0886_
rlabel metal1 26588 17646 26588 17646 0 _0887_
rlabel metal1 25990 17782 25990 17782 0 _0888_
rlabel metal2 26082 17340 26082 17340 0 _0889_
rlabel metal2 25070 16558 25070 16558 0 _0890_
rlabel metal2 26082 20434 26082 20434 0 _0891_
rlabel metal1 37122 24140 37122 24140 0 _0892_
rlabel metal1 25944 20910 25944 20910 0 _0893_
rlabel metal1 35880 20910 35880 20910 0 _0894_
rlabel metal1 40304 20502 40304 20502 0 _0895_
rlabel metal1 35696 20570 35696 20570 0 _0896_
rlabel metal1 37398 20910 37398 20910 0 _0897_
rlabel metal2 35926 20876 35926 20876 0 _0898_
rlabel metal1 35834 20502 35834 20502 0 _0899_
rlabel metal1 35006 20298 35006 20298 0 _0900_
rlabel metal1 32062 23698 32062 23698 0 _0901_
rlabel metal1 32062 23086 32062 23086 0 _0902_
rlabel metal2 37306 24378 37306 24378 0 _0903_
rlabel metal1 28290 23562 28290 23562 0 _0904_
rlabel metal2 27830 23562 27830 23562 0 _0905_
rlabel metal2 29118 20672 29118 20672 0 _0906_
rlabel metal1 35236 23086 35236 23086 0 _0907_
rlabel metal1 33212 22134 33212 22134 0 _0908_
rlabel metal1 33810 21862 33810 21862 0 _0909_
rlabel metal1 33258 20026 33258 20026 0 _0910_
rlabel metal1 31004 22066 31004 22066 0 _0911_
rlabel metal2 27922 23460 27922 23460 0 _0912_
rlabel metal1 27048 21998 27048 21998 0 _0913_
rlabel metal1 37582 13260 37582 13260 0 _0914_
rlabel metal1 39238 20978 39238 20978 0 _0915_
rlabel metal1 39560 22406 39560 22406 0 _0916_
rlabel metal1 38134 19380 38134 19380 0 _0917_
rlabel metal1 40618 19380 40618 19380 0 _0918_
rlabel metal2 40526 19652 40526 19652 0 _0919_
rlabel metal2 40618 20026 40618 20026 0 _0920_
rlabel metal2 40066 20332 40066 20332 0 _0921_
rlabel metal1 30222 21012 30222 21012 0 _0922_
rlabel metal1 29348 20366 29348 20366 0 _0923_
rlabel metal2 27002 21318 27002 21318 0 _0924_
rlabel metal1 36984 21930 36984 21930 0 _0925_
rlabel metal2 25714 21794 25714 21794 0 _0926_
rlabel metal2 25622 21828 25622 21828 0 _0927_
rlabel metal2 25806 21556 25806 21556 0 _0928_
rlabel metal1 25622 23698 25622 23698 0 _0929_
rlabel metal1 25346 23596 25346 23596 0 _0930_
rlabel metal1 25116 16762 25116 16762 0 _0931_
rlabel metal2 26450 23664 26450 23664 0 _0932_
rlabel metal1 27002 23630 27002 23630 0 _0933_
rlabel metal1 27048 23562 27048 23562 0 _0934_
rlabel metal1 31832 21998 31832 21998 0 _0935_
rlabel metal2 32798 22848 32798 22848 0 _0936_
rlabel metal1 34454 21590 34454 21590 0 _0937_
rlabel metal1 34316 21658 34316 21658 0 _0938_
rlabel metal2 32430 22950 32430 22950 0 _0939_
rlabel metal1 30314 23018 30314 23018 0 _0940_
rlabel metal2 29118 24004 29118 24004 0 _0941_
rlabel metal1 36432 22610 36432 22610 0 _0942_
rlabel via1 35926 22627 35926 22627 0 _0943_
rlabel metal1 33718 22610 33718 22610 0 _0944_
rlabel metal2 29026 23460 29026 23460 0 _0945_
rlabel metal2 31234 21318 31234 21318 0 _0946_
rlabel metal1 29854 24174 29854 24174 0 _0947_
rlabel metal1 35320 17238 35320 17238 0 _0948_
rlabel metal2 33994 16762 33994 16762 0 _0949_
rlabel metal2 33810 17136 33810 17136 0 _0950_
rlabel metal2 34086 17408 34086 17408 0 _0951_
rlabel metal2 33442 19040 33442 19040 0 _0952_
rlabel metal1 32292 20026 32292 20026 0 _0953_
rlabel metal1 31602 20468 31602 20468 0 _0954_
rlabel metal1 30774 20434 30774 20434 0 _0955_
rlabel via1 30311 19822 30311 19822 0 _0956_
rlabel metal1 45310 24072 45310 24072 0 _0957_
rlabel metal1 30636 23562 30636 23562 0 _0958_
rlabel metal1 27692 23698 27692 23698 0 _0959_
rlabel metal2 25438 23426 25438 23426 0 _0960_
rlabel metal1 25208 23086 25208 23086 0 _0961_
rlabel metal1 24748 23766 24748 23766 0 _0962_
rlabel metal2 24978 24310 24978 24310 0 _0963_
rlabel metal1 36202 19788 36202 19788 0 _0964_
rlabel metal1 30360 19958 30360 19958 0 _0965_
rlabel metal2 27278 20230 27278 20230 0 _0966_
rlabel metal1 44712 17170 44712 17170 0 _0967_
rlabel metal2 27554 20536 27554 20536 0 _0968_
rlabel metal2 25714 20604 25714 20604 0 _0969_
rlabel metal1 34178 18768 34178 18768 0 _0970_
rlabel metal2 34362 18938 34362 18938 0 _0971_
rlabel metal1 32246 18768 32246 18768 0 _0972_
rlabel metal2 31142 18462 31142 18462 0 _0973_
rlabel metal1 31234 18700 31234 18700 0 _0974_
rlabel metal2 25622 19516 25622 19516 0 _0975_
rlabel metal1 23782 20366 23782 20366 0 _0976_
rlabel metal1 32154 17306 32154 17306 0 _0977_
rlabel metal1 44666 21556 44666 21556 0 _0978_
rlabel metal2 42918 17476 42918 17476 0 _0979_
rlabel metal1 42688 16422 42688 16422 0 _0980_
rlabel metal2 36938 15742 36938 15742 0 _0981_
rlabel metal2 40526 17476 40526 17476 0 _0982_
rlabel metal1 30452 17714 30452 17714 0 _0983_
rlabel metal1 30176 17782 30176 17782 0 _0984_
rlabel metal1 23046 19754 23046 19754 0 _0985_
rlabel metal1 23644 20502 23644 20502 0 _0986_
rlabel metal1 30728 23154 30728 23154 0 _0987_
rlabel metal1 23506 23256 23506 23256 0 _0988_
rlabel metal1 35604 21522 35604 21522 0 _0989_
rlabel metal2 16146 1520 16146 1520 0 addI[0]
rlabel metal3 1188 51748 1188 51748 0 addI[1]
rlabel via2 58282 22491 58282 22491 0 addI[2]
rlabel metal2 27094 1520 27094 1520 0 addI[3]
rlabel metal2 58282 57103 58282 57103 0 addI[4]
rlabel metal1 57822 57562 57822 57562 0 addI[5]
rlabel metal1 19458 57562 19458 57562 0 addQ[0]
rlabel metal1 24610 57562 24610 57562 0 addQ[1]
rlabel metal2 38042 1520 38042 1520 0 addQ[2]
rlabel metal3 1188 28628 1188 28628 0 addQ[3]
rlabel metal2 1702 57715 1702 57715 0 addQ[4]
rlabel metal1 58098 29002 58098 29002 0 addQ[5]
rlabel metal2 27462 27166 27462 27166 0 gen_sym.Reg_2M.data_in
rlabel metal2 29486 26350 29486 26350 0 gen_sym.Reg_2M.data_out
rlabel metal1 26910 26010 26910 26010 0 gen_sym.Reg_2M.enable
rlabel metal1 29670 26486 29670 26486 0 gen_sym.Reg_Sym.data_out\[0\]
rlabel metal2 30958 25534 30958 25534 0 gen_sym.Reg_Sym.data_out\[1\]
rlabel metal2 31510 27166 31510 27166 0 mapper.bit_Q\[1\]
rlabel via3 30613 56644 30613 56644 0 net1
rlabel metal1 57684 40358 57684 40358 0 net10
rlabel metal1 24265 7174 24265 7174 0 net11
rlabel metal1 32384 7174 32384 7174 0 net12
rlabel metal1 46276 57426 46276 57426 0 net13
rlabel metal1 2484 23494 2484 23494 0 net14
rlabel metal1 57454 45798 57454 45798 0 net15
rlabel metal1 2208 34918 2208 34918 0 net16
rlabel metal1 12282 2414 12282 2414 0 net17
rlabel metal1 1932 40494 1932 40494 0 net18
rlabel metal1 2162 17170 2162 17170 0 net19
rlabel metal2 2898 42398 2898 42398 0 net2
rlabel metal1 35420 57018 35420 57018 0 net20
rlabel metal1 52624 57426 52624 57426 0 net21
rlabel via2 57454 17085 57454 17085 0 net22
rlabel metal1 57362 51782 57362 51782 0 net23
rlabel metal1 14030 57426 14030 57426 0 net24
rlabel metal1 1886 2380 1886 2380 0 net25
rlabel metal1 2162 11730 2162 11730 0 net26
rlabel metal2 18906 30940 18906 30940 0 net27
rlabel metal1 9660 57426 9660 57426 0 net28
rlabel metal1 2162 5678 2162 5678 0 net29
rlabel via2 36846 26741 36846 26741 0 net3
rlabel metal2 34454 2655 34454 2655 0 net30
rlabel metal1 41124 57426 41124 57426 0 net31
rlabel via2 17710 2499 17710 2499 0 net32
rlabel metal1 2254 51782 2254 51782 0 net33
rlabel metal1 57776 22610 57776 22610 0 net34
rlabel via2 37490 20859 37490 20859 0 net35
rlabel metal1 57868 56814 57868 56814 0 net36
rlabel metal1 57316 57222 57316 57222 0 net37
rlabel metal1 19734 57392 19734 57392 0 net38
rlabel metal1 25116 57426 25116 57426 0 net39
rlabel metal2 58190 18938 58190 18938 0 net4
rlabel metal1 37352 2618 37352 2618 0 net40
rlabel metal1 2162 29138 2162 29138 0 net41
rlabel metal1 1932 56678 1932 56678 0 net42
rlabel metal1 58098 29104 58098 29104 0 net43
rlabel metal1 33718 43214 33718 43214 0 net44
rlabel metal1 44252 21998 44252 21998 0 net45
rlabel metal1 23552 26554 23552 26554 0 net46
rlabel metal1 36255 29206 36255 29206 0 net47
rlabel metal1 36156 36006 36156 36006 0 net48
rlabel metal1 24978 12274 24978 12274 0 net49
rlabel metal1 6325 2482 6325 2482 0 net5
rlabel metal2 33442 24718 33442 24718 0 net50
rlabel metal2 35742 39644 35742 39644 0 net51
rlabel metal1 57822 5678 57822 5678 0 net6
rlabel metal1 2116 46546 2116 46546 0 net7
rlabel metal1 57776 2414 57776 2414 0 net8
rlabel metal1 55361 2414 55361 2414 0 net9
rlabel metal1 27600 10710 27600 10710 0 p_shaping_I.p_shaping_I.bit_in
rlabel metal1 29486 10710 29486 10710 0 p_shaping_I.p_shaping_I.bit_in_1
rlabel metal1 33350 12818 33350 12818 0 p_shaping_I.p_shaping_I.bit_in_2
rlabel metal2 28934 9860 28934 9860 0 p_shaping_I.p_shaping_I.counter\[0\]
rlabel metal1 31280 10030 31280 10030 0 p_shaping_I.p_shaping_I.counter\[1\]
rlabel metal1 27554 12274 27554 12274 0 p_shaping_I.p_shaping_I.ctl_1
rlabel metal2 19274 32674 19274 32674 0 p_shaping_Q.p_shaping_I.bit_in
rlabel metal1 22586 35632 22586 35632 0 p_shaping_Q.p_shaping_I.bit_in_1
rlabel metal2 21666 34442 21666 34442 0 p_shaping_Q.p_shaping_I.bit_in_2
rlabel metal1 28474 28526 28474 28526 0 p_shaping_Q.p_shaping_I.counter\[0\]
rlabel metal2 17802 34986 17802 34986 0 p_shaping_Q.p_shaping_I.counter\[1\]
rlabel via1 27454 31382 27454 31382 0 p_shaping_Q.p_shaping_I.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
