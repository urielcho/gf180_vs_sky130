// This is the unpowered netlist.
module OQPSK_RCOSINE_ALL (ACK,
    Bit_In,
    EN,
    REQ_SAMPLE,
    RST,
    I,
    Q,
    addI,
    addQ);
 input ACK;
 input Bit_In;
 input EN;
 input REQ_SAMPLE;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire \gen_sym.Reg_2M.data_in ;
 wire \gen_sym.Reg_2M.data_out ;
 wire \gen_sym.Reg_2M.enable ;
 wire \gen_sym.Reg_Sym.data_out[0] ;
 wire \gen_sym.Reg_Sym.data_out[1] ;
 wire \mapper.bit_Q[1] ;
 wire \p_shaping_I.p_shaping_I.bit_in ;
 wire \p_shaping_I.p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.p_shaping_I.counter[0] ;
 wire \p_shaping_I.p_shaping_I.counter[1] ;
 wire \p_shaping_I.p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in ;
 wire \p_shaping_Q.p_shaping_I.bit_in_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in_2 ;
 wire \p_shaping_Q.p_shaping_I.counter[0] ;
 wire \p_shaping_Q.p_shaping_I.counter[1] ;
 wire \p_shaping_Q.p_shaping_I.ctl_1 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;

 sky130_fd_sc_hd__clkbuf_4 _0990_ (.A(net35),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _0991_ (.A(net45),
    .X(_0828_));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(_0817_),
    .B(_0828_),
    .Y(_0839_));
 sky130_fd_sc_hd__buf_4 _0993_ (.A(net33),
    .X(_0850_));
 sky130_fd_sc_hd__a31o_1 _0994_ (.A1(_0850_),
    .A2(net32),
    .A3(net45),
    .B1(net35),
    .X(_0861_));
 sky130_fd_sc_hd__nand2b_4 _0995_ (.A_N(net36),
    .B(net37),
    .Y(_0871_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(_0839_),
    .A2(_0861_),
    .B1(_0871_),
    .Y(_0882_));
 sky130_fd_sc_hd__o21a_2 _0997_ (.A1(_0850_),
    .A2(net45),
    .B1(net35),
    .X(_0892_));
 sky130_fd_sc_hd__and2b_1 _0998_ (.A_N(net37),
    .B(net36),
    .X(_0903_));
 sky130_fd_sc_hd__o31ai_4 _0999_ (.A1(_0850_),
    .A2(net35),
    .A3(net45),
    .B1(net36),
    .Y(_0914_));
 sky130_fd_sc_hd__clkbuf_4 _1000_ (.A(net37),
    .X(_0925_));
 sky130_fd_sc_hd__a22oi_2 _1001_ (.A1(_0892_),
    .A2(_0903_),
    .B1(_0914_),
    .B2(_0925_),
    .Y(_0935_));
 sky130_fd_sc_hd__or2_1 _1002_ (.A(_0882_),
    .B(_0935_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_4 _1003_ (.A(_0850_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_4 _1004_ (.A(net45),
    .X(_0967_));
 sky130_fd_sc_hd__buf_4 _1005_ (.A(net32),
    .X(_0978_));
 sky130_fd_sc_hd__or4b_2 _1006_ (.A(_0957_),
    .B(_0817_),
    .C(_0967_),
    .D_N(_0978_),
    .X(_0989_));
 sky130_fd_sc_hd__or2_1 _1007_ (.A(_0946_),
    .B(_0989_),
    .X(_0031_));
 sky130_fd_sc_hd__buf_4 _1008_ (.A(_0031_),
    .X(_0042_));
 sky130_fd_sc_hd__clkinv_2 _1009_ (.A(_0042_),
    .Y(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _1010_ (.A(net43),
    .X(_0062_));
 sky130_fd_sc_hd__buf_2 _1011_ (.A(net41),
    .X(_0072_));
 sky130_fd_sc_hd__buf_2 _1012_ (.A(_0072_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _1013_ (.A(net40),
    .X(_0090_));
 sky130_fd_sc_hd__a21oi_1 _1014_ (.A1(_0083_),
    .A2(_0090_),
    .B1(net42),
    .Y(_0098_));
 sky130_fd_sc_hd__clkbuf_4 _1015_ (.A(net44),
    .X(_0105_));
 sky130_fd_sc_hd__buf_4 _1016_ (.A(net38),
    .X(_0112_));
 sky130_fd_sc_hd__buf_2 _1017_ (.A(net40),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_4 _1018_ (.A(net41),
    .X(_0115_));
 sky130_fd_sc_hd__a31o_2 _1019_ (.A1(_0105_),
    .A2(_0112_),
    .A3(_0114_),
    .B1(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__nand2_1 _1020_ (.A(_0098_),
    .B(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(net42),
    .Y(_0118_));
 sky130_fd_sc_hd__or3_2 _1022_ (.A(net44),
    .B(net41),
    .C(net40),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(_0118_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(net38),
    .Y(_0121_));
 sky130_fd_sc_hd__or2_1 _1025_ (.A(_0121_),
    .B(_0119_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_4 _1026_ (.A(net42),
    .X(_0123_));
 sky130_fd_sc_hd__o21a_1 _1027_ (.A1(_0105_),
    .A2(_0090_),
    .B1(_0115_),
    .X(_0124_));
 sky130_fd_sc_hd__a21oi_2 _1028_ (.A1(_0123_),
    .A2(_0124_),
    .B1(_0062_),
    .Y(_0125_));
 sky130_fd_sc_hd__a311o_4 _1029_ (.A1(_0062_),
    .A2(_0117_),
    .A3(_0120_),
    .B1(_0122_),
    .C1(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__clkinv_2 _1030_ (.A(_0126_),
    .Y(_0005_));
 sky130_fd_sc_hd__nor2b_2 _1031_ (.A(net1),
    .B_N(\gen_sym.Reg_Sym.data_out[1] ),
    .Y(_0127_));
 sky130_fd_sc_hd__buf_2 _1032_ (.A(_0127_),
    .X(\p_shaping_I.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__and2b_1 _1033_ (.A_N(net1),
    .B(\gen_sym.Reg_Sym.data_out[0] ),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(_0128_),
    .X(\mapper.bit_Q[1] ));
 sky130_fd_sc_hd__buf_2 _1035_ (.A(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(\p_shaping_I.p_shaping_I.bit_in ),
    .A1(\p_shaping_I.p_shaping_I.ctl_1 ),
    .S(net49),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(_0129_),
    .A1(_0130_),
    .S(_0042_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0131_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_2 _1039_ (.A(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_4 _1040_ (.A(\p_shaping_Q.p_shaping_I.bit_in ),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1041_ (.A0(_0133_),
    .A1(\p_shaping_Q.p_shaping_I.ctl_1 ),
    .S(net46),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(_0132_),
    .A1(_0134_),
    .S(_0126_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _1043_ (.A(_0135_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1044_ (.A(net3),
    .B(net2),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1045_ (.A(_0136_),
    .X(\gen_sym.Reg_2M.data_in ));
 sky130_fd_sc_hd__xnor2_1 _1046_ (.A(_0042_),
    .B(_0005_),
    .Y(\gen_sym.Reg_2M.enable ));
 sky130_fd_sc_hd__and2_1 _1047_ (.A(net49),
    .B(_0042_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _1048_ (.A(_0137_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1049_ (.A(net46),
    .B(_0126_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1050_ (.A(_0138_),
    .X(_0003_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(net41),
    .Y(_0139_));
 sky130_fd_sc_hd__clkbuf_4 _1052_ (.A(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_4 _1053_ (.A(net44),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_4 _1054_ (.A(net38),
    .X(_0142_));
 sky130_fd_sc_hd__nor2_4 _1055_ (.A(_0141_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__buf_2 _1056_ (.A(_0115_),
    .X(_0144_));
 sky130_fd_sc_hd__or2_2 _1057_ (.A(_0144_),
    .B(_0123_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_4 _1058_ (.A(_0062_),
    .X(_0146_));
 sky130_fd_sc_hd__a21bo_2 _1059_ (.A1(_0141_),
    .A2(net40),
    .B1_N(net41),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _1060_ (.A(_0121_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__buf_4 _1061_ (.A(net40),
    .X(_0149_));
 sky130_fd_sc_hd__a211o_1 _1062_ (.A1(_0141_),
    .A2(_0142_),
    .B1(_0072_),
    .C1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0123_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0083_),
    .B(_0062_),
    .Y(_0152_));
 sky130_fd_sc_hd__clkbuf_4 _1065_ (.A(_0114_),
    .X(_0153_));
 sky130_fd_sc_hd__o21a_1 _1066_ (.A1(_0143_),
    .A2(_0152_),
    .B1(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_4 _1067_ (.A(_0141_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2b_4 _1068_ (.A_N(_0142_),
    .B(net40),
    .Y(_0156_));
 sky130_fd_sc_hd__a31o_1 _1069_ (.A1(_0155_),
    .A2(_0144_),
    .A3(_0156_),
    .B1(_0123_),
    .X(_0157_));
 sky130_fd_sc_hd__o22a_1 _1070_ (.A1(_0148_),
    .A2(_0151_),
    .B1(_0154_),
    .B2(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a221oi_4 _1071_ (.A1(_0140_),
    .A2(_0143_),
    .B1(_0145_),
    .B2(_0146_),
    .C1(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _1072_ (.A(\p_shaping_Q.p_shaping_I.counter[1] ),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__a21oi_4 _1073_ (.A1(_0141_),
    .A2(_0112_),
    .B1(_0149_),
    .Y(_0161_));
 sky130_fd_sc_hd__or2_1 _1074_ (.A(net44),
    .B(_0142_),
    .X(_0162_));
 sky130_fd_sc_hd__and3_1 _1075_ (.A(_0141_),
    .B(_0112_),
    .C(_0149_),
    .X(_0163_));
 sky130_fd_sc_hd__a21o_1 _1076_ (.A1(_0161_),
    .A2(_0162_),
    .B1(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__nand2b_4 _1077_ (.A_N(net44),
    .B(_0149_),
    .Y(_0165_));
 sky130_fd_sc_hd__nor2_1 _1078_ (.A(_0083_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__a211o_1 _1079_ (.A1(_0144_),
    .A2(_0164_),
    .B1(_0166_),
    .C1(_0123_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_4 _1080_ (.A(_0123_),
    .X(_0168_));
 sky130_fd_sc_hd__clkinv_2 _1081_ (.A(net43),
    .Y(_0169_));
 sky130_fd_sc_hd__a21oi_1 _1082_ (.A1(_0168_),
    .A2(_0119_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__buf_2 _1083_ (.A(_0142_),
    .X(_0171_));
 sky130_fd_sc_hd__or2b_1 _1084_ (.A(_0090_),
    .B_N(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_1 _1085_ (.A(_0083_),
    .B(_0143_),
    .Y(_0173_));
 sky130_fd_sc_hd__and3_1 _1086_ (.A(_0172_),
    .B(_0156_),
    .C(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_4 _1087_ (.A(_0118_),
    .X(_0175_));
 sky130_fd_sc_hd__o21ai_2 _1088_ (.A1(_0112_),
    .A2(_0149_),
    .B1(_0072_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand2_1 _1089_ (.A(_0105_),
    .B(_0112_),
    .Y(_0177_));
 sky130_fd_sc_hd__o21a_1 _1090_ (.A1(_0112_),
    .A2(_0149_),
    .B1(_0072_),
    .X(_0178_));
 sky130_fd_sc_hd__and3_1 _1091_ (.A(_0177_),
    .B(_0165_),
    .C(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__a211o_1 _1092_ (.A1(_0175_),
    .A2(_0176_),
    .B1(_0179_),
    .C1(_0062_),
    .X(_0180_));
 sky130_fd_sc_hd__o2bb2a_2 _1093_ (.A1_N(_0167_),
    .A2_N(_0170_),
    .B1(_0174_),
    .B2(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__nor2b_2 _1094_ (.A(_0141_),
    .B_N(_0149_),
    .Y(_0182_));
 sky130_fd_sc_hd__and2b_1 _1095_ (.A_N(_0114_),
    .B(_0105_),
    .X(_0183_));
 sky130_fd_sc_hd__or3_1 _1096_ (.A(_0083_),
    .B(_0182_),
    .C(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(_0144_),
    .B(_0183_),
    .Y(_0185_));
 sky130_fd_sc_hd__o41a_1 _1098_ (.A1(_0141_),
    .A2(_0112_),
    .A3(_0072_),
    .A4(_0114_),
    .B1(net42),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _1099_ (.A(_0169_),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _1100_ (.A1(_0184_),
    .A2(_0185_),
    .B1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__nand4_1 _1101_ (.A(_0155_),
    .B(_0140_),
    .C(_0172_),
    .D(_0156_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21boi_1 _1102_ (.A1(_0105_),
    .A2(_0114_),
    .B1_N(_0072_),
    .Y(_0190_));
 sky130_fd_sc_hd__xnor2_2 _1103_ (.A(_0105_),
    .B(_0112_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0190_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__a21o_1 _1105_ (.A1(_0105_),
    .A2(_0114_),
    .B1(_0072_),
    .X(_0193_));
 sky130_fd_sc_hd__nand3_1 _1106_ (.A(_0171_),
    .B(_0115_),
    .C(_0090_),
    .Y(_0194_));
 sky130_fd_sc_hd__o211a_1 _1107_ (.A1(_0143_),
    .A2(_0193_),
    .B1(_0194_),
    .C1(_0123_),
    .X(_0195_));
 sky130_fd_sc_hd__a311o_1 _1108_ (.A1(_0175_),
    .A2(_0189_),
    .A3(_0192_),
    .B1(_0195_),
    .C1(_0146_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _1109_ (.A(_0188_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_2 _1110_ (.A(\p_shaping_Q.p_shaping_I.counter[0] ),
    .B(\p_shaping_Q.p_shaping_I.counter[1] ),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_1 _1111_ (.A(_0197_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__xnor2_1 _1112_ (.A(_0181_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__xnor2_2 _1113_ (.A(_0160_),
    .B(_0200_),
    .Y(net19));
 sky130_fd_sc_hd__a21o_1 _1114_ (.A1(_0188_),
    .A2(_0196_),
    .B1(_0132_),
    .X(_0201_));
 sky130_fd_sc_hd__buf_4 _1115_ (.A(_0169_),
    .X(_0202_));
 sky130_fd_sc_hd__and3b_1 _1116_ (.A_N(_0072_),
    .B(_0149_),
    .C(_0141_),
    .X(_0203_));
 sky130_fd_sc_hd__xor2_4 _1117_ (.A(net44),
    .B(net38),
    .X(_0204_));
 sky130_fd_sc_hd__o21ai_4 _1118_ (.A1(net44),
    .A2(_0142_),
    .B1(net40),
    .Y(_0205_));
 sky130_fd_sc_hd__o21a_1 _1119_ (.A1(_0114_),
    .A2(_0204_),
    .B1(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__o31a_1 _1120_ (.A1(_0168_),
    .A2(_0203_),
    .A3(_0206_),
    .B1(_0120_),
    .X(_0207_));
 sky130_fd_sc_hd__nor2b_2 _1121_ (.A(_0142_),
    .B_N(net44),
    .Y(_0208_));
 sky130_fd_sc_hd__o211a_1 _1122_ (.A1(_0153_),
    .A2(_0208_),
    .B1(_0156_),
    .C1(_0144_),
    .X(_0209_));
 sky130_fd_sc_hd__or2b_1 _1123_ (.A(net40),
    .B_N(net44),
    .X(_0210_));
 sky130_fd_sc_hd__a31o_1 _1124_ (.A1(_0121_),
    .A2(_0165_),
    .A3(_0210_),
    .B1(_0083_),
    .X(_0211_));
 sky130_fd_sc_hd__nor3b_1 _1125_ (.A(_0168_),
    .B(_0209_),
    .C_N(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(_0144_),
    .B(_0183_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _1127_ (.A(_0139_),
    .B(_0163_),
    .Y(_0214_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(net42),
    .B(_0062_),
    .X(_0215_));
 sky130_fd_sc_hd__o31a_1 _1129_ (.A1(_0062_),
    .A2(_0213_),
    .A3(_0214_),
    .B1(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o22a_2 _1130_ (.A1(_0202_),
    .A2(_0207_),
    .B1(_0212_),
    .B2(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _1131_ (.A(_0201_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _1132_ (.A(_0201_),
    .B(_0217_),
    .Y(_0219_));
 sky130_fd_sc_hd__or3b_1 _1133_ (.A(_0198_),
    .B(_0218_),
    .C_N(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_2 _1134_ (.A1(_0105_),
    .A2(_0149_),
    .B1(_0072_),
    .Y(_0221_));
 sky130_fd_sc_hd__and2b_1 _1135_ (.A_N(net44),
    .B(_0142_),
    .X(_0222_));
 sky130_fd_sc_hd__or3_1 _1136_ (.A(_0083_),
    .B(_0222_),
    .C(_0182_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _1137_ (.A(_0105_),
    .B(_0114_),
    .Y(_0224_));
 sky130_fd_sc_hd__o32a_1 _1138_ (.A1(_0115_),
    .A2(_0224_),
    .A3(_0204_),
    .B1(_0176_),
    .B2(_0182_),
    .X(_0225_));
 sky130_fd_sc_hd__a21oi_1 _1139_ (.A1(_0175_),
    .A2(_0225_),
    .B1(_0169_),
    .Y(_0226_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(_0083_),
    .B(_0208_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_4 _1141_ (.A(net42),
    .B(net43),
    .Y(_0228_));
 sky130_fd_sc_hd__o21a_1 _1142_ (.A1(_0214_),
    .A2(_0227_),
    .B1(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__a311o_2 _1143_ (.A1(_0168_),
    .A2(_0221_),
    .A3(_0223_),
    .B1(_0226_),
    .C1(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _1144_ (.A(\p_shaping_Q.p_shaping_I.bit_in ),
    .B(_0181_),
    .X(_0231_));
 sky130_fd_sc_hd__xnor2_1 _1145_ (.A(_0230_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__or2_1 _1146_ (.A(_0220_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__xnor2_1 _1147_ (.A(_0220_),
    .B(_0232_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .Y(_0235_));
 sky130_fd_sc_hd__buf_2 _1149_ (.A(_0083_),
    .X(_0236_));
 sky130_fd_sc_hd__or2_2 _1150_ (.A(_0153_),
    .B(_0222_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(_0144_),
    .B(_0182_),
    .Y(_0238_));
 sky130_fd_sc_hd__o22a_1 _1152_ (.A1(_0236_),
    .A2(_0237_),
    .B1(_0238_),
    .B2(_0171_),
    .X(_0239_));
 sky130_fd_sc_hd__a21o_1 _1153_ (.A1(_0141_),
    .A2(_0142_),
    .B1(net41),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_1 _1154_ (.A(_0240_),
    .B(_0205_),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2b_1 _1155_ (.A(_0090_),
    .B_N(_0112_),
    .Y(_0242_));
 sky130_fd_sc_hd__nor2_1 _1156_ (.A(_0147_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__or3_1 _1157_ (.A(_0139_),
    .B(_0118_),
    .C(_0191_),
    .X(_0244_));
 sky130_fd_sc_hd__o31a_1 _1158_ (.A1(_0168_),
    .A2(_0241_),
    .A3(_0243_),
    .B1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__a2bb2o_2 _1159_ (.A1_N(_0187_),
    .A2_N(_0239_),
    .B1(_0245_),
    .B2(_0202_),
    .X(_0246_));
 sky130_fd_sc_hd__a21o_1 _1160_ (.A1(_0235_),
    .A2(_0159_),
    .B1(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _1161_ (.A(\p_shaping_Q.p_shaping_I.counter[1] ),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__a31o_1 _1162_ (.A1(_0235_),
    .A2(_0159_),
    .A3(_0246_),
    .B1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _1163_ (.A(_0234_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_4 _1164_ (.A(_0146_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_1 _1165_ (.A(_0105_),
    .B(_0176_),
    .Y(_0252_));
 sky130_fd_sc_hd__a211o_1 _1166_ (.A1(_0123_),
    .A2(_0122_),
    .B1(_0241_),
    .C1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_2 _1167_ (.A(_0142_),
    .B(net41),
    .X(_0254_));
 sky130_fd_sc_hd__o22ai_4 _1168_ (.A1(_0114_),
    .A2(_0254_),
    .B1(_0205_),
    .B2(_0240_),
    .Y(_0255_));
 sky130_fd_sc_hd__or3_1 _1169_ (.A(net42),
    .B(_0252_),
    .C(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__nor2_1 _1170_ (.A(_0190_),
    .B(_0203_),
    .Y(_0257_));
 sky130_fd_sc_hd__o31ai_1 _1171_ (.A1(_0171_),
    .A2(_0062_),
    .A3(_0257_),
    .B1(_0215_),
    .Y(_0258_));
 sky130_fd_sc_hd__a22oi_1 _1172_ (.A1(_0251_),
    .A2(_0253_),
    .B1(_0256_),
    .B2(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__a211o_1 _1173_ (.A1(_0197_),
    .A2(_0217_),
    .B1(_0259_),
    .C1(_0132_),
    .X(_0260_));
 sky130_fd_sc_hd__a21oi_1 _1174_ (.A1(net46),
    .A2(\p_shaping_Q.p_shaping_I.ctl_1 ),
    .B1(\p_shaping_Q.p_shaping_I.bit_in ),
    .Y(_0261_));
 sky130_fd_sc_hd__and3_1 _1175_ (.A(net46),
    .B(\p_shaping_Q.p_shaping_I.bit_in ),
    .C(\p_shaping_Q.p_shaping_I.ctl_1 ),
    .X(_0262_));
 sky130_fd_sc_hd__or3_1 _1176_ (.A(_0126_),
    .B(_0261_),
    .C(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_4 _1177_ (.A(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__o211ai_1 _1178_ (.A1(_0132_),
    .A2(_0217_),
    .B1(_0201_),
    .C1(_0259_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor3_1 _1179_ (.A(_0126_),
    .B(_0261_),
    .C(_0262_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_2 _1180_ (.A(_0118_),
    .B(_0062_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21o_1 _1181_ (.A1(_0176_),
    .A2(_0211_),
    .B1(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__o21a_1 _1182_ (.A1(_0171_),
    .A2(_0147_),
    .B1(_0150_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _1183_ (.A(_0228_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_2 _1184_ (.A(_0115_),
    .B(_0156_),
    .Y(_0271_));
 sky130_fd_sc_hd__a211o_1 _1185_ (.A1(_0090_),
    .A2(_0222_),
    .B1(_0208_),
    .C1(_0115_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(net42),
    .B(_0169_),
    .Y(_0273_));
 sky130_fd_sc_hd__a211o_1 _1187_ (.A1(_0271_),
    .A2(_0272_),
    .B1(_0273_),
    .C1(_0269_),
    .X(_0274_));
 sky130_fd_sc_hd__a31o_1 _1188_ (.A1(_0268_),
    .A2(_0270_),
    .A3(_0274_),
    .B1(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .X(_0275_));
 sky130_fd_sc_hd__a221o_1 _1189_ (.A1(_0146_),
    .A2(_0253_),
    .B1(_0256_),
    .B2(_0258_),
    .C1(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .X(_0276_));
 sky130_fd_sc_hd__a211o_1 _1190_ (.A1(_0144_),
    .A2(_0206_),
    .B1(_0186_),
    .C1(_0166_),
    .X(_0277_));
 sky130_fd_sc_hd__a21o_1 _1191_ (.A1(_0090_),
    .A2(_0204_),
    .B1(_0221_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_2 _1192_ (.A(_0112_),
    .B(_0149_),
    .Y(_0279_));
 sky130_fd_sc_hd__a31o_1 _1193_ (.A1(_0165_),
    .A2(_0210_),
    .A3(_0279_),
    .B1(_0115_),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _1194_ (.A1(_0278_),
    .A2(_0280_),
    .B1(_0123_),
    .X(_0281_));
 sky130_fd_sc_hd__o21ai_1 _1195_ (.A1(_0115_),
    .A2(_0279_),
    .B1(net42),
    .Y(_0282_));
 sky130_fd_sc_hd__o21a_1 _1196_ (.A1(_0148_),
    .A2(_0282_),
    .B1(_0169_),
    .X(_0283_));
 sky130_fd_sc_hd__a221o_1 _1197_ (.A1(_0146_),
    .A2(_0277_),
    .B1(_0281_),
    .B2(_0283_),
    .C1(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .X(_0284_));
 sky130_fd_sc_hd__a41o_1 _1198_ (.A1(_0266_),
    .A2(_0275_),
    .A3(_0276_),
    .A4(_0284_),
    .B1(_0198_),
    .X(_0285_));
 sky130_fd_sc_hd__a31o_1 _1199_ (.A1(_0260_),
    .A2(_0264_),
    .A3(_0265_),
    .B1(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__a21oi_1 _1200_ (.A1(_0181_),
    .A2(_0230_),
    .B1(_0133_),
    .Y(_0287_));
 sky130_fd_sc_hd__nor2_1 _1201_ (.A(_0222_),
    .B(_0242_),
    .Y(_0288_));
 sky130_fd_sc_hd__or2_1 _1202_ (.A(_0155_),
    .B(_0121_),
    .X(_0289_));
 sky130_fd_sc_hd__o2bb2a_1 _1203_ (.A1_N(_0288_),
    .A2_N(_0254_),
    .B1(_0144_),
    .B2(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__o221a_1 _1204_ (.A1(_0271_),
    .A2(_0182_),
    .B1(_0204_),
    .B2(_0153_),
    .C1(_0169_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _1205_ (.A(_0155_),
    .B(_0090_),
    .X(_0292_));
 sky130_fd_sc_hd__a31o_1 _1206_ (.A1(_0171_),
    .A2(_0292_),
    .A3(_0257_),
    .B1(_0215_),
    .X(_0293_));
 sky130_fd_sc_hd__o221ai_4 _1207_ (.A1(_0202_),
    .A2(_0290_),
    .B1(_0291_),
    .B2(_0175_),
    .C1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__xnor2_1 _1208_ (.A(_0287_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__xor2_1 _1209_ (.A(_0286_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__or2_1 _1210_ (.A(_0159_),
    .B(_0246_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _1211_ (.A(_0153_),
    .X(_0298_));
 sky130_fd_sc_hd__o31a_1 _1212_ (.A1(_0236_),
    .A2(_0298_),
    .A3(_0208_),
    .B1(_0194_),
    .X(_0299_));
 sky130_fd_sc_hd__nor2b_1 _1213_ (.A(_0153_),
    .B_N(_0083_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _1214_ (.A(_0177_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__a211o_1 _1215_ (.A1(_0161_),
    .A2(_0254_),
    .B1(_0273_),
    .C1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _1216_ (.A(_0236_),
    .B(_0298_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _1217_ (.A(_0140_),
    .B(_0279_),
    .Y(_0304_));
 sky130_fd_sc_hd__o2111ai_4 _1218_ (.A1(_0289_),
    .A2(_0303_),
    .B1(_0237_),
    .C1(_0228_),
    .D1(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o211ai_4 _1219_ (.A1(_0267_),
    .A2(_0299_),
    .B1(_0302_),
    .C1(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__a21oi_1 _1220_ (.A1(_0235_),
    .A2(_0297_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__and3_1 _1221_ (.A(_0235_),
    .B(_0297_),
    .C(_0306_),
    .X(_0308_));
 sky130_fd_sc_hd__or3b_1 _1222_ (.A(_0307_),
    .B(_0308_),
    .C_N(\p_shaping_Q.p_shaping_I.counter[1] ),
    .X(_0309_));
 sky130_fd_sc_hd__xor2_1 _1223_ (.A(_0296_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__a21bo_1 _1224_ (.A1(_0233_),
    .A2(_0250_),
    .B1_N(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__nand3b_1 _1225_ (.A_N(_0310_),
    .B(_0233_),
    .C(_0250_),
    .Y(_0312_));
 sky130_fd_sc_hd__or2b_1 _1226_ (.A(_0160_),
    .B_N(_0200_),
    .X(_0313_));
 sky130_fd_sc_hd__o31ai_1 _1227_ (.A1(_0181_),
    .A2(_0197_),
    .A3(_0198_),
    .B1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__xor2_1 _1228_ (.A(_0234_),
    .B(_0249_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(_0314_),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__and3_1 _1230_ (.A(_0311_),
    .B(_0312_),
    .C(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__a21oi_1 _1231_ (.A1(_0311_),
    .A2(_0312_),
    .B1(_0316_),
    .Y(_0318_));
 sky130_fd_sc_hd__nor2_1 _1232_ (.A(_0317_),
    .B(_0318_),
    .Y(net24));
 sky130_fd_sc_hd__and2b_1 _1233_ (.A_N(_0286_),
    .B(_0295_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0296_),
    .B(_0309_),
    .Y(_0320_));
 sky130_fd_sc_hd__a22o_1 _1235_ (.A1(_0251_),
    .A2(_0277_),
    .B1(_0281_),
    .B2(_0283_),
    .X(_0321_));
 sky130_fd_sc_hd__o211a_1 _1236_ (.A1(_0132_),
    .A2(_0217_),
    .B1(_0276_),
    .C1(_0201_),
    .X(_0322_));
 sky130_fd_sc_hd__xnor2_1 _1237_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__a21o_1 _1238_ (.A1(_0155_),
    .A2(_0171_),
    .B1(_0153_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _1239_ (.A(_0236_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__a22o_1 _1240_ (.A1(_0146_),
    .A2(_0145_),
    .B1(_0228_),
    .B2(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _1241_ (.A(_0132_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a41o_1 _1242_ (.A1(_0275_),
    .A2(_0276_),
    .A3(_0284_),
    .A4(_0326_),
    .B1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__inv_2 _1243_ (.A(_0198_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21ai_2 _1244_ (.A1(_0264_),
    .A2(_0328_),
    .B1(_0007_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21oi_1 _1245_ (.A1(_0264_),
    .A2(_0323_),
    .B1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__a31o_1 _1246_ (.A1(_0181_),
    .A2(_0230_),
    .A3(_0294_),
    .B1(_0133_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(_0090_),
    .B(_0204_),
    .Y(_0332_));
 sky130_fd_sc_hd__a221o_1 _1248_ (.A1(_0204_),
    .A2(_0178_),
    .B1(_0332_),
    .B2(_0140_),
    .C1(_0123_),
    .X(_0333_));
 sky130_fd_sc_hd__or3b_1 _1249_ (.A(_0072_),
    .B(_0208_),
    .C_N(_0114_),
    .X(_0334_));
 sky130_fd_sc_hd__and3b_1 _1250_ (.A_N(_0148_),
    .B(_0228_),
    .C(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__or2_2 _1251_ (.A(_0090_),
    .B(_0162_),
    .X(_0336_));
 sky130_fd_sc_hd__nor2_1 _1252_ (.A(_0118_),
    .B(_0062_),
    .Y(_0337_));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(_0143_),
    .A1(_0156_),
    .S(_0115_),
    .X(_0338_));
 sky130_fd_sc_hd__and3_1 _1254_ (.A(_0336_),
    .B(_0337_),
    .C(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__a311o_1 _1255_ (.A1(_0146_),
    .A2(_0122_),
    .A3(_0333_),
    .B1(_0335_),
    .C1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__xor2_1 _1256_ (.A(_0331_),
    .B(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__xor2_1 _1257_ (.A(_0330_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _1258_ (.A(_0297_),
    .B(_0306_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _1259_ (.A1(_0153_),
    .A2(_0204_),
    .B1(_0242_),
    .Y(_0344_));
 sky130_fd_sc_hd__and2_1 _1260_ (.A(_0223_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o21bai_1 _1261_ (.A1(_0223_),
    .A2(_0344_),
    .B1_N(_0267_),
    .Y(_0346_));
 sky130_fd_sc_hd__o21ai_1 _1262_ (.A1(_0242_),
    .A2(_0193_),
    .B1(_0228_),
    .Y(_0347_));
 sky130_fd_sc_hd__a31o_1 _1263_ (.A1(_0165_),
    .A2(_0164_),
    .A3(_0178_),
    .B1(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__or3b_1 _1264_ (.A(_0182_),
    .B(_0183_),
    .C_N(_0279_),
    .X(_0349_));
 sky130_fd_sc_hd__and3_1 _1265_ (.A(_0144_),
    .B(_0165_),
    .C(_0279_),
    .X(_0350_));
 sky130_fd_sc_hd__a221o_1 _1266_ (.A1(_0173_),
    .A2(_0349_),
    .B1(_0350_),
    .B2(_0210_),
    .C1(_0273_),
    .X(_0351_));
 sky130_fd_sc_hd__o211a_1 _1267_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0348_),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__o21ai_1 _1268_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .A2(_0343_),
    .B1(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__or3_1 _1269_ (.A(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .B(_0352_),
    .C(_0343_),
    .X(_0354_));
 sky130_fd_sc_hd__and3_1 _1270_ (.A(\p_shaping_Q.p_shaping_I.counter[1] ),
    .B(_0353_),
    .C(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__xor2_1 _1271_ (.A(_0342_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _1272_ (.A1(_0319_),
    .A2(_0320_),
    .B1(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__or3_1 _1273_ (.A(_0319_),
    .B(_0320_),
    .C(_0356_),
    .X(_0358_));
 sky130_fd_sc_hd__and2b_1 _1274_ (.A_N(_0357_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__a21bo_1 _1275_ (.A1(_0312_),
    .A2(_0316_),
    .B1_N(_0311_),
    .X(_0360_));
 sky130_fd_sc_hd__xor2_4 _1276_ (.A(_0359_),
    .B(_0360_),
    .X(net25));
 sky130_fd_sc_hd__a21oi_1 _1277_ (.A1(_0358_),
    .A2(_0360_),
    .B1(_0357_),
    .Y(_0361_));
 sky130_fd_sc_hd__buf_2 _1278_ (.A(\p_shaping_Q.p_shaping_I.counter[1] ),
    .X(_0362_));
 sky130_fd_sc_hd__o211ai_2 _1279_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0348_),
    .C1(_0351_),
    .Y(_0363_));
 sky130_fd_sc_hd__o41ai_4 _1280_ (.A1(_0159_),
    .A2(_0246_),
    .A3(_0306_),
    .A4(_0363_),
    .B1(_0235_),
    .Y(_0364_));
 sky130_fd_sc_hd__buf_2 _1281_ (.A(_0236_),
    .X(_0365_));
 sky130_fd_sc_hd__o211a_1 _1282_ (.A1(_0298_),
    .A2(_0177_),
    .B1(_0162_),
    .C1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a211o_1 _1283_ (.A1(_0124_),
    .A2(_0288_),
    .B1(_0255_),
    .C1(_0175_),
    .X(_0367_));
 sky130_fd_sc_hd__buf_2 _1284_ (.A(_0168_),
    .X(_0368_));
 sky130_fd_sc_hd__a311o_1 _1285_ (.A1(_0155_),
    .A2(_0171_),
    .A3(_0236_),
    .B1(_0368_),
    .C1(_0203_),
    .X(_0369_));
 sky130_fd_sc_hd__nand3_1 _1286_ (.A(_0202_),
    .B(_0367_),
    .C(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__o31a_2 _1287_ (.A1(_0267_),
    .A2(_0241_),
    .A3(_0366_),
    .B1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__xor2_1 _1288_ (.A(_0364_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__o21a_1 _1289_ (.A1(_0132_),
    .A2(_0217_),
    .B1(_0201_),
    .X(_0373_));
 sky130_fd_sc_hd__and2_1 _1290_ (.A(_0276_),
    .B(_0284_),
    .X(_0374_));
 sky130_fd_sc_hd__a221o_1 _1291_ (.A1(_0236_),
    .A2(_0164_),
    .B1(_0205_),
    .B2(_0292_),
    .C1(_0168_),
    .X(_0375_));
 sky130_fd_sc_hd__and2b_1 _1292_ (.A_N(_0186_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _1293_ (.A(_0155_),
    .B(_0300_),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _1294_ (.A1(_0254_),
    .A2(_0210_),
    .B1(_0337_),
    .C1(_0289_),
    .X(_0378_));
 sky130_fd_sc_hd__a31o_1 _1295_ (.A1(_0185_),
    .A2(_0228_),
    .A3(_0377_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__a21o_1 _1296_ (.A1(_0251_),
    .A2(_0376_),
    .B1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__and3_1 _1297_ (.A(_0373_),
    .B(_0374_),
    .C(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__a21oi_1 _1298_ (.A1(_0373_),
    .A2(_0374_),
    .B1(_0380_),
    .Y(_0382_));
 sky130_fd_sc_hd__o21a_1 _1299_ (.A1(_0264_),
    .A2(_0328_),
    .B1(_0007_),
    .X(_0383_));
 sky130_fd_sc_hd__o31a_1 _1300_ (.A1(_0266_),
    .A2(_0381_),
    .A3(_0382_),
    .B1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__and4_1 _1301_ (.A(_0181_),
    .B(_0230_),
    .C(_0294_),
    .D(_0340_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _1302_ (.A(_0133_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a31o_1 _1303_ (.A1(_0236_),
    .A2(_0165_),
    .A3(_0336_),
    .B1(_0282_),
    .X(_0387_));
 sky130_fd_sc_hd__nand3_1 _1304_ (.A(_0155_),
    .B(_0175_),
    .C(_0193_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _1305_ (.A1(_0324_),
    .A2(_0205_),
    .B1(_0140_),
    .Y(_0389_));
 sky130_fd_sc_hd__o21ba_1 _1306_ (.A1(_0171_),
    .A2(_0153_),
    .B1_N(_0240_),
    .X(_0390_));
 sky130_fd_sc_hd__o31a_1 _1307_ (.A1(_0168_),
    .A2(_0389_),
    .A3(_0390_),
    .B1(_0146_),
    .X(_0391_));
 sky130_fd_sc_hd__a31o_1 _1308_ (.A1(_0202_),
    .A2(_0387_),
    .A3(_0388_),
    .B1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__xnor2_1 _1309_ (.A(_0386_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__xor2_1 _1310_ (.A(_0384_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a21oi_1 _1311_ (.A1(_0362_),
    .A2(_0372_),
    .B1(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__and3_1 _1312_ (.A(_0362_),
    .B(_0394_),
    .C(_0372_),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _1313_ (.A(_0395_),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _1314_ (.A(_0330_),
    .B(_0341_),
    .X(_0398_));
 sky130_fd_sc_hd__a21oi_2 _1315_ (.A1(_0342_),
    .A2(_0355_),
    .B1(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__xor2_1 _1316_ (.A(_0397_),
    .B(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__and2b_1 _1317_ (.A_N(_0361_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__and2b_1 _1318_ (.A_N(_0400_),
    .B(_0361_),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_2 _1319_ (.A(_0401_),
    .B(_0402_),
    .Y(net26));
 sky130_fd_sc_hd__and2_1 _1320_ (.A(_0384_),
    .B(_0393_),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _1321_ (.A(_0268_),
    .B(_0270_),
    .C(_0274_),
    .X(_0404_));
 sky130_fd_sc_hd__a21bo_1 _1322_ (.A1(_0404_),
    .A2(_0374_),
    .B1_N(_0275_),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _1323_ (.A1(_0264_),
    .A2(_0405_),
    .B1(_0329_),
    .X(_0406_));
 sky130_fd_sc_hd__a21o_1 _1324_ (.A1(_0385_),
    .A2(_0392_),
    .B1(_0133_),
    .X(_0407_));
 sky130_fd_sc_hd__nor3_1 _1325_ (.A(_0175_),
    .B(_0203_),
    .C(_0209_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _1326_ (.A(_0368_),
    .B(_0300_),
    .Y(_0409_));
 sky130_fd_sc_hd__and2_1 _1327_ (.A(_0236_),
    .B(_0153_),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _1328_ (.A(_0140_),
    .B(_0177_),
    .C(_0279_),
    .X(_0411_));
 sky130_fd_sc_hd__o21a_1 _1329_ (.A1(_0410_),
    .A2(_0411_),
    .B1(_0336_),
    .X(_0412_));
 sky130_fd_sc_hd__o32a_1 _1330_ (.A1(_0146_),
    .A2(_0408_),
    .A3(_0409_),
    .B1(_0187_),
    .B2(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__xnor2_1 _1331_ (.A(_0407_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__xnor2_1 _1332_ (.A(_0406_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__o32a_1 _1333_ (.A1(_0224_),
    .A2(_0143_),
    .A3(_0193_),
    .B1(_0204_),
    .B2(_0147_),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _1334_ (.A(_0146_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0116_),
    .B(_0325_),
    .Y(_0418_));
 sky130_fd_sc_hd__a22o_1 _1336_ (.A1(_0368_),
    .A2(_0417_),
    .B1(_0418_),
    .B2(_0251_),
    .X(_0419_));
 sky130_fd_sc_hd__a31o_1 _1337_ (.A1(_0271_),
    .A2(_0189_),
    .A3(_0228_),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__o21a_1 _1338_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .A2(_0371_),
    .B1(_0364_),
    .X(_0421_));
 sky130_fd_sc_hd__a21boi_1 _1339_ (.A1(_0420_),
    .A2(_0421_),
    .B1_N(\p_shaping_Q.p_shaping_I.counter[1] ),
    .Y(_0422_));
 sky130_fd_sc_hd__o21a_1 _1340_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__xnor2_1 _1341_ (.A(_0415_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_1 _1342_ (.A1(_0403_),
    .A2(_0396_),
    .B1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__or3_1 _1343_ (.A(_0403_),
    .B(_0396_),
    .C(_0424_),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _1344_ (.A(_0425_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__o21ba_1 _1345_ (.A1(_0397_),
    .A2(_0399_),
    .B1_N(_0401_),
    .X(_0428_));
 sky130_fd_sc_hd__xnor2_2 _1346_ (.A(_0427_),
    .B(_0428_),
    .Y(net27));
 sky130_fd_sc_hd__and3_1 _1347_ (.A(_0275_),
    .B(_0276_),
    .C(_0284_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_2 _1348_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _1349_ (.A(_0298_),
    .B(_0191_),
    .Y(_0431_));
 sky130_fd_sc_hd__nor2_1 _1350_ (.A(_0163_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__o21a_1 _1351_ (.A1(_0140_),
    .A2(_0164_),
    .B1(_0288_),
    .X(_0433_));
 sky130_fd_sc_hd__a211o_1 _1352_ (.A1(_0148_),
    .A2(_0432_),
    .B1(_0433_),
    .C1(_0368_),
    .X(_0434_));
 sky130_fd_sc_hd__a311o_1 _1353_ (.A1(_0368_),
    .A2(_0237_),
    .A3(_0205_),
    .B1(_0156_),
    .C1(_0365_),
    .X(_0435_));
 sky130_fd_sc_hd__o2111ai_1 _1354_ (.A1(_0236_),
    .A2(_0156_),
    .B1(_0237_),
    .C1(_0205_),
    .D1(_0168_),
    .Y(_0436_));
 sky130_fd_sc_hd__o311a_1 _1355_ (.A1(_0368_),
    .A2(_0271_),
    .A3(_0332_),
    .B1(_0436_),
    .C1(_0202_),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _1356_ (.A1(_0251_),
    .A2(_0434_),
    .B1(_0435_),
    .B2(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__xnor2_1 _1357_ (.A(_0430_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1358_ (.A1(_0264_),
    .A2(_0439_),
    .B1(_0329_),
    .Y(_0440_));
 sky130_fd_sc_hd__a21o_1 _1359_ (.A1(_0298_),
    .A2(_0191_),
    .B1(_0221_),
    .X(_0441_));
 sky130_fd_sc_hd__a31o_1 _1360_ (.A1(_0368_),
    .A2(_0193_),
    .A3(_0441_),
    .B1(_0098_),
    .X(_0442_));
 sky130_fd_sc_hd__a21o_1 _1361_ (.A1(_0271_),
    .A2(_0272_),
    .B1(_0267_),
    .X(_0443_));
 sky130_fd_sc_hd__o21a_1 _1362_ (.A1(_0251_),
    .A2(_0442_),
    .B1(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a31o_2 _1363_ (.A1(_0385_),
    .A2(_0392_),
    .A3(_0413_),
    .B1(_0133_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _1364_ (.A(_0133_),
    .B(_0444_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21oi_1 _1365_ (.A1(_0444_),
    .A2(_0445_),
    .B1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__xor2_1 _1366_ (.A(_0440_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_2 _1367_ (.A(_0368_),
    .X(_0449_));
 sky130_fd_sc_hd__and3_1 _1368_ (.A(_0368_),
    .B(_0336_),
    .C(_0205_),
    .X(_0450_));
 sky130_fd_sc_hd__xnor2_1 _1369_ (.A(_0411_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__buf_2 _1370_ (.A(_0251_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_1 _1371_ (.A1(_0449_),
    .A2(_0116_),
    .B1(_0251_),
    .Y(_0453_));
 sky130_fd_sc_hd__o221a_1 _1372_ (.A1(_0449_),
    .A2(_0238_),
    .B1(_0451_),
    .B2(_0452_),
    .C1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__a31o_2 _1373_ (.A1(_0364_),
    .A2(_0371_),
    .A3(_0420_),
    .B1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .X(_0455_));
 sky130_fd_sc_hd__xnor2_1 _1374_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _1375_ (.A(\p_shaping_Q.p_shaping_I.counter[1] ),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__xor2_1 _1376_ (.A(_0448_),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__nand2_1 _1377_ (.A(_0406_),
    .B(_0414_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_0406_),
    .B(_0414_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _1379_ (.A1(_0459_),
    .A2(_0423_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__xnor2_1 _1380_ (.A(_0458_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nor3_1 _1381_ (.A(_0403_),
    .B(_0396_),
    .C(_0424_),
    .Y(_0463_));
 sky130_fd_sc_hd__o31a_1 _1382_ (.A1(_0397_),
    .A2(_0399_),
    .A3(_0463_),
    .B1(_0425_),
    .X(_0464_));
 sky130_fd_sc_hd__a21bo_1 _1383_ (.A1(_0401_),
    .A2(_0427_),
    .B1_N(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__xnor2_2 _1384_ (.A(_0462_),
    .B(_0465_),
    .Y(net28));
 sky130_fd_sc_hd__nand2_1 _1385_ (.A(_0298_),
    .B(_0204_),
    .Y(_0466_));
 sky130_fd_sc_hd__o211a_1 _1386_ (.A1(_0208_),
    .A2(_0237_),
    .B1(_0466_),
    .C1(_0140_),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_1 _1387_ (.A1(_0350_),
    .A2(_0467_),
    .B1(_0337_),
    .Y(_0468_));
 sky130_fd_sc_hd__xnor2_1 _1388_ (.A(_0155_),
    .B(_0271_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(_0168_),
    .B(_0122_),
    .Y(_0470_));
 sky130_fd_sc_hd__or3b_1 _1390_ (.A(_0469_),
    .B(_0202_),
    .C_N(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a31o_1 _1391_ (.A1(_0365_),
    .A2(_0336_),
    .A3(_0466_),
    .B1(_0347_),
    .X(_0472_));
 sky130_fd_sc_hd__a31o_1 _1392_ (.A1(_0468_),
    .A2(_0471_),
    .A3(_0472_),
    .B1(_0266_),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_1 _1393_ (.A(_0132_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__a211o_1 _1394_ (.A1(_0430_),
    .A2(_0473_),
    .B1(_0474_),
    .C1(_0198_),
    .X(_0475_));
 sky130_fd_sc_hd__o2111a_1 _1395_ (.A1(_0116_),
    .A2(_0161_),
    .B1(_0470_),
    .C1(_0238_),
    .D1(_0251_),
    .X(_0476_));
 sky130_fd_sc_hd__a31o_1 _1396_ (.A1(_0124_),
    .A2(_0205_),
    .A3(_0337_),
    .B1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__xor2_2 _1397_ (.A(_0445_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__xor2_2 _1398_ (.A(_0475_),
    .B(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _1399_ (.A(_0365_),
    .B(_0336_),
    .X(_0480_));
 sky130_fd_sc_hd__a211o_1 _1400_ (.A1(_0171_),
    .A2(_0183_),
    .B1(_0182_),
    .C1(_0175_),
    .X(_0481_));
 sky130_fd_sc_hd__o32a_1 _1401_ (.A1(_0449_),
    .A2(_0410_),
    .A3(_0255_),
    .B1(_0480_),
    .B2(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_1 _1402_ (.A(_0452_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__xnor2_1 _1403_ (.A(_0455_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_0362_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__xor2_2 _1405_ (.A(_0479_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__and2_1 _1406_ (.A(_0440_),
    .B(_0447_),
    .X(_0487_));
 sky130_fd_sc_hd__a31o_1 _1407_ (.A1(_0362_),
    .A2(_0448_),
    .A3(_0456_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__xor2_2 _1408_ (.A(_0486_),
    .B(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _1409_ (.A(_0458_),
    .B(_0461_),
    .Y(_0490_));
 sky130_fd_sc_hd__or2_1 _1410_ (.A(_0458_),
    .B(_0461_),
    .X(_0491_));
 sky130_fd_sc_hd__a21bo_1 _1411_ (.A1(_0490_),
    .A2(_0465_),
    .B1_N(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__xnor2_2 _1412_ (.A(_0489_),
    .B(_0492_),
    .Y(net29));
 sky130_fd_sc_hd__a21oi_1 _1413_ (.A1(_0324_),
    .A2(_0205_),
    .B1(_0365_),
    .Y(_0493_));
 sky130_fd_sc_hd__or2_1 _1414_ (.A(_0157_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__a41o_1 _1415_ (.A1(_0385_),
    .A2(_0392_),
    .A3(_0413_),
    .A4(_0494_),
    .B1(_0133_),
    .X(_0495_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(_0133_),
    .Y(_0496_));
 sky130_fd_sc_hd__a31oi_1 _1417_ (.A1(_0452_),
    .A2(_0117_),
    .A3(_0120_),
    .B1(_0125_),
    .Y(_0497_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(_0495_),
    .A1(_0496_),
    .S(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__and3_1 _1419_ (.A(_0165_),
    .B(_0178_),
    .C(_0279_),
    .X(_0499_));
 sky130_fd_sc_hd__or3_1 _1420_ (.A(_0186_),
    .B(_0467_),
    .C(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a211o_1 _1421_ (.A1(_0213_),
    .A2(_0466_),
    .B1(_0499_),
    .C1(_0368_),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(_0172_),
    .B(_0173_),
    .Y(_0502_));
 sky130_fd_sc_hd__a31o_1 _1423_ (.A1(_0202_),
    .A2(_0147_),
    .A3(_0502_),
    .B1(_0228_),
    .X(_0503_));
 sky130_fd_sc_hd__a22oi_2 _1424_ (.A1(_0251_),
    .A2(_0500_),
    .B1(_0501_),
    .B2(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__or2_1 _1425_ (.A(_0430_),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _1426_ (.A(_0132_),
    .B(_0504_),
    .Y(_0506_));
 sky130_fd_sc_hd__a31o_1 _1427_ (.A1(_0264_),
    .A2(_0505_),
    .A3(_0506_),
    .B1(_0329_),
    .X(_0507_));
 sky130_fd_sc_hd__or2_1 _1428_ (.A(_0498_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_0498_),
    .B(_0507_),
    .Y(_0509_));
 sky130_fd_sc_hd__and2_1 _1430_ (.A(_0508_),
    .B(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__mux4_1 _1431_ (.A0(_0298_),
    .A1(_0432_),
    .A2(_0336_),
    .A3(_0161_),
    .S0(_0140_),
    .S1(_0449_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_1 _1432_ (.A(_0452_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__inv_2 _1433_ (.A(_0376_),
    .Y(_0513_));
 sky130_fd_sc_hd__o211ai_1 _1434_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .A2(_0513_),
    .B1(_0455_),
    .C1(_0512_),
    .Y(_0514_));
 sky130_fd_sc_hd__o211a_1 _1435_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .A2(_0512_),
    .B1(_0514_),
    .C1(_0362_),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _1436_ (.A(_0510_),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(_0510_),
    .B(_0515_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_2 _1438_ (.A(_0516_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand3_1 _1439_ (.A(_0362_),
    .B(_0479_),
    .C(_0484_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_2 _1440_ (.A1(_0475_),
    .A2(_0478_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__xor2_4 _1441_ (.A(_0518_),
    .B(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__and2b_1 _1442_ (.A_N(_0488_),
    .B(_0486_),
    .X(_0522_));
 sky130_fd_sc_hd__or2b_1 _1443_ (.A(_0486_),
    .B_N(_0488_),
    .X(_0523_));
 sky130_fd_sc_hd__o21a_1 _1444_ (.A1(_0491_),
    .A2(_0522_),
    .B1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__or2_1 _1445_ (.A(_0462_),
    .B(_0489_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _1446_ (.A(_0464_),
    .B(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_1 _1447_ (.A(_0425_),
    .B(_0426_),
    .Y(_0527_));
 sky130_fd_sc_hd__or4b_1 _1448_ (.A(_0361_),
    .B(_0527_),
    .C(_0525_),
    .D_N(_0400_),
    .X(_0528_));
 sky130_fd_sc_hd__and3_1 _1449_ (.A(_0524_),
    .B(_0526_),
    .C(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__xor2_4 _1450_ (.A(_0521_),
    .B(_0529_),
    .X(net30));
 sky130_fd_sc_hd__nand2_1 _1451_ (.A(_0508_),
    .B(_0517_),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _1452_ (.A(_0147_),
    .B(_0431_),
    .Y(_0531_));
 sky130_fd_sc_hd__a31o_1 _1453_ (.A1(_0140_),
    .A2(_0156_),
    .A3(_0165_),
    .B1(_0449_),
    .X(_0532_));
 sky130_fd_sc_hd__o211a_1 _1454_ (.A1(_0531_),
    .A2(_0532_),
    .B1(_0202_),
    .C1(_0151_),
    .X(_0533_));
 sky130_fd_sc_hd__a21oi_1 _1455_ (.A1(_0452_),
    .A2(_0494_),
    .B1(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__or2_1 _1456_ (.A(_0430_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(_0132_),
    .B(_0534_),
    .Y(_0536_));
 sky130_fd_sc_hd__a31o_1 _1458_ (.A1(_0264_),
    .A2(_0535_),
    .A3(_0536_),
    .B1(_0329_),
    .X(_0537_));
 sky130_fd_sc_hd__clkinv_2 _1459_ (.A(_0445_),
    .Y(_0538_));
 sky130_fd_sc_hd__a31o_1 _1460_ (.A1(_0452_),
    .A2(_0303_),
    .A3(_0116_),
    .B1(_0125_),
    .X(_0539_));
 sky130_fd_sc_hd__a31o_1 _1461_ (.A1(_0449_),
    .A2(_0452_),
    .A3(_0119_),
    .B1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(_0133_),
    .A1(_0538_),
    .S(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__xnor2_1 _1463_ (.A(_0537_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__o21ai_1 _1464_ (.A1(_0365_),
    .A2(_0177_),
    .B1(_0298_),
    .Y(_0543_));
 sky130_fd_sc_hd__o311a_1 _1465_ (.A1(_0365_),
    .A2(_0298_),
    .A3(_0143_),
    .B1(_0543_),
    .C1(_0175_),
    .X(_0544_));
 sky130_fd_sc_hd__a31o_1 _1466_ (.A1(_0365_),
    .A2(_0449_),
    .A3(_0336_),
    .B1(_0452_),
    .X(_0545_));
 sky130_fd_sc_hd__o21ai_1 _1467_ (.A1(_0544_),
    .A2(_0545_),
    .B1(_0455_),
    .Y(_0546_));
 sky130_fd_sc_hd__or3_1 _1468_ (.A(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .B(_0544_),
    .C(_0545_),
    .X(_0547_));
 sky130_fd_sc_hd__nand4_2 _1469_ (.A(_0362_),
    .B(_0542_),
    .C(_0546_),
    .D(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a31o_1 _1470_ (.A1(_0362_),
    .A2(_0546_),
    .A3(_0547_),
    .B1(_0542_),
    .X(_0549_));
 sky130_fd_sc_hd__and3_1 _1471_ (.A(_0530_),
    .B(_0548_),
    .C(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0548_),
    .B(_0549_),
    .Y(_0551_));
 sky130_fd_sc_hd__and3_1 _1473_ (.A(_0508_),
    .B(_0517_),
    .C(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _1474_ (.A(_0550_),
    .B(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__or2b_1 _1475_ (.A(_0518_),
    .B_N(_0520_),
    .X(_0554_));
 sky130_fd_sc_hd__a31o_1 _1476_ (.A1(_0524_),
    .A2(_0526_),
    .A3(_0528_),
    .B1(_0521_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _1477_ (.A(_0554_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__xnor2_2 _1478_ (.A(_0553_),
    .B(_0556_),
    .Y(net31));
 sky130_fd_sc_hd__or2b_1 _1479_ (.A(_0551_),
    .B_N(_0530_),
    .X(_0557_));
 sky130_fd_sc_hd__and2_1 _1480_ (.A(_0554_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__or2b_1 _1481_ (.A(_0537_),
    .B_N(_0541_),
    .X(_0559_));
 sky130_fd_sc_hd__xnor2_1 _1482_ (.A(_0264_),
    .B(_0430_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_1 _1483_ (.A1(_0300_),
    .A2(_0161_),
    .B1(_0175_),
    .Y(_0561_));
 sky130_fd_sc_hd__a22o_1 _1484_ (.A1(_0228_),
    .A2(_0418_),
    .B1(_0561_),
    .B2(_0452_),
    .X(_0562_));
 sky130_fd_sc_hd__xor2_1 _1485_ (.A(_0560_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(_0007_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__a31o_1 _1487_ (.A1(_0449_),
    .A2(_0452_),
    .A3(_0119_),
    .B1(_0496_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(_0565_),
    .A1(_0445_),
    .S(_0125_),
    .X(_0566_));
 sky130_fd_sc_hd__xor2_1 _1489_ (.A(_0564_),
    .B(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_1 _1490_ (.A(_0145_),
    .B(_0336_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_1 _1491_ (.A1(_0545_),
    .A2(_0568_),
    .B1(_0455_),
    .Y(_0569_));
 sky130_fd_sc_hd__o311a_1 _1492_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .A2(_0545_),
    .A3(_0568_),
    .B1(_0569_),
    .C1(_0362_),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(_0567_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__or2_1 _1494_ (.A(_0567_),
    .B(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _1495_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__a21o_1 _1496_ (.A1(_0559_),
    .A2(_0548_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__nand3_1 _1497_ (.A(_0559_),
    .B(_0548_),
    .C(_0573_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a211o_1 _1499_ (.A1(_0555_),
    .A2(_0558_),
    .B1(_0576_),
    .C1(_0552_),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_1 _1500_ (.A1(_0555_),
    .A2(_0558_),
    .B1(_0552_),
    .X(_0578_));
 sky130_fd_sc_hd__nand2_1 _1501_ (.A(_0576_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__and2_1 _1502_ (.A(_0577_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _1503_ (.A(_0580_),
    .X(net20));
 sky130_fd_sc_hd__or2_1 _1504_ (.A(_0564_),
    .B(_0566_),
    .X(_0581_));
 sky130_fd_sc_hd__a21o_1 _1505_ (.A1(_0264_),
    .A2(_0328_),
    .B1(_0329_),
    .X(_0582_));
 sky130_fd_sc_hd__xor2_1 _1506_ (.A(_0570_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_1 _1507_ (.A(_0566_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__a21oi_1 _1508_ (.A1(_0581_),
    .A2(_0571_),
    .B1(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__and3_1 _1509_ (.A(_0581_),
    .B(_0571_),
    .C(_0584_),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _1510_ (.A(_0585_),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__nand2_1 _1511_ (.A(_0574_),
    .B(_0577_),
    .Y(_0588_));
 sky130_fd_sc_hd__xnor2_2 _1512_ (.A(_0587_),
    .B(_0588_),
    .Y(net21));
 sky130_fd_sc_hd__nor2_1 _1513_ (.A(_0198_),
    .B(_0560_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21bo_1 _1514_ (.A1(_0570_),
    .A2(_0582_),
    .B1_N(_0566_),
    .X(_0590_));
 sky130_fd_sc_hd__o21a_1 _1515_ (.A1(_0570_),
    .A2(_0582_),
    .B1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__and2_1 _1516_ (.A(_0589_),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _1517_ (.A1(_0581_),
    .A2(_0571_),
    .B1(_0584_),
    .X(_0593_));
 sky130_fd_sc_hd__a31o_1 _1518_ (.A1(_0574_),
    .A2(_0577_),
    .A3(_0593_),
    .B1(_0586_),
    .X(_0594_));
 sky130_fd_sc_hd__or2_1 _1519_ (.A(_0589_),
    .B(_0591_),
    .X(_0595_));
 sky130_fd_sc_hd__o21a_1 _1520_ (.A1(_0592_),
    .A2(_0594_),
    .B1(_0595_),
    .X(net22));
 sky130_fd_sc_hd__nor2_1 _1521_ (.A(_0314_),
    .B(_0315_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_2 _1522_ (.A(_0316_),
    .B(_0596_),
    .Y(net23));
 sky130_fd_sc_hd__clkbuf_4 _1523_ (.A(_0925_),
    .X(_0597_));
 sky130_fd_sc_hd__buf_4 _1524_ (.A(net32),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_4 _1525_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_4 _1526_ (.A(_0828_),
    .X(_0600_));
 sky130_fd_sc_hd__a21boi_2 _1527_ (.A1(_0599_),
    .A2(_0600_),
    .B1_N(_0817_),
    .Y(_0601_));
 sky130_fd_sc_hd__buf_4 _1528_ (.A(_0850_),
    .X(_0602_));
 sky130_fd_sc_hd__xnor2_4 _1529_ (.A(_0602_),
    .B(_0978_),
    .Y(_0603_));
 sky130_fd_sc_hd__clkbuf_4 _1530_ (.A(_0957_),
    .X(_0604_));
 sky130_fd_sc_hd__inv_2 _1531_ (.A(net35),
    .Y(_0605_));
 sky130_fd_sc_hd__buf_2 _1532_ (.A(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__or2b_1 _1533_ (.A(_0967_),
    .B_N(_0978_),
    .X(_0607_));
 sky130_fd_sc_hd__nand2b_2 _1534_ (.A_N(_0978_),
    .B(_0967_),
    .Y(_0608_));
 sky130_fd_sc_hd__clkbuf_4 _1535_ (.A(net36),
    .X(_0609_));
 sky130_fd_sc_hd__a41o_1 _1536_ (.A1(_0604_),
    .A2(_0606_),
    .A3(_0607_),
    .A4(_0608_),
    .B1(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__a21oi_1 _1537_ (.A1(_0601_),
    .A2(_0603_),
    .B1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__clkbuf_4 _1538_ (.A(_0817_),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_2 _1539_ (.A(_0602_),
    .B(net45),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_1 _1540_ (.A(_0612_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_2 _1541_ (.A(_0957_),
    .B(_0599_),
    .Y(_0615_));
 sky130_fd_sc_hd__clkbuf_4 _1542_ (.A(_0609_),
    .X(_0616_));
 sky130_fd_sc_hd__o31a_1 _1543_ (.A1(_0614_),
    .A2(_0615_),
    .A3(_0601_),
    .B1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2b_1 _1544_ (.A_N(_0967_),
    .B(_0957_),
    .Y(_0618_));
 sky130_fd_sc_hd__clkbuf_4 _1545_ (.A(_0817_),
    .X(_0619_));
 sky130_fd_sc_hd__and2b_1 _1546_ (.A_N(net45),
    .B(net33),
    .X(_0620_));
 sky130_fd_sc_hd__buf_2 _1547_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__and2b_2 _1548_ (.A_N(_0850_),
    .B(net45),
    .X(_0622_));
 sky130_fd_sc_hd__or3_1 _1549_ (.A(_0619_),
    .B(_0621_),
    .C(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__o21a_1 _1550_ (.A1(_0606_),
    .A2(_0618_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__inv_2 _1551_ (.A(_0925_),
    .Y(_0625_));
 sky130_fd_sc_hd__or3_4 _1552_ (.A(_0850_),
    .B(_0598_),
    .C(net45),
    .X(_0626_));
 sky130_fd_sc_hd__o21a_1 _1553_ (.A1(_0619_),
    .A2(_0626_),
    .B1(_0609_),
    .X(_0627_));
 sky130_fd_sc_hd__or2_1 _1554_ (.A(_0625_),
    .B(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__o32a_1 _1555_ (.A1(_0597_),
    .A2(_0611_),
    .A3(_0617_),
    .B1(_0624_),
    .B2(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__or2_1 _1556_ (.A(\p_shaping_I.p_shaping_I.counter[1] ),
    .B(\p_shaping_I.p_shaping_I.counter[0] ),
    .X(_0630_));
 sky130_fd_sc_hd__buf_2 _1557_ (.A(_0630_),
    .X(_0021_));
 sky130_fd_sc_hd__or2b_1 _1558_ (.A(_0629_),
    .B_N(_0021_),
    .X(_0631_));
 sky130_fd_sc_hd__xor2_4 _1559_ (.A(_0850_),
    .B(_0598_),
    .X(_0632_));
 sky130_fd_sc_hd__a21bo_1 _1560_ (.A1(_0602_),
    .A2(_0978_),
    .B1_N(_0828_),
    .X(_0633_));
 sky130_fd_sc_hd__o211a_1 _1561_ (.A1(_0600_),
    .A2(_0632_),
    .B1(_0633_),
    .C1(_0619_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2b_2 _1562_ (.A_N(_0957_),
    .B(_0967_),
    .Y(_0635_));
 sky130_fd_sc_hd__nor2_1 _1563_ (.A(_0612_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__o31a_1 _1564_ (.A1(_0616_),
    .A2(_0634_),
    .A3(_0636_),
    .B1(_0914_),
    .X(_0637_));
 sky130_fd_sc_hd__a21oi_4 _1565_ (.A1(_0957_),
    .A2(_0978_),
    .B1(_0967_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_2 _1566_ (.A(_0609_),
    .B(_0625_),
    .Y(_0639_));
 sky130_fd_sc_hd__o31a_1 _1567_ (.A1(_0606_),
    .A2(_0925_),
    .A3(_0638_),
    .B1(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a21bo_2 _1568_ (.A1(_0602_),
    .A2(_0598_),
    .B1_N(net35),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _1569_ (.A(_0602_),
    .B(_0828_),
    .X(_0642_));
 sky130_fd_sc_hd__and2b_1 _1570_ (.A_N(_0828_),
    .B(_0598_),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_2 _1571_ (.A(_0642_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2b_2 _1572_ (.A(_0598_),
    .B_N(_0602_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21a_1 _1573_ (.A1(_0600_),
    .A2(_0645_),
    .B1(_0606_),
    .X(_0646_));
 sky130_fd_sc_hd__a2bb2o_1 _1574_ (.A1_N(_0641_),
    .A2_N(_0644_),
    .B1(_0646_),
    .B2(_0608_),
    .X(_0647_));
 sky130_fd_sc_hd__o2bb2a_2 _1575_ (.A1_N(_0597_),
    .A2_N(_0637_),
    .B1(_0640_),
    .B2(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_4 _1576_ (.A(_0606_),
    .X(_0649_));
 sky130_fd_sc_hd__or2_2 _1577_ (.A(_0612_),
    .B(_0609_),
    .X(_0650_));
 sky130_fd_sc_hd__a21oi_1 _1578_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0609_),
    .Y(_0651_));
 sky130_fd_sc_hd__inv_2 _1579_ (.A(_0828_),
    .Y(_0652_));
 sky130_fd_sc_hd__a211o_1 _1580_ (.A1(_0817_),
    .A2(_0632_),
    .B1(_0925_),
    .C1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__clkinv_2 _1581_ (.A(_0609_),
    .Y(_0654_));
 sky130_fd_sc_hd__a211oi_4 _1582_ (.A1(_0850_),
    .A2(_0598_),
    .B1(net35),
    .C1(_0828_),
    .Y(_0655_));
 sky130_fd_sc_hd__or2_1 _1583_ (.A(_0654_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__and3_1 _1584_ (.A(_0978_),
    .B(_0817_),
    .C(_0613_),
    .X(_0657_));
 sky130_fd_sc_hd__o2bb2a_1 _1585_ (.A1_N(_0651_),
    .A2_N(_0653_),
    .B1(_0656_),
    .B2(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a221oi_4 _1586_ (.A1(_0649_),
    .A2(_0615_),
    .B1(_0650_),
    .B2(_0597_),
    .C1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _1587_ (.A(\p_shaping_I.p_shaping_I.counter[1] ),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__xor2_1 _1588_ (.A(_0648_),
    .B(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__xnor2_1 _1589_ (.A(_0631_),
    .B(_0661_),
    .Y(net6));
 sky130_fd_sc_hd__clkbuf_4 _1590_ (.A(\p_shaping_I.p_shaping_I.counter[1] ),
    .X(_0662_));
 sky130_fd_sc_hd__buf_2 _1591_ (.A(_0817_),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _1592_ (.A(_0605_),
    .B(_0600_),
    .C(_0632_),
    .X(_0664_));
 sky130_fd_sc_hd__or2_4 _1593_ (.A(_0609_),
    .B(_0925_),
    .X(_0665_));
 sky130_fd_sc_hd__a211o_1 _1594_ (.A1(_0663_),
    .A2(_0644_),
    .B1(_0664_),
    .C1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__buf_2 _1595_ (.A(_0967_),
    .X(_0667_));
 sky130_fd_sc_hd__nor2b_2 _1596_ (.A(_0602_),
    .B_N(_0598_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand3b_2 _1597_ (.A_N(_0957_),
    .B(_0817_),
    .C(_0600_),
    .Y(_0669_));
 sky130_fd_sc_hd__o32a_1 _1598_ (.A1(_0619_),
    .A2(_0667_),
    .A3(_0668_),
    .B1(_0669_),
    .B2(_0599_),
    .X(_0670_));
 sky130_fd_sc_hd__o21ai_1 _1599_ (.A1(_0627_),
    .A2(_0670_),
    .B1(_0925_),
    .Y(_0671_));
 sky130_fd_sc_hd__o311a_1 _1600_ (.A1(_0649_),
    .A2(_0639_),
    .A3(_0603_),
    .B1(_0666_),
    .C1(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _1601_ (.A(_0659_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_4 _1602_ (.A(_0616_),
    .B(_0925_),
    .Y(_0674_));
 sky130_fd_sc_hd__buf_2 _1603_ (.A(_0599_),
    .X(_0675_));
 sky130_fd_sc_hd__or2_1 _1604_ (.A(_0600_),
    .B(_0668_),
    .X(_0676_));
 sky130_fd_sc_hd__a32o_1 _1605_ (.A1(_0675_),
    .A2(_0667_),
    .A3(_0641_),
    .B1(_0676_),
    .B2(_0601_),
    .X(_0677_));
 sky130_fd_sc_hd__and2_1 _1606_ (.A(_0599_),
    .B(_0621_),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _1607_ (.A(_0602_),
    .B(_0978_),
    .C(_0828_),
    .X(_0679_));
 sky130_fd_sc_hd__o32a_1 _1608_ (.A1(_0619_),
    .A2(_0600_),
    .A3(_0668_),
    .B1(_0638_),
    .B2(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__a211oi_1 _1609_ (.A1(_0606_),
    .A2(_0678_),
    .B1(_0680_),
    .C1(_0639_),
    .Y(_0681_));
 sky130_fd_sc_hd__nor2_1 _1610_ (.A(_0609_),
    .B(_0625_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _1611_ (.A(_0978_),
    .B(_0967_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1612_ (.A(_0612_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__and3b_1 _1613_ (.A_N(_0646_),
    .B(_0682_),
    .C(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__a211oi_2 _1614_ (.A1(_0674_),
    .A2(_0677_),
    .B1(_0681_),
    .C1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__o21ai_1 _1615_ (.A1(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .A2(_0673_),
    .B1(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__or3_1 _1616_ (.A(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .B(_0673_),
    .C(_0686_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _1617_ (.A(_0604_),
    .B(_0683_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2b_2 _1618_ (.A_N(_0967_),
    .B(_0817_),
    .Y(_0690_));
 sky130_fd_sc_hd__o311a_1 _1619_ (.A1(_0663_),
    .A2(_0678_),
    .A3(_0689_),
    .B1(_0690_),
    .C1(_0641_),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_2 _1620_ (.A(_0612_),
    .B(_0608_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _1621_ (.A(_0652_),
    .B(_0603_),
    .Y(_0693_));
 sky130_fd_sc_hd__clkbuf_4 _1622_ (.A(_0903_),
    .X(_0694_));
 sky130_fd_sc_hd__o211a_1 _1623_ (.A1(_0622_),
    .A2(_0692_),
    .B1(_0693_),
    .C1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__nor2_2 _1624_ (.A(_0599_),
    .B(_0619_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _1625_ (.A(_0663_),
    .B(_0618_),
    .Y(_0697_));
 sky130_fd_sc_hd__o31a_1 _1626_ (.A1(_0696_),
    .A2(_0657_),
    .A3(_0697_),
    .B1(_0682_),
    .X(_0698_));
 sky130_fd_sc_hd__a211o_1 _1627_ (.A1(_0674_),
    .A2(_0691_),
    .B1(_0695_),
    .C1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__inv_2 _1628_ (.A(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__a211o_1 _1629_ (.A1(_0663_),
    .A2(_0644_),
    .B1(_0655_),
    .C1(_0664_),
    .X(_0701_));
 sky130_fd_sc_hd__o211a_1 _1630_ (.A1(_0663_),
    .A2(_0645_),
    .B1(_0641_),
    .C1(_0690_),
    .X(_0702_));
 sky130_fd_sc_hd__o21ba_1 _1631_ (.A1(_0978_),
    .A2(_0967_),
    .B1_N(_0602_),
    .X(_0703_));
 sky130_fd_sc_hd__nor2_1 _1632_ (.A(_0612_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__o21a_1 _1633_ (.A1(_0892_),
    .A2(_0704_),
    .B1(_0694_),
    .X(_0705_));
 sky130_fd_sc_hd__a221oi_4 _1634_ (.A1(_0682_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0674_),
    .C1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__a21oi_1 _1635_ (.A1(_0648_),
    .A2(_0706_),
    .B1(_0127_),
    .Y(_0707_));
 sky130_fd_sc_hd__xnor2_1 _1636_ (.A(_0700_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__and4_1 _1637_ (.A(_0662_),
    .B(_0687_),
    .C(_0688_),
    .D(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__a31oi_2 _1638_ (.A1(_0662_),
    .A2(_0687_),
    .A3(_0688_),
    .B1(_0708_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _1639_ (.A(_0616_),
    .B(_0989_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _1640_ (.A(_0663_),
    .B(_0703_),
    .Y(_0712_));
 sky130_fd_sc_hd__nand3b_1 _1641_ (.A_N(_0664_),
    .B(_0711_),
    .C(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21o_1 _1642_ (.A1(_0957_),
    .A2(_0600_),
    .B1(_0619_),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _1643_ (.A(_0616_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__nor2_1 _1644_ (.A(_0606_),
    .B(_0613_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor4_1 _1645_ (.A(_0675_),
    .B(_0925_),
    .C(_0715_),
    .D(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__a211o_1 _1646_ (.A1(_0667_),
    .A2(_0603_),
    .B1(_0643_),
    .C1(_0612_),
    .X(_0718_));
 sky130_fd_sc_hd__a21oi_1 _1647_ (.A1(_0712_),
    .A2(_0718_),
    .B1(_0665_),
    .Y(_0719_));
 sky130_fd_sc_hd__a211o_2 _1648_ (.A1(_0597_),
    .A2(_0713_),
    .B1(_0717_),
    .C1(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(_0667_),
    .B(_0632_),
    .Y(_0721_));
 sky130_fd_sc_hd__o21ai_2 _1650_ (.A1(_0957_),
    .A2(_0599_),
    .B1(_0667_),
    .Y(_0722_));
 sky130_fd_sc_hd__a21oi_1 _1651_ (.A1(_0604_),
    .A2(_0606_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o311a_1 _1652_ (.A1(_0616_),
    .A2(_0721_),
    .A3(_0723_),
    .B1(_0925_),
    .C1(_0914_),
    .X(_0724_));
 sky130_fd_sc_hd__a31oi_1 _1653_ (.A1(_0696_),
    .A2(_0618_),
    .A3(_0635_),
    .B1(_0616_),
    .Y(_0725_));
 sky130_fd_sc_hd__o21ai_1 _1654_ (.A1(_0675_),
    .A2(_0618_),
    .B1(_0601_),
    .Y(_0726_));
 sky130_fd_sc_hd__o2111a_1 _1655_ (.A1(_0612_),
    .A2(_0621_),
    .B1(_0641_),
    .C1(_0690_),
    .D1(_0694_),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_1 _1656_ (.A1(_0625_),
    .A2(_0725_),
    .A3(_0726_),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1657_ (.A(_0724_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__a21oi_1 _1658_ (.A1(_0629_),
    .A2(_0729_),
    .B1(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .Y(_0730_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(_0720_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__a21oi_2 _1660_ (.A1(\p_shaping_I.p_shaping_I.ctl_1 ),
    .A2(net49),
    .B1(_0127_),
    .Y(_0732_));
 sky130_fd_sc_hd__and3_1 _1661_ (.A(\p_shaping_I.p_shaping_I.ctl_1 ),
    .B(net49),
    .C(_0127_),
    .X(_0733_));
 sky130_fd_sc_hd__nor3_4 _1662_ (.A(_0042_),
    .B(_0732_),
    .C(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21o_1 _1663_ (.A1(_0720_),
    .A2(_0730_),
    .B1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_4 _1664_ (.A(_0612_),
    .X(_0736_));
 sky130_fd_sc_hd__a21oi_1 _1665_ (.A1(_0604_),
    .A2(_0667_),
    .B1(_0599_),
    .Y(_0737_));
 sky130_fd_sc_hd__a21oi_2 _1666_ (.A1(_0736_),
    .A2(_0737_),
    .B1(_0655_),
    .Y(_0738_));
 sky130_fd_sc_hd__a211o_1 _1667_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0645_),
    .C1(_0663_),
    .X(_0739_));
 sky130_fd_sc_hd__a21oi_1 _1668_ (.A1(_0692_),
    .A2(_0739_),
    .B1(_0738_),
    .Y(_0740_));
 sky130_fd_sc_hd__or2_1 _1669_ (.A(_0675_),
    .B(_0690_),
    .X(_0741_));
 sky130_fd_sc_hd__a21o_1 _1670_ (.A1(_0725_),
    .A2(_0741_),
    .B1(_0625_),
    .X(_0742_));
 sky130_fd_sc_hd__o221ai_4 _1671_ (.A1(_0665_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(_0639_),
    .C1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__a311o_1 _1672_ (.A1(_0736_),
    .A2(_0693_),
    .A3(_0722_),
    .B1(_0636_),
    .C1(_0627_),
    .X(_0744_));
 sky130_fd_sc_hd__nor2_1 _1673_ (.A(_0652_),
    .B(_0603_),
    .Y(_0745_));
 sky130_fd_sc_hd__nor2_2 _1674_ (.A(_0602_),
    .B(_0828_),
    .Y(_0746_));
 sky130_fd_sc_hd__o221a_1 _1675_ (.A1(_0736_),
    .A2(_0635_),
    .B1(_0745_),
    .B2(_0746_),
    .C1(_0674_),
    .X(_0747_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_0663_),
    .B(_0683_),
    .Y(_0748_));
 sky130_fd_sc_hd__o21a_1 _1677_ (.A1(_0657_),
    .A2(_0748_),
    .B1(_0694_),
    .X(_0749_));
 sky130_fd_sc_hd__a211o_1 _1678_ (.A1(_0597_),
    .A2(_0744_),
    .B1(_0747_),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__a31o_2 _1679_ (.A1(_0720_),
    .A2(_0743_),
    .A3(_0750_),
    .B1(_0129_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _1680_ (.A(_0734_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__o211a_1 _1681_ (.A1(_0731_),
    .A2(_0735_),
    .B1(_0752_),
    .C1(_0021_),
    .X(_0753_));
 sky130_fd_sc_hd__o21bai_1 _1682_ (.A1(_0709_),
    .A2(_0710_),
    .B1_N(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__or3b_1 _1683_ (.A(_0709_),
    .B(_0710_),
    .C_N(_0753_),
    .X(_0755_));
 sky130_fd_sc_hd__clkinv_2 _1684_ (.A(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .Y(_0756_));
 sky130_fd_sc_hd__a21oi_1 _1685_ (.A1(_0756_),
    .A2(_0659_),
    .B1(_0672_),
    .Y(_0757_));
 sky130_fd_sc_hd__inv_2 _1686_ (.A(\p_shaping_I.p_shaping_I.counter[1] ),
    .Y(_0758_));
 sky130_fd_sc_hd__a31o_1 _1687_ (.A1(_0756_),
    .A2(_0659_),
    .A3(_0672_),
    .B1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__or2_1 _1688_ (.A(_0757_),
    .B(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__or2_1 _1689_ (.A(_0127_),
    .B(_0648_),
    .X(_0761_));
 sky130_fd_sc_hd__xnor2_1 _1690_ (.A(_0706_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _1691_ (.A(_0760_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ai_1 _1692_ (.A1(_0129_),
    .A2(_0629_),
    .B1(_0729_),
    .Y(_0764_));
 sky130_fd_sc_hd__or3_1 _1693_ (.A(_0129_),
    .B(_0629_),
    .C(_0729_),
    .X(_0765_));
 sky130_fd_sc_hd__and3_1 _1694_ (.A(_0021_),
    .B(_0764_),
    .C(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1695_ (.A(_0760_),
    .B(_0762_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21o_1 _1696_ (.A1(_0763_),
    .A2(_0766_),
    .B1(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__and3_1 _1697_ (.A(_0754_),
    .B(_0755_),
    .C(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__a21o_1 _1698_ (.A1(_0754_),
    .A2(_0755_),
    .B1(_0768_),
    .X(_0770_));
 sky130_fd_sc_hd__and2b_1 _1699_ (.A_N(_0769_),
    .B(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__and2b_1 _1700_ (.A_N(_0631_),
    .B(_0661_),
    .X(_0772_));
 sky130_fd_sc_hd__o21ba_1 _1701_ (.A1(_0648_),
    .A2(_0660_),
    .B1_N(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__xnor2_1 _1702_ (.A(_0760_),
    .B(_0762_),
    .Y(_0774_));
 sky130_fd_sc_hd__xnor2_2 _1703_ (.A(_0774_),
    .B(_0766_),
    .Y(_0775_));
 sky130_fd_sc_hd__and2b_1 _1704_ (.A_N(_0773_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__xor2_1 _1705_ (.A(_0771_),
    .B(_0776_),
    .X(net11));
 sky130_fd_sc_hd__nor3b_1 _1706_ (.A(_0709_),
    .B(_0710_),
    .C_N(_0753_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor3b_1 _1707_ (.A(_0659_),
    .B(_0672_),
    .C_N(_0686_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21o_1 _1708_ (.A1(_0600_),
    .A2(_0632_),
    .B1(_0643_),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _1709_ (.A(_0704_),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__nor2_1 _1710_ (.A(_0704_),
    .B(_0779_),
    .Y(_0781_));
 sky130_fd_sc_hd__and2b_1 _1711_ (.A_N(_0598_),
    .B(_0828_),
    .X(_0782_));
 sky130_fd_sc_hd__o31a_1 _1712_ (.A1(_0619_),
    .A2(_0746_),
    .A3(_0782_),
    .B1(_0609_),
    .X(_0783_));
 sky130_fd_sc_hd__or3_1 _1713_ (.A(_0621_),
    .B(_0622_),
    .C(_0641_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(_0598_),
    .A1(_0850_),
    .S(net45),
    .X(_0785_));
 sky130_fd_sc_hd__o21ai_1 _1715_ (.A1(_0612_),
    .A2(_0785_),
    .B1(_0654_),
    .Y(_0786_));
 sky130_fd_sc_hd__o2111a_1 _1716_ (.A1(_0600_),
    .A2(_0632_),
    .B1(_0633_),
    .C1(_0785_),
    .D1(_0619_),
    .X(_0787_));
 sky130_fd_sc_hd__o2bb2a_1 _1717_ (.A1_N(_0783_),
    .A2_N(_0784_),
    .B1(_0786_),
    .B2(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__o32a_1 _1718_ (.A1(_0871_),
    .A2(_0780_),
    .A3(_0781_),
    .B1(_0788_),
    .B2(_0597_),
    .X(_0789_));
 sky130_fd_sc_hd__o21ai_1 _1719_ (.A1(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .A2(_0778_),
    .B1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__or3_1 _1720_ (.A(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .B(_0789_),
    .C(_0778_),
    .X(_0791_));
 sky130_fd_sc_hd__and3_1 _1721_ (.A(\p_shaping_I.p_shaping_I.counter[1] ),
    .B(_0790_),
    .C(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__a31o_1 _1722_ (.A1(_0648_),
    .A2(_0700_),
    .A3(_0706_),
    .B1(_0127_),
    .X(_0793_));
 sky130_fd_sc_hd__nor4_1 _1723_ (.A(_0663_),
    .B(_0667_),
    .C(_0668_),
    .D(_0645_),
    .Y(_0794_));
 sky130_fd_sc_hd__nor2_1 _1724_ (.A(_0641_),
    .B(_0737_),
    .Y(_0795_));
 sky130_fd_sc_hd__o311a_1 _1725_ (.A1(_0616_),
    .A2(_0794_),
    .A3(_0795_),
    .B1(_0597_),
    .C1(_0989_),
    .X(_0796_));
 sky130_fd_sc_hd__nor2_1 _1726_ (.A(_0606_),
    .B(_0782_),
    .Y(_0797_));
 sky130_fd_sc_hd__or2_1 _1727_ (.A(_0599_),
    .B(_0669_),
    .X(_0798_));
 sky130_fd_sc_hd__o2111a_1 _1728_ (.A1(_0615_),
    .A2(_0797_),
    .B1(_0798_),
    .C1(_0626_),
    .D1(_0694_),
    .X(_0799_));
 sky130_fd_sc_hd__nor2_1 _1729_ (.A(_0663_),
    .B(_0645_),
    .Y(_0800_));
 sky130_fd_sc_hd__a211o_1 _1730_ (.A1(_0667_),
    .A2(_0800_),
    .B1(_0657_),
    .C1(_0665_),
    .X(_0801_));
 sky130_fd_sc_hd__or3b_2 _1731_ (.A(_0796_),
    .B(_0799_),
    .C_N(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__xor2_1 _1732_ (.A(_0793_),
    .B(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__xnor2_1 _1733_ (.A(_0792_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__or3_1 _1734_ (.A(_0042_),
    .B(_0732_),
    .C(_0733_),
    .X(_0805_));
 sky130_fd_sc_hd__a31o_1 _1735_ (.A1(_0629_),
    .A2(_0720_),
    .A3(_0729_),
    .B1(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .X(_0806_));
 sky130_fd_sc_hd__xnor2_1 _1736_ (.A(_0750_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__o21a_2 _1737_ (.A1(_0805_),
    .A2(_0807_),
    .B1(_0021_),
    .X(_0808_));
 sky130_fd_sc_hd__a21bo_1 _1738_ (.A1(_0805_),
    .A2(_0807_),
    .B1_N(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__xor2_1 _1739_ (.A(_0804_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__o21a_1 _1740_ (.A1(_0709_),
    .A2(_0777_),
    .B1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__or3_1 _1741_ (.A(_0709_),
    .B(_0777_),
    .C(_0810_),
    .X(_0812_));
 sky130_fd_sc_hd__and2b_1 _1742_ (.A_N(_0811_),
    .B(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__a21o_1 _1743_ (.A1(_0770_),
    .A2(_0776_),
    .B1(_0769_),
    .X(_0814_));
 sky130_fd_sc_hd__xor2_1 _1744_ (.A(_0813_),
    .B(_0814_),
    .X(net12));
 sky130_fd_sc_hd__and2_1 _1745_ (.A(_0792_),
    .B(_0803_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _1746_ (.A(_0804_),
    .B(_0809_),
    .Y(_0816_));
 sky130_fd_sc_hd__or4bb_1 _1747_ (.A(_0659_),
    .B(_0672_),
    .C_N(_0686_),
    .D_N(_0789_),
    .X(_0818_));
 sky130_fd_sc_hd__or2_1 _1748_ (.A(_0957_),
    .B(_0599_),
    .X(_0819_));
 sky130_fd_sc_hd__nand2_1 _1749_ (.A(_0675_),
    .B(_0621_),
    .Y(_0820_));
 sky130_fd_sc_hd__a31o_1 _1750_ (.A1(_0736_),
    .A2(_0819_),
    .A3(_0820_),
    .B1(_0871_),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _1751_ (.A(_0675_),
    .B(_0613_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21bo_1 _1752_ (.A1(_0892_),
    .A2(_0822_),
    .B1_N(_0718_),
    .X(_0823_));
 sky130_fd_sc_hd__a2bb2o_1 _1753_ (.A1_N(_0664_),
    .A2_N(_0821_),
    .B1(_0823_),
    .B2(_0694_),
    .X(_0824_));
 sky130_fd_sc_hd__a31o_1 _1754_ (.A1(_0714_),
    .A2(_0674_),
    .A3(_0641_),
    .B1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__a21oi_1 _1755_ (.A1(_0756_),
    .A2(_0818_),
    .B1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a31o_1 _1756_ (.A1(_0756_),
    .A2(_0818_),
    .A3(_0825_),
    .B1(_0758_),
    .X(_0827_));
 sky130_fd_sc_hd__or2_1 _1757_ (.A(_0826_),
    .B(_0827_),
    .X(_0829_));
 sky130_fd_sc_hd__nand4b_2 _1758_ (.A_N(_0699_),
    .B(_0802_),
    .C(_0706_),
    .D(_0648_),
    .Y(_0830_));
 sky130_fd_sc_hd__and2b_1 _1759_ (.A_N(\p_shaping_I.p_shaping_I.bit_in ),
    .B(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and3_1 _1760_ (.A(_0736_),
    .B(_0635_),
    .C(_0626_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_2 _1761_ (.A(_0616_),
    .X(_0833_));
 sky130_fd_sc_hd__o21ai_1 _1762_ (.A1(_0748_),
    .A2(_0832_),
    .B1(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__buf_2 _1763_ (.A(_0625_),
    .X(_0835_));
 sky130_fd_sc_hd__a31o_1 _1764_ (.A1(_0604_),
    .A2(_0835_),
    .A3(_0714_),
    .B1(_0694_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _1765_ (.A(_0606_),
    .B(_0608_),
    .Y(_0837_));
 sky130_fd_sc_hd__o211a_1 _1766_ (.A1(_0668_),
    .A2(_0837_),
    .B1(_0798_),
    .C1(_0820_),
    .X(_0838_));
 sky130_fd_sc_hd__o2bb2a_1 _1767_ (.A1_N(_0834_),
    .A2_N(_0836_),
    .B1(_0838_),
    .B2(_0871_),
    .X(_0840_));
 sky130_fd_sc_hd__xnor2_1 _1768_ (.A(_0831_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__xnor2_1 _1769_ (.A(_0829_),
    .B(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a21oi_1 _1770_ (.A1(_0720_),
    .A2(_0750_),
    .B1(_0129_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _1771_ (.A(_0730_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__buf_2 _1772_ (.A(_0597_),
    .X(_0845_));
 sky130_fd_sc_hd__or2_1 _1773_ (.A(_0604_),
    .B(_0608_),
    .X(_0846_));
 sky130_fd_sc_hd__or4b_1 _1774_ (.A(_0833_),
    .B(_0621_),
    .C(_0634_),
    .D_N(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__or2b_1 _1775_ (.A(_0627_),
    .B_N(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__or2b_1 _1776_ (.A(_0604_),
    .B_N(_0690_),
    .X(_0849_));
 sky130_fd_sc_hd__a21oi_1 _1777_ (.A1(_0696_),
    .A2(_0621_),
    .B1(_0668_),
    .Y(_0851_));
 sky130_fd_sc_hd__a221o_1 _1778_ (.A1(_0651_),
    .A2(_0849_),
    .B1(_0851_),
    .B2(_0833_),
    .C1(_0845_),
    .X(_0852_));
 sky130_fd_sc_hd__a21boi_1 _1779_ (.A1(_0845_),
    .A2(_0848_),
    .B1_N(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__nor2_1 _1780_ (.A(_0844_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__a21o_1 _1781_ (.A1(_0844_),
    .A2(_0853_),
    .B1(_0734_),
    .X(_0855_));
 sky130_fd_sc_hd__o21a_1 _1782_ (.A1(_0854_),
    .A2(_0855_),
    .B1(_0808_),
    .X(_0856_));
 sky130_fd_sc_hd__xor2_1 _1783_ (.A(_0842_),
    .B(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__o21a_1 _1784_ (.A1(_0815_),
    .A2(_0816_),
    .B1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__or3_1 _1785_ (.A(_0815_),
    .B(_0816_),
    .C(_0857_),
    .X(_0859_));
 sky130_fd_sc_hd__or2b_2 _1786_ (.A(_0858_),
    .B_N(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a21o_2 _1787_ (.A1(_0812_),
    .A2(_0814_),
    .B1(_0811_),
    .X(_0862_));
 sky130_fd_sc_hd__xnor2_4 _1788_ (.A(_0860_),
    .B(_0862_),
    .Y(net13));
 sky130_fd_sc_hd__and2b_1 _1789_ (.A_N(_0829_),
    .B(_0841_),
    .X(_0863_));
 sky130_fd_sc_hd__and2_1 _1790_ (.A(_0842_),
    .B(_0856_),
    .X(_0864_));
 sky130_fd_sc_hd__nor2_1 _1791_ (.A(_0818_),
    .B(_0825_),
    .Y(_0865_));
 sky130_fd_sc_hd__o21ai_1 _1792_ (.A1(_0649_),
    .A2(_0638_),
    .B1(_0861_),
    .Y(_0866_));
 sky130_fd_sc_hd__o32a_1 _1793_ (.A1(_0642_),
    .A2(_0746_),
    .A3(_0837_),
    .B1(_0632_),
    .B2(_0684_),
    .X(_0867_));
 sky130_fd_sc_hd__o2bb2a_1 _1794_ (.A1_N(_0616_),
    .A2_N(_0867_),
    .B1(_0797_),
    .B2(_0610_),
    .X(_0868_));
 sky130_fd_sc_hd__a2bb2o_1 _1795_ (.A1_N(_0871_),
    .A2_N(_0866_),
    .B1(_0868_),
    .B2(_0835_),
    .X(_0869_));
 sky130_fd_sc_hd__inv_2 _1796_ (.A(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__o21a_1 _1797_ (.A1(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .A2(_0865_),
    .B1(_0870_),
    .X(_0872_));
 sky130_fd_sc_hd__or3_1 _1798_ (.A(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .B(_0870_),
    .C(_0865_),
    .X(_0873_));
 sky130_fd_sc_hd__or3b_1 _1799_ (.A(_0872_),
    .B(_0758_),
    .C_N(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__and2b_1 _1800_ (.A_N(_0830_),
    .B(_0840_),
    .X(_0875_));
 sky130_fd_sc_hd__nor2_1 _1801_ (.A(\p_shaping_I.p_shaping_I.bit_in ),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand3_1 _1802_ (.A(_0714_),
    .B(_0694_),
    .C(_0726_),
    .Y(_0877_));
 sky130_fd_sc_hd__or3b_1 _1803_ (.A(_0736_),
    .B(_0746_),
    .C_N(_0675_),
    .X(_0878_));
 sky130_fd_sc_hd__a31o_1 _1804_ (.A1(_0690_),
    .A2(_0626_),
    .A3(_0878_),
    .B1(_0628_),
    .X(_0879_));
 sky130_fd_sc_hd__o211a_1 _1805_ (.A1(_0690_),
    .A2(_0665_),
    .B1(_0877_),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__xnor2_1 _1806_ (.A(_0876_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__xor2_1 _1807_ (.A(_0874_),
    .B(_0881_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(_0129_),
    .A1(_0843_),
    .S(_0743_),
    .X(_0884_));
 sky130_fd_sc_hd__o21ai_1 _1809_ (.A1(_0734_),
    .A2(_0884_),
    .B1(_0808_),
    .Y(_0885_));
 sky130_fd_sc_hd__xor2_1 _1810_ (.A(_0883_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__nor3_1 _1811_ (.A(_0863_),
    .B(_0864_),
    .C(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__o21a_1 _1812_ (.A1(_0863_),
    .A2(_0864_),
    .B1(_0886_),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_1 _1813_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__a21oi_1 _1814_ (.A1(_0859_),
    .A2(_0862_),
    .B1(_0858_),
    .Y(_0890_));
 sky130_fd_sc_hd__xnor2_2 _1815_ (.A(_0889_),
    .B(_0890_),
    .Y(net14));
 sky130_fd_sc_hd__and2b_1 _1816_ (.A_N(_0874_),
    .B(_0881_),
    .X(_0891_));
 sky130_fd_sc_hd__nor2_1 _1817_ (.A(_0883_),
    .B(_0885_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_1 _1818_ (.A(_0667_),
    .B(_0819_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _1819_ (.A(_0833_),
    .B(_0722_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_1 _1820_ (.A(_0894_),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__a21oi_1 _1821_ (.A1(_0649_),
    .A2(_0746_),
    .B1(_0696_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_1 _1822_ (.A1(_0833_),
    .A2(_0669_),
    .B1(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__a41o_1 _1823_ (.A1(_0833_),
    .A2(_0626_),
    .A3(_0722_),
    .A4(_0897_),
    .B1(_0597_),
    .X(_0899_));
 sky130_fd_sc_hd__a21oi_1 _1824_ (.A1(_0896_),
    .A2(_0898_),
    .B1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__o21ba_1 _1825_ (.A1(_0871_),
    .A2(_0861_),
    .B1_N(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__o31a_2 _1826_ (.A1(_0818_),
    .A2(_0825_),
    .A3(_0869_),
    .B1(_0756_),
    .X(_0902_));
 sky130_fd_sc_hd__xnor2_1 _1827_ (.A(_0901_),
    .B(_0902_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _1828_ (.A(_0662_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21oi_2 _1829_ (.A1(_0875_),
    .A2(_0880_),
    .B1(\p_shaping_I.p_shaping_I.bit_in ),
    .Y(_0906_));
 sky130_fd_sc_hd__o21a_1 _1830_ (.A1(_0652_),
    .A2(_0632_),
    .B1(_0892_),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _1831_ (.A(_0715_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__and2_1 _1832_ (.A(_0654_),
    .B(_0839_),
    .X(_0909_));
 sky130_fd_sc_hd__a21o_1 _1833_ (.A1(_0692_),
    .A2(_0739_),
    .B1(_0871_),
    .X(_0910_));
 sky130_fd_sc_hd__o31a_1 _1834_ (.A1(_0845_),
    .A2(_0908_),
    .A3(_0909_),
    .B1(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(\p_shaping_I.p_shaping_I.bit_in ),
    .A1(_0906_),
    .S(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__xor2_1 _1836_ (.A(_0905_),
    .B(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__o31a_1 _1837_ (.A1(_0649_),
    .A2(_0679_),
    .A3(_0621_),
    .B1(_0822_),
    .X(_0915_));
 sky130_fd_sc_hd__a31o_1 _1838_ (.A1(_0675_),
    .A2(_0613_),
    .A3(_0892_),
    .B1(_0871_),
    .X(_0916_));
 sky130_fd_sc_hd__nor2_1 _1839_ (.A(_0833_),
    .B(_0721_),
    .Y(_0917_));
 sky130_fd_sc_hd__o21ai_1 _1840_ (.A1(_0736_),
    .A2(_0608_),
    .B1(_0676_),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_1 _1841_ (.A(_0895_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__and3_1 _1842_ (.A(_0649_),
    .B(_0782_),
    .C(_0895_),
    .X(_0920_));
 sky130_fd_sc_hd__a211o_1 _1843_ (.A1(_0797_),
    .A2(_0917_),
    .B1(_0919_),
    .C1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a2bb2o_1 _1844_ (.A1_N(_0915_),
    .A2_N(_0916_),
    .B1(_0921_),
    .B2(_0835_),
    .X(_0922_));
 sky130_fd_sc_hd__xnor2_1 _1845_ (.A(_0751_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__o21ai_1 _1846_ (.A1(_0734_),
    .A2(_0923_),
    .B1(_0808_),
    .Y(_0924_));
 sky130_fd_sc_hd__xor2_1 _1847_ (.A(_0913_),
    .B(_0924_),
    .X(_0926_));
 sky130_fd_sc_hd__o21a_1 _1848_ (.A1(_0891_),
    .A2(_0893_),
    .B1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nor3_1 _1849_ (.A(_0891_),
    .B(_0893_),
    .C(_0926_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_2 _1850_ (.A(_0927_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(_0887_),
    .Y(_0930_));
 sky130_fd_sc_hd__a211o_1 _1852_ (.A1(_0859_),
    .A2(_0862_),
    .B1(_0888_),
    .C1(_0858_),
    .X(_0931_));
 sky130_fd_sc_hd__nand2_2 _1853_ (.A(_0930_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__xnor2_4 _1854_ (.A(_0929_),
    .B(_0932_),
    .Y(net15));
 sky130_fd_sc_hd__and3_1 _1855_ (.A(_0662_),
    .B(_0904_),
    .C(_0912_),
    .X(_0933_));
 sky130_fd_sc_hd__nor2_1 _1856_ (.A(_0913_),
    .B(_0924_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _1857_ (.A(_0718_),
    .B(_0909_),
    .Y(_0936_));
 sky130_fd_sc_hd__nor2_1 _1858_ (.A(_0649_),
    .B(_0894_),
    .Y(_0937_));
 sky130_fd_sc_hd__or4_1 _1859_ (.A(_0654_),
    .B(_0622_),
    .C(_0678_),
    .D(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__a21o_1 _1860_ (.A1(_0936_),
    .A2(_0938_),
    .B1(_0845_),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_2 _1861_ (.A(_0902_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _1862_ (.A(_0662_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__or3_1 _1863_ (.A(_0736_),
    .B(_0679_),
    .C(_0638_),
    .X(_0942_));
 sky130_fd_sc_hd__and3_1 _1864_ (.A(_0892_),
    .B(_0694_),
    .C(_0722_),
    .X(_0943_));
 sky130_fd_sc_hd__a41o_1 _1865_ (.A1(_0845_),
    .A2(_0669_),
    .A3(_0711_),
    .A4(_0942_),
    .B1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__xor2_2 _1866_ (.A(_0906_),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_1 _1867_ (.A(_0941_),
    .B(_0945_),
    .X(_0947_));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(_0745_),
    .Y(_0948_));
 sky130_fd_sc_hd__and3_1 _1869_ (.A(_0649_),
    .B(_0693_),
    .C(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__a21oi_1 _1870_ (.A1(_0635_),
    .A2(_0601_),
    .B1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a22o_1 _1871_ (.A1(_0649_),
    .A2(_0644_),
    .B1(_0948_),
    .B2(_0937_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _1872_ (.A0(_0950_),
    .A1(_0951_),
    .S(_0654_),
    .X(_0952_));
 sky130_fd_sc_hd__xnor2_1 _1873_ (.A(_0604_),
    .B(_0692_),
    .Y(_0953_));
 sky130_fd_sc_hd__o211a_1 _1874_ (.A1(_0833_),
    .A2(_0953_),
    .B1(_0989_),
    .C1(_0845_),
    .X(_0954_));
 sky130_fd_sc_hd__a211o_1 _1875_ (.A1(_0835_),
    .A2(_0952_),
    .B1(_0954_),
    .C1(_0734_),
    .X(_0955_));
 sky130_fd_sc_hd__nand2_1 _1876_ (.A(_0751_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__o211a_1 _1877_ (.A1(_0129_),
    .A2(_0955_),
    .B1(_0956_),
    .C1(_0021_),
    .X(_0958_));
 sky130_fd_sc_hd__xnor2_1 _1878_ (.A(_0947_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__o21a_1 _1879_ (.A1(_0933_),
    .A2(_0934_),
    .B1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__nor3_1 _1880_ (.A(_0933_),
    .B(_0934_),
    .C(_0959_),
    .Y(_0961_));
 sky130_fd_sc_hd__nor2_1 _1881_ (.A(_0960_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a31o_1 _1882_ (.A1(_0930_),
    .A2(_0929_),
    .A3(_0931_),
    .B1(_0927_),
    .X(_0963_));
 sky130_fd_sc_hd__xor2_2 _1883_ (.A(_0962_),
    .B(_0963_),
    .X(net16));
 sky130_fd_sc_hd__a22o_1 _1884_ (.A1(_0604_),
    .A2(_0797_),
    .B1(_0820_),
    .B2(_0649_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _1885_ (.A1(_0846_),
    .A2(_0964_),
    .B1(_0833_),
    .Y(_0965_));
 sky130_fd_sc_hd__and3b_1 _1886_ (.A_N(_0965_),
    .B(_0880_),
    .C(_0875_),
    .X(_0966_));
 sky130_fd_sc_hd__nor2_1 _1887_ (.A(\p_shaping_I.p_shaping_I.bit_in ),
    .B(_0966_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux2_1 _1888_ (.A0(\p_shaping_I.p_shaping_I.bit_in ),
    .A1(_0968_),
    .S(_0946_),
    .X(_0969_));
 sky130_fd_sc_hd__o311a_1 _1889_ (.A1(_0622_),
    .A2(_0721_),
    .A3(_0837_),
    .B1(_0690_),
    .C1(_0654_),
    .X(_0970_));
 sky130_fd_sc_hd__o31a_1 _1890_ (.A1(_0597_),
    .A2(_0655_),
    .A3(_0937_),
    .B1(_0665_),
    .X(_0971_));
 sky130_fd_sc_hd__or2_1 _1891_ (.A(_0970_),
    .B(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__o21ai_1 _1892_ (.A1(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .A2(_0848_),
    .B1(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__or2_1 _1893_ (.A(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .B(_0972_),
    .X(_0974_));
 sky130_fd_sc_hd__o211a_1 _1894_ (.A1(_0902_),
    .A2(_0973_),
    .B1(_0974_),
    .C1(_0662_),
    .X(_0975_));
 sky130_fd_sc_hd__xor2_2 _1895_ (.A(_0969_),
    .B(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__o21ai_1 _1896_ (.A1(_0627_),
    .A2(_0949_),
    .B1(_0845_),
    .Y(_0977_));
 sky130_fd_sc_hd__a21oi_1 _1897_ (.A1(_0683_),
    .A2(_0800_),
    .B1(_0716_),
    .Y(_0979_));
 sky130_fd_sc_hd__or3_1 _1898_ (.A(_0694_),
    .B(_0684_),
    .C(_0737_),
    .X(_0980_));
 sky130_fd_sc_hd__or4_1 _1899_ (.A(_0845_),
    .B(_0621_),
    .C(_0650_),
    .D(_0745_),
    .X(_0981_));
 sky130_fd_sc_hd__o211a_1 _1900_ (.A1(_0639_),
    .A2(_0979_),
    .B1(_0980_),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a21oi_1 _1901_ (.A1(_0977_),
    .A2(_0982_),
    .B1(_0751_),
    .Y(_0983_));
 sky130_fd_sc_hd__and3_1 _1902_ (.A(_0129_),
    .B(_0977_),
    .C(_0982_),
    .X(_0984_));
 sky130_fd_sc_hd__o31a_1 _1903_ (.A1(_0734_),
    .A2(_0983_),
    .A3(_0984_),
    .B1(_0808_),
    .X(_0985_));
 sky130_fd_sc_hd__xor2_2 _1904_ (.A(_0976_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__and2b_1 _1905_ (.A_N(_0947_),
    .B(_0958_),
    .X(_0987_));
 sky130_fd_sc_hd__a31oi_4 _1906_ (.A1(_0662_),
    .A2(_0940_),
    .A3(_0945_),
    .B1(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__xnor2_2 _1907_ (.A(_0986_),
    .B(_0988_),
    .Y(_0022_));
 sky130_fd_sc_hd__o21ba_1 _1908_ (.A1(_0927_),
    .A2(_0960_),
    .B1_N(_0961_),
    .X(_0023_));
 sky130_fd_sc_hd__a41o_1 _1909_ (.A1(_0930_),
    .A2(_0929_),
    .A3(_0931_),
    .A4(_0962_),
    .B1(_0023_),
    .X(_0024_));
 sky130_fd_sc_hd__xor2_2 _1910_ (.A(_0022_),
    .B(_0024_),
    .X(net17));
 sky130_fd_sc_hd__and2_1 _1911_ (.A(_0969_),
    .B(_0975_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _1912_ (.A(_0976_),
    .B(_0985_),
    .X(_0026_));
 sky130_fd_sc_hd__o21ai_1 _1913_ (.A1(_0861_),
    .A2(_0894_),
    .B1(_0909_),
    .Y(_0027_));
 sky130_fd_sc_hd__a21oi_1 _1914_ (.A1(_0833_),
    .A2(_0937_),
    .B1(_0845_),
    .Y(_0028_));
 sky130_fd_sc_hd__a21oi_1 _1915_ (.A1(_0027_),
    .A2(_0028_),
    .B1(_0902_),
    .Y(_0029_));
 sky130_fd_sc_hd__a311oi_2 _1916_ (.A1(_0756_),
    .A2(_0027_),
    .A3(_0028_),
    .B1(_0029_),
    .C1(_0758_),
    .Y(_0030_));
 sky130_fd_sc_hd__a31o_1 _1917_ (.A1(_0845_),
    .A2(_0839_),
    .A3(_0861_),
    .B1(_0935_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(\p_shaping_I.p_shaping_I.bit_in ),
    .A1(_0906_),
    .S(_0032_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(_0030_),
    .B(_0033_),
    .Y(_0034_));
 sky130_fd_sc_hd__or2_1 _1920_ (.A(_0030_),
    .B(_0033_),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(_0034_),
    .B(_0035_),
    .Y(_0036_));
 sky130_fd_sc_hd__o211a_1 _1922_ (.A1(_0622_),
    .A2(_0837_),
    .B1(_0669_),
    .C1(_0917_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_0835_),
    .B(_0656_),
    .Y(_0038_));
 sky130_fd_sc_hd__o22a_1 _1924_ (.A1(_0835_),
    .A2(_0965_),
    .B1(_0037_),
    .B2(_0038_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_1 _1925_ (.A(_0751_),
    .B(_0039_),
    .Y(_0040_));
 sky130_fd_sc_hd__a211o_1 _1926_ (.A1(_0129_),
    .A2(_0039_),
    .B1(_0040_),
    .C1(_0734_),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _1927_ (.A(_0808_),
    .B(_0041_),
    .X(_0043_));
 sky130_fd_sc_hd__xnor2_1 _1928_ (.A(_0036_),
    .B(_0043_),
    .Y(_0044_));
 sky130_fd_sc_hd__o21ai_1 _1929_ (.A1(_0025_),
    .A2(_0026_),
    .B1(_0044_),
    .Y(_0045_));
 sky130_fd_sc_hd__or3_1 _1930_ (.A(_0025_),
    .B(_0026_),
    .C(_0044_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _1931_ (.A(_0045_),
    .B(_0046_),
    .X(_0047_));
 sky130_fd_sc_hd__or2b_1 _1932_ (.A(_0988_),
    .B_N(_0986_),
    .X(_0048_));
 sky130_fd_sc_hd__a21bo_1 _1933_ (.A1(_0022_),
    .A2(_0024_),
    .B1_N(_0048_),
    .X(_0049_));
 sky130_fd_sc_hd__xor2_2 _1934_ (.A(_0047_),
    .B(_0049_),
    .X(net18));
 sky130_fd_sc_hd__o21a_1 _1935_ (.A1(_0626_),
    .A2(_0650_),
    .B1(_0028_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _1936_ (.A(_0902_),
    .B(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _1937_ (.A(_0756_),
    .B(_0050_),
    .Y(_0052_));
 sky130_fd_sc_hd__mux2_1 _1938_ (.A0(\p_shaping_I.p_shaping_I.bit_in ),
    .A1(_0906_),
    .S(_0935_),
    .X(_0053_));
 sky130_fd_sc_hd__nand4_2 _1939_ (.A(_0662_),
    .B(_0051_),
    .C(_0052_),
    .D(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__a31o_1 _1940_ (.A1(_0662_),
    .A2(_0051_),
    .A3(_0052_),
    .B1(_0053_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_2 _1941_ (.A(_0054_),
    .B(_0055_),
    .Y(_0056_));
 sky130_fd_sc_hd__o21a_1 _1942_ (.A1(_0736_),
    .A2(_0638_),
    .B1(_0909_),
    .X(_0057_));
 sky130_fd_sc_hd__o2bb2a_1 _1943_ (.A1_N(_0674_),
    .A2_N(_0866_),
    .B1(_0057_),
    .B2(_0835_),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _1944_ (.A(_0734_),
    .B(_0751_),
    .X(_0059_));
 sky130_fd_sc_hd__nand2_1 _1945_ (.A(_0752_),
    .B(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__o21ai_1 _1946_ (.A1(_0058_),
    .A2(_0060_),
    .B1(_0021_),
    .Y(_0061_));
 sky130_fd_sc_hd__a21oi_2 _1947_ (.A1(_0058_),
    .A2(_0060_),
    .B1(_0061_),
    .Y(_0063_));
 sky130_fd_sc_hd__xor2_4 _1948_ (.A(_0056_),
    .B(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__a21boi_4 _1949_ (.A1(_0035_),
    .A2(_0043_),
    .B1_N(_0034_),
    .Y(_0065_));
 sky130_fd_sc_hd__xnor2_4 _1950_ (.A(_0064_),
    .B(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__a21boi_1 _1951_ (.A1(_0048_),
    .A2(_0045_),
    .B1_N(_0046_),
    .Y(_0067_));
 sky130_fd_sc_hd__a31o_2 _1952_ (.A1(_0022_),
    .A2(_0024_),
    .A3(_0047_),
    .B1(_0067_),
    .X(_0068_));
 sky130_fd_sc_hd__xnor2_4 _1953_ (.A(_0066_),
    .B(_0068_),
    .Y(net7));
 sky130_fd_sc_hd__or2b_1 _1954_ (.A(_0056_),
    .B_N(_0063_),
    .X(_0069_));
 sky130_fd_sc_hd__clkinv_2 _1955_ (.A(_0129_),
    .Y(_0070_));
 sky130_fd_sc_hd__o21a_1 _1956_ (.A1(_0835_),
    .A2(_0650_),
    .B1(_0640_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1957_ (.A0(_0070_),
    .A1(_0751_),
    .S(_0071_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _1958_ (.A(_0808_),
    .Y(_0074_));
 sky130_fd_sc_hd__a21o_1 _1959_ (.A1(_0805_),
    .A2(_0073_),
    .B1(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__xnor2_1 _1960_ (.A(_0056_),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__a21o_1 _1961_ (.A1(_0054_),
    .A2(_0069_),
    .B1(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__nand3_1 _1962_ (.A(_0054_),
    .B(_0069_),
    .C(_0076_),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_2 _1963_ (.A(_0077_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1964_ (.A(_0066_),
    .Y(_0080_));
 sky130_fd_sc_hd__nor2_1 _1965_ (.A(_0064_),
    .B(_0065_),
    .Y(_0081_));
 sky130_fd_sc_hd__a21o_1 _1966_ (.A1(_0080_),
    .A2(_0068_),
    .B1(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__xnor2_4 _1967_ (.A(_0079_),
    .B(_0082_),
    .Y(net8));
 sky130_fd_sc_hd__nand4_1 _1968_ (.A(_0080_),
    .B(_0068_),
    .C(_0077_),
    .D(_0078_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand2_1 _1969_ (.A(_0081_),
    .B(_0078_),
    .Y(_0085_));
 sky130_fd_sc_hd__a21bo_1 _1970_ (.A1(_0055_),
    .A2(_0075_),
    .B1_N(_0054_),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_1 _1971_ (.A1(_0021_),
    .A2(_0060_),
    .B1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__and3_1 _1972_ (.A(_0021_),
    .B(_0060_),
    .C(_0086_),
    .X(_0088_));
 sky130_fd_sc_hd__a41o_1 _1973_ (.A1(_0077_),
    .A2(_0084_),
    .A3(_0085_),
    .A4(_0087_),
    .B1(_0088_),
    .X(net9));
 sky130_fd_sc_hd__xnor2_4 _1974_ (.A(_0775_),
    .B(_0773_),
    .Y(net10));
 sky130_fd_sc_hd__nand2_1 _1975_ (.A(\p_shaping_Q.p_shaping_I.counter[0] ),
    .B(_0362_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _1976_ (.A(_0007_),
    .B(_0089_),
    .Y(_0006_));
 sky130_fd_sc_hd__and2_1 _1977_ (.A(net50),
    .B(net3),
    .X(_0091_));
 sky130_fd_sc_hd__buf_2 _1978_ (.A(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _1979_ (.A(_0675_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__and3_1 _1980_ (.A(_0675_),
    .B(net50),
    .C(net3),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _1981_ (.A(_0093_),
    .B(_0094_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_2 _1982_ (.A(net50),
    .B(net3),
    .Y(_0095_));
 sky130_fd_sc_hd__nor2_1 _1983_ (.A(_0603_),
    .B(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__a22o_1 _1984_ (.A1(_0604_),
    .A2(_0095_),
    .B1(_0096_),
    .B2(_0042_),
    .X(_0009_));
 sky130_fd_sc_hd__or3_1 _1985_ (.A(_0679_),
    .B(_0638_),
    .C(_0095_),
    .X(_0097_));
 sky130_fd_sc_hd__o21ai_1 _1986_ (.A1(_0652_),
    .A2(_0092_),
    .B1(_0097_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(_0716_),
    .B(_0094_),
    .Y(_0099_));
 sky130_fd_sc_hd__o211a_1 _1988_ (.A1(_0736_),
    .A2(_0094_),
    .B1(_0099_),
    .C1(_0714_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1989_ (.A(_0654_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _1990_ (.A(_0654_),
    .B(_0099_),
    .Y(_0101_));
 sky130_fd_sc_hd__o211a_1 _1991_ (.A1(_0042_),
    .A2(_0095_),
    .B1(_0100_),
    .C1(_0101_),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_1 _1992_ (.A(_0835_),
    .B(_0100_),
    .Y(_0102_));
 sky130_fd_sc_hd__or2_1 _1993_ (.A(_0835_),
    .B(_0100_),
    .X(_0103_));
 sky130_fd_sc_hd__o211a_1 _1994_ (.A1(_0042_),
    .A2(_0095_),
    .B1(_0102_),
    .C1(_0103_),
    .X(_0013_));
 sky130_fd_sc_hd__xnor2_1 _1995_ (.A(_0121_),
    .B(_0092_),
    .Y(_0014_));
 sky130_fd_sc_hd__and2_1 _1996_ (.A(_0155_),
    .B(_0095_),
    .X(_0104_));
 sky130_fd_sc_hd__a31o_1 _1997_ (.A1(_0126_),
    .A2(_0204_),
    .A3(_0092_),
    .B1(_0104_),
    .X(_0015_));
 sky130_fd_sc_hd__or3_1 _1998_ (.A(_0163_),
    .B(_0161_),
    .C(_0095_),
    .X(_0106_));
 sky130_fd_sc_hd__a21bo_1 _1999_ (.A1(_0298_),
    .A2(_0095_),
    .B1_N(_0106_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_1 _2000_ (.A(_0365_),
    .B(_0163_),
    .C(_0092_),
    .X(_0107_));
 sky130_fd_sc_hd__a21oi_1 _2001_ (.A1(_0163_),
    .A2(_0092_),
    .B1(_0365_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_1 _2002_ (.A(_0107_),
    .B(_0108_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _2003_ (.A(_0449_),
    .B(_0107_),
    .Y(_0109_));
 sky130_fd_sc_hd__or2_1 _2004_ (.A(_0449_),
    .B(_0107_),
    .X(_0110_));
 sky130_fd_sc_hd__o211a_1 _2005_ (.A1(_0126_),
    .A2(_0095_),
    .B1(_0109_),
    .C1(_0110_),
    .X(_0018_));
 sky130_fd_sc_hd__xnor2_1 _2006_ (.A(_0202_),
    .B(_0109_),
    .Y(_0111_));
 sky130_fd_sc_hd__a21oi_1 _2007_ (.A1(_0005_),
    .A2(_0092_),
    .B1(_0111_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_1 _2008_ (.A(_0662_),
    .B(\p_shaping_I.p_shaping_I.counter[0] ),
    .Y(_0113_));
 sky130_fd_sc_hd__nand2_1 _2009_ (.A(_0021_),
    .B(_0113_),
    .Y(_0020_));
 sky130_fd_sc_hd__dfrtp_1 _2010_ (.CLK(_0005_),
    .D(_0006_),
    .RESET_B(net46),
    .Q(\p_shaping_Q.p_shaping_I.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2011_ (.CLK(_0005_),
    .D(_0007_),
    .RESET_B(net46),
    .Q(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2012_ (.CLK(_0004_),
    .D(\gen_sym.Reg_2M.data_in ),
    .RESET_B(net46),
    .Q(\gen_sym.Reg_Sym.data_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2013_ (.CLK(_0004_),
    .D(\gen_sym.Reg_2M.data_out ),
    .RESET_B(net47),
    .Q(\gen_sym.Reg_Sym.data_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2014_ (.CLK(\gen_sym.Reg_2M.enable ),
    .D(\gen_sym.Reg_2M.data_in ),
    .RESET_B(net46),
    .Q(\gen_sym.Reg_2M.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _2015_ (.CLK(_0005_),
    .D(\mapper.bit_Q[1] ),
    .RESET_B(net47),
    .Q(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__dfrtp_4 _2016_ (.CLK(_0004_),
    .D(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .RESET_B(net49),
    .Q(\p_shaping_I.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__dlxtn_1 _2017_ (.D(_0000_),
    .GATE_N(_0001_),
    .Q(\p_shaping_I.p_shaping_I.ctl_1 ));
 sky130_fd_sc_hd__dfrtp_4 _2018_ (.CLK(net50),
    .D(_0008_),
    .RESET_B(net47),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_4 _2019_ (.CLK(net50),
    .D(_0009_),
    .RESET_B(net47),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _2020_ (.CLK(net50),
    .D(_0010_),
    .RESET_B(net47),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_4 _2021_ (.CLK(net50),
    .D(_0011_),
    .RESET_B(net47),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_4 _2022_ (.CLK(net50),
    .D(_0012_),
    .RESET_B(net47),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_4 _2023_ (.CLK(net50),
    .D(_0013_),
    .RESET_B(net47),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _2024_ (.CLK(_0004_),
    .D(\p_shaping_I.p_shaping_I.bit_in ),
    .RESET_B(net49),
    .Q(\p_shaping_I.p_shaping_I.bit_in_1 ));
 sky130_fd_sc_hd__dfrtp_4 _2025_ (.CLK(_0005_),
    .D(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .RESET_B(net46),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__dlxtn_1 _2026_ (.D(_0002_),
    .GATE_N(_0003_),
    .Q(\p_shaping_Q.p_shaping_I.ctl_1 ));
 sky130_fd_sc_hd__dfstp_4 _2027_ (.CLK(net51),
    .D(_0014_),
    .SET_B(net48),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _2028_ (.CLK(net51),
    .D(_0015_),
    .RESET_B(net48),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_4 _2029_ (.CLK(net51),
    .D(_0016_),
    .RESET_B(net48),
    .Q(net40));
 sky130_fd_sc_hd__dfstp_4 _2030_ (.CLK(net51),
    .D(_0017_),
    .SET_B(net48),
    .Q(net41));
 sky130_fd_sc_hd__dfstp_4 _2031_ (.CLK(net51),
    .D(_0018_),
    .SET_B(net48),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_4 _2032_ (.CLK(net50),
    .D(_0019_),
    .RESET_B(net47),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _2033_ (.CLK(_0005_),
    .D(\p_shaping_Q.p_shaping_I.bit_in ),
    .RESET_B(net46),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 sky130_fd_sc_hd__dfrtp_1 _2034_ (.CLK(_0004_),
    .D(_0020_),
    .RESET_B(net49),
    .Q(\p_shaping_I.p_shaping_I.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2035_ (.CLK(_0004_),
    .D(_0021_),
    .RESET_B(net49),
    .Q(\p_shaping_I.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ACK),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(Bit_In),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(EN),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(REQ_SAMPLE),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(RST),
    .X(net5));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(I[0]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(I[10]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(I[11]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(I[12]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(I[1]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(I[2]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(I[3]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(I[4]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(I[5]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(I[6]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(I[7]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(I[8]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(I[9]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(Q[0]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(Q[10]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(Q[11]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(Q[12]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(Q[1]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(Q[2]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(Q[3]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(Q[4]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(Q[5]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(Q[6]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(Q[7]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(Q[8]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(Q[9]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(addI[0]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(addI[1]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(addI[2]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(addI[3]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(addI[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(addI[5]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(addQ[0]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(addQ[1]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(addQ[2]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(addQ[3]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(addQ[4]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(addQ[5]));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net39),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net34),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net48),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net5),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net4),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout51 (.A(net4),
    .X(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ACK));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(Bit_In));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(EN));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(REQ_SAMPLE));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(RST));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__D (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__A1 (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__B1 (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__C1 (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__B1 (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__C1 (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__B_N (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1 (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__A1 (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__B2 (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__A (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__B (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__A (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__S (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A (.DIODE(_0042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A2 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__A2 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__C (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A3 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__B (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A2 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__B (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A3 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A3 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A2 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A1 (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A1 (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__A (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__S (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__B1 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__A (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__C (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__B1 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__B1 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__B (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__A2 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__A1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__A (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__A (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__B2 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A1 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__A1 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__A1 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__B1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__C1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__C1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__C1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__B2 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__A1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__C1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__A3 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__B (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__A (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__B1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__B (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__C1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__B2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__B1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__A2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__B1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__A2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A3 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__A2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__C (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__C1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__A3 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__A2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__B1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__B1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__B (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__B1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__A1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__A (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A3 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__A (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__A (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__A (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__B (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__C1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__A (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__C1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__A (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A2 (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__A2 (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__B (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__C1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__B (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A2 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__C (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__A2 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__B1 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A3 (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A3 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__C (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__B1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__C1 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A3 (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__A1_N (.DIODE(_0641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__C1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__C_N (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A1 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__D_N (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__B (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__B1 (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A_N (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__B (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__B2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__B2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__B2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__D (.DIODE(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__B (.DIODE(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__B1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A (.DIODE(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__A (.DIODE(\p_shaping_Q.p_shaping_I.bit_in ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__A1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__A (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__A1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__B1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__A1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A1 (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (.DIODE(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__B1_N (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__C_N (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__B (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__A (.DIODE(\p_shaping_Q.p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__C (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output6_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_output7_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_output8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_output9_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__B1_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__A_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__C (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__B1_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__SET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__SET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__SET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__S (.DIODE(net49));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
endmodule

