magic
tech sky130A
magscale 1 2
timestamp 1671750181
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 14 2128 59970 57712
<< metal2 >>
rect 2594 59200 2650 59800
rect 8390 59200 8446 59800
rect 13542 59200 13598 59800
rect 19338 59200 19394 59800
rect 24490 59200 24546 59800
rect 30286 59200 30342 59800
rect 35438 59200 35494 59800
rect 41234 59200 41290 59800
rect 46386 59200 46442 59800
rect 52182 59200 52238 59800
rect 57334 59200 57390 59800
rect 18 200 74 800
rect 5170 200 5226 800
rect 10966 200 11022 800
rect 16118 200 16174 800
rect 21914 200 21970 800
rect 27066 200 27122 800
rect 32862 200 32918 800
rect 38014 200 38070 800
rect 43810 200 43866 800
rect 48962 200 49018 800
rect 54758 200 54814 800
rect 59910 200 59966 800
<< obsm2 >>
rect 20 59144 2538 59200
rect 2706 59144 8334 59200
rect 8502 59144 13486 59200
rect 13654 59144 19282 59200
rect 19450 59144 24434 59200
rect 24602 59144 30230 59200
rect 30398 59144 35382 59200
rect 35550 59144 41178 59200
rect 41346 59144 46330 59200
rect 46498 59144 52126 59200
rect 52294 59144 57278 59200
rect 57446 59144 59964 59200
rect 20 856 59964 59144
rect 130 734 5114 856
rect 5282 734 10910 856
rect 11078 734 16062 856
rect 16230 734 21858 856
rect 22026 734 27010 856
rect 27178 734 32806 856
rect 32974 734 37958 856
rect 38126 734 43754 856
rect 43922 734 48906 856
rect 49074 734 54702 856
rect 54870 734 59854 856
<< metal3 >>
rect 200 57808 800 57928
rect 59200 57128 59800 57248
rect 200 51688 800 51808
rect 59200 51688 59800 51808
rect 200 46248 800 46368
rect 59200 45568 59800 45688
rect 200 40128 800 40248
rect 59200 40128 59800 40248
rect 200 34688 800 34808
rect 59200 34008 59800 34128
rect 200 28568 800 28688
rect 59200 28568 59800 28688
rect 200 23128 800 23248
rect 59200 22448 59800 22568
rect 200 17008 800 17128
rect 59200 17008 59800 17128
rect 200 11568 800 11688
rect 59200 10888 59800 11008
rect 200 5448 800 5568
rect 59200 5448 59800 5568
<< obsm3 >>
rect 880 57728 59200 57901
rect 800 57328 59200 57728
rect 800 57048 59120 57328
rect 800 51888 59200 57048
rect 880 51608 59120 51888
rect 800 46448 59200 51608
rect 880 46168 59200 46448
rect 800 45768 59200 46168
rect 800 45488 59120 45768
rect 800 40328 59200 45488
rect 880 40048 59120 40328
rect 800 34888 59200 40048
rect 880 34608 59200 34888
rect 800 34208 59200 34608
rect 800 33928 59120 34208
rect 800 28768 59200 33928
rect 880 28488 59120 28768
rect 800 23328 59200 28488
rect 880 23048 59200 23328
rect 800 22648 59200 23048
rect 800 22368 59120 22648
rect 800 17208 59200 22368
rect 880 16928 59120 17208
rect 800 11768 59200 16928
rect 880 11488 59200 11768
rect 800 11088 59200 11488
rect 800 10808 59120 11088
rect 800 5648 59200 10808
rect 880 5368 59120 5648
rect 800 2143 59200 5368
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 22139 2483 34848 56677
rect 35328 2483 44653 56677
<< labels >>
rlabel metal2 s 30286 59200 30342 59800 6 ACK
port 1 nsew signal input
rlabel metal2 s 2594 59200 2650 59800 6 Bit_In
port 2 nsew signal input
rlabel metal2 s 43810 200 43866 800 6 EN
port 3 nsew signal input
rlabel metal3 s 59200 5448 59800 5568 6 I[0]
port 4 nsew signal output
rlabel metal3 s 200 46248 800 46368 6 I[10]
port 5 nsew signal output
rlabel metal2 s 59910 200 59966 800 6 I[11]
port 6 nsew signal output
rlabel metal2 s 54758 200 54814 800 6 I[12]
port 7 nsew signal output
rlabel metal3 s 59200 40128 59800 40248 6 I[1]
port 8 nsew signal output
rlabel metal2 s 21914 200 21970 800 6 I[2]
port 9 nsew signal output
rlabel metal2 s 32862 200 32918 800 6 I[3]
port 10 nsew signal output
rlabel metal2 s 46386 59200 46442 59800 6 I[4]
port 11 nsew signal output
rlabel metal3 s 200 23128 800 23248 6 I[5]
port 12 nsew signal output
rlabel metal3 s 59200 45568 59800 45688 6 I[6]
port 13 nsew signal output
rlabel metal3 s 200 34688 800 34808 6 I[7]
port 14 nsew signal output
rlabel metal2 s 10966 200 11022 800 6 I[8]
port 15 nsew signal output
rlabel metal3 s 200 40128 800 40248 6 I[9]
port 16 nsew signal output
rlabel metal3 s 200 17008 800 17128 6 Q[0]
port 17 nsew signal output
rlabel metal2 s 35438 59200 35494 59800 6 Q[10]
port 18 nsew signal output
rlabel metal2 s 52182 59200 52238 59800 6 Q[11]
port 19 nsew signal output
rlabel metal3 s 59200 17008 59800 17128 6 Q[12]
port 20 nsew signal output
rlabel metal3 s 59200 51688 59800 51808 6 Q[1]
port 21 nsew signal output
rlabel metal2 s 13542 59200 13598 59800 6 Q[2]
port 22 nsew signal output
rlabel metal2 s 18 200 74 800 6 Q[3]
port 23 nsew signal output
rlabel metal3 s 200 11568 800 11688 6 Q[4]
port 24 nsew signal output
rlabel metal3 s 59200 34008 59800 34128 6 Q[5]
port 25 nsew signal output
rlabel metal2 s 8390 59200 8446 59800 6 Q[6]
port 26 nsew signal output
rlabel metal3 s 200 5448 800 5568 6 Q[7]
port 27 nsew signal output
rlabel metal2 s 48962 200 49018 800 6 Q[8]
port 28 nsew signal output
rlabel metal2 s 41234 59200 41290 59800 6 Q[9]
port 29 nsew signal output
rlabel metal3 s 59200 10888 59800 11008 6 REQ_SAMPLE
port 30 nsew signal input
rlabel metal2 s 5170 200 5226 800 6 RST
port 31 nsew signal input
rlabel metal2 s 16118 200 16174 800 6 addI[0]
port 32 nsew signal output
rlabel metal3 s 200 51688 800 51808 6 addI[1]
port 33 nsew signal output
rlabel metal3 s 59200 22448 59800 22568 6 addI[2]
port 34 nsew signal output
rlabel metal2 s 27066 200 27122 800 6 addI[3]
port 35 nsew signal output
rlabel metal3 s 59200 57128 59800 57248 6 addI[4]
port 36 nsew signal output
rlabel metal2 s 57334 59200 57390 59800 6 addI[5]
port 37 nsew signal output
rlabel metal2 s 19338 59200 19394 59800 6 addQ[0]
port 38 nsew signal output
rlabel metal2 s 24490 59200 24546 59800 6 addQ[1]
port 39 nsew signal output
rlabel metal2 s 38014 200 38070 800 6 addQ[2]
port 40 nsew signal output
rlabel metal3 s 200 28568 800 28688 6 addQ[3]
port 41 nsew signal output
rlabel metal3 s 200 57808 800 57928 6 addQ[4]
port 42 nsew signal output
rlabel metal3 s 59200 28568 59800 28688 6 addQ[5]
port 43 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4765790
string GDS_FILE /home/urielcho/Proyectos_caravel/MPW8/gf180_vs_sky130/openlane/modulador_a/runs/22_12_22_17_00/results/signoff/OQPSK_RCOSINE_ALL.magic.gds
string GDS_START 948680
<< end >>

