magic
tech sky130A
magscale 1 2
timestamp 1671747965
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 14 1844 299538 297696
<< metal2 >>
rect 1950 299200 2006 299800
rect 4526 299200 4582 299800
rect 7746 299200 7802 299800
rect 10966 299200 11022 299800
rect 13542 299200 13598 299800
rect 16762 299200 16818 299800
rect 19338 299200 19394 299800
rect 22558 299200 22614 299800
rect 25134 299200 25190 299800
rect 28354 299200 28410 299800
rect 30930 299200 30986 299800
rect 34150 299200 34206 299800
rect 36726 299200 36782 299800
rect 39946 299200 40002 299800
rect 42522 299200 42578 299800
rect 45742 299200 45798 299800
rect 48318 299200 48374 299800
rect 51538 299200 51594 299800
rect 54758 299200 54814 299800
rect 57334 299200 57390 299800
rect 60554 299200 60610 299800
rect 63130 299200 63186 299800
rect 66350 299200 66406 299800
rect 68926 299200 68982 299800
rect 72146 299200 72202 299800
rect 74722 299200 74778 299800
rect 77942 299200 77998 299800
rect 80518 299200 80574 299800
rect 83738 299200 83794 299800
rect 86314 299200 86370 299800
rect 89534 299200 89590 299800
rect 92754 299200 92810 299800
rect 95330 299200 95386 299800
rect 98550 299200 98606 299800
rect 101126 299200 101182 299800
rect 104346 299200 104402 299800
rect 106922 299200 106978 299800
rect 110142 299200 110198 299800
rect 112718 299200 112774 299800
rect 115938 299200 115994 299800
rect 118514 299200 118570 299800
rect 121734 299200 121790 299800
rect 124310 299200 124366 299800
rect 127530 299200 127586 299800
rect 130106 299200 130162 299800
rect 133326 299200 133382 299800
rect 136546 299200 136602 299800
rect 139122 299200 139178 299800
rect 142342 299200 142398 299800
rect 144918 299200 144974 299800
rect 148138 299200 148194 299800
rect 150714 299200 150770 299800
rect 153934 299200 153990 299800
rect 156510 299200 156566 299800
rect 159730 299200 159786 299800
rect 162306 299200 162362 299800
rect 165526 299200 165582 299800
rect 168102 299200 168158 299800
rect 171322 299200 171378 299800
rect 173898 299200 173954 299800
rect 177118 299200 177174 299800
rect 180338 299200 180394 299800
rect 182914 299200 182970 299800
rect 186134 299200 186190 299800
rect 188710 299200 188766 299800
rect 191930 299200 191986 299800
rect 194506 299200 194562 299800
rect 197726 299200 197782 299800
rect 200302 299200 200358 299800
rect 203522 299200 203578 299800
rect 206098 299200 206154 299800
rect 209318 299200 209374 299800
rect 211894 299200 211950 299800
rect 215114 299200 215170 299800
rect 218334 299200 218390 299800
rect 220910 299200 220966 299800
rect 224130 299200 224186 299800
rect 226706 299200 226762 299800
rect 229926 299200 229982 299800
rect 232502 299200 232558 299800
rect 235722 299200 235778 299800
rect 238298 299200 238354 299800
rect 241518 299200 241574 299800
rect 244094 299200 244150 299800
rect 247314 299200 247370 299800
rect 249890 299200 249946 299800
rect 253110 299200 253166 299800
rect 255686 299200 255742 299800
rect 258906 299200 258962 299800
rect 262126 299200 262182 299800
rect 264702 299200 264758 299800
rect 267922 299200 267978 299800
rect 270498 299200 270554 299800
rect 273718 299200 273774 299800
rect 276294 299200 276350 299800
rect 279514 299200 279570 299800
rect 282090 299200 282146 299800
rect 285310 299200 285366 299800
rect 287886 299200 287942 299800
rect 291106 299200 291162 299800
rect 293682 299200 293738 299800
rect 296902 299200 296958 299800
rect 299478 299200 299534 299800
rect 18 200 74 800
rect 2594 200 2650 800
rect 5814 200 5870 800
rect 8390 200 8446 800
rect 11610 200 11666 800
rect 14186 200 14242 800
rect 17406 200 17462 800
rect 19982 200 20038 800
rect 23202 200 23258 800
rect 25778 200 25834 800
rect 28998 200 29054 800
rect 31574 200 31630 800
rect 34794 200 34850 800
rect 37370 200 37426 800
rect 40590 200 40646 800
rect 43810 200 43866 800
rect 46386 200 46442 800
rect 49606 200 49662 800
rect 52182 200 52238 800
rect 55402 200 55458 800
rect 57978 200 58034 800
rect 61198 200 61254 800
rect 63774 200 63830 800
rect 66994 200 67050 800
rect 69570 200 69626 800
rect 72790 200 72846 800
rect 75366 200 75422 800
rect 78586 200 78642 800
rect 81162 200 81218 800
rect 84382 200 84438 800
rect 87602 200 87658 800
rect 90178 200 90234 800
rect 93398 200 93454 800
rect 95974 200 96030 800
rect 99194 200 99250 800
rect 101770 200 101826 800
rect 104990 200 105046 800
rect 107566 200 107622 800
rect 110786 200 110842 800
rect 113362 200 113418 800
rect 116582 200 116638 800
rect 119158 200 119214 800
rect 122378 200 122434 800
rect 125598 200 125654 800
rect 128174 200 128230 800
rect 131394 200 131450 800
rect 133970 200 134026 800
rect 137190 200 137246 800
rect 139766 200 139822 800
rect 142986 200 143042 800
rect 145562 200 145618 800
rect 148782 200 148838 800
rect 151358 200 151414 800
rect 154578 200 154634 800
rect 157154 200 157210 800
rect 160374 200 160430 800
rect 162950 200 163006 800
rect 166170 200 166226 800
rect 169390 200 169446 800
rect 171966 200 172022 800
rect 175186 200 175242 800
rect 177762 200 177818 800
rect 180982 200 181038 800
rect 183558 200 183614 800
rect 186778 200 186834 800
rect 189354 200 189410 800
rect 192574 200 192630 800
rect 195150 200 195206 800
rect 198370 200 198426 800
rect 200946 200 201002 800
rect 204166 200 204222 800
rect 206742 200 206798 800
rect 209962 200 210018 800
rect 213182 200 213238 800
rect 215758 200 215814 800
rect 218978 200 219034 800
rect 221554 200 221610 800
rect 224774 200 224830 800
rect 227350 200 227406 800
rect 230570 200 230626 800
rect 233146 200 233202 800
rect 236366 200 236422 800
rect 238942 200 238998 800
rect 242162 200 242218 800
rect 244738 200 244794 800
rect 247958 200 248014 800
rect 251178 200 251234 800
rect 253754 200 253810 800
rect 256974 200 257030 800
rect 259550 200 259606 800
rect 262770 200 262826 800
rect 265346 200 265402 800
rect 268566 200 268622 800
rect 271142 200 271198 800
rect 274362 200 274418 800
rect 276938 200 276994 800
rect 280158 200 280214 800
rect 282734 200 282790 800
rect 285954 200 286010 800
rect 288530 200 288586 800
rect 291750 200 291806 800
rect 294970 200 295026 800
rect 297546 200 297602 800
<< obsm2 >>
rect 20 299144 1894 299282
rect 2062 299144 4470 299282
rect 4638 299144 7690 299282
rect 7858 299144 10910 299282
rect 11078 299144 13486 299282
rect 13654 299144 16706 299282
rect 16874 299144 19282 299282
rect 19450 299144 22502 299282
rect 22670 299144 25078 299282
rect 25246 299144 28298 299282
rect 28466 299144 30874 299282
rect 31042 299144 34094 299282
rect 34262 299144 36670 299282
rect 36838 299144 39890 299282
rect 40058 299144 42466 299282
rect 42634 299144 45686 299282
rect 45854 299144 48262 299282
rect 48430 299144 51482 299282
rect 51650 299144 54702 299282
rect 54870 299144 57278 299282
rect 57446 299144 60498 299282
rect 60666 299144 63074 299282
rect 63242 299144 66294 299282
rect 66462 299144 68870 299282
rect 69038 299144 72090 299282
rect 72258 299144 74666 299282
rect 74834 299144 77886 299282
rect 78054 299144 80462 299282
rect 80630 299144 83682 299282
rect 83850 299144 86258 299282
rect 86426 299144 89478 299282
rect 89646 299144 92698 299282
rect 92866 299144 95274 299282
rect 95442 299144 98494 299282
rect 98662 299144 101070 299282
rect 101238 299144 104290 299282
rect 104458 299144 106866 299282
rect 107034 299144 110086 299282
rect 110254 299144 112662 299282
rect 112830 299144 115882 299282
rect 116050 299144 118458 299282
rect 118626 299144 121678 299282
rect 121846 299144 124254 299282
rect 124422 299144 127474 299282
rect 127642 299144 130050 299282
rect 130218 299144 133270 299282
rect 133438 299144 136490 299282
rect 136658 299144 139066 299282
rect 139234 299144 142286 299282
rect 142454 299144 144862 299282
rect 145030 299144 148082 299282
rect 148250 299144 150658 299282
rect 150826 299144 153878 299282
rect 154046 299144 156454 299282
rect 156622 299144 159674 299282
rect 159842 299144 162250 299282
rect 162418 299144 165470 299282
rect 165638 299144 168046 299282
rect 168214 299144 171266 299282
rect 171434 299144 173842 299282
rect 174010 299144 177062 299282
rect 177230 299144 180282 299282
rect 180450 299144 182858 299282
rect 183026 299144 186078 299282
rect 186246 299144 188654 299282
rect 188822 299144 191874 299282
rect 192042 299144 194450 299282
rect 194618 299144 197670 299282
rect 197838 299144 200246 299282
rect 200414 299144 203466 299282
rect 203634 299144 206042 299282
rect 206210 299144 209262 299282
rect 209430 299144 211838 299282
rect 212006 299144 215058 299282
rect 215226 299144 218278 299282
rect 218446 299144 220854 299282
rect 221022 299144 224074 299282
rect 224242 299144 226650 299282
rect 226818 299144 229870 299282
rect 230038 299144 232446 299282
rect 232614 299144 235666 299282
rect 235834 299144 238242 299282
rect 238410 299144 241462 299282
rect 241630 299144 244038 299282
rect 244206 299144 247258 299282
rect 247426 299144 249834 299282
rect 250002 299144 253054 299282
rect 253222 299144 255630 299282
rect 255798 299144 258850 299282
rect 259018 299144 262070 299282
rect 262238 299144 264646 299282
rect 264814 299144 267866 299282
rect 268034 299144 270442 299282
rect 270610 299144 273662 299282
rect 273830 299144 276238 299282
rect 276406 299144 279458 299282
rect 279626 299144 282034 299282
rect 282202 299144 285254 299282
rect 285422 299144 287830 299282
rect 287998 299144 291050 299282
rect 291218 299144 293626 299282
rect 293794 299144 296846 299282
rect 297014 299144 299422 299282
rect 20 856 299532 299144
rect 130 711 2538 856
rect 2706 711 5758 856
rect 5926 711 8334 856
rect 8502 711 11554 856
rect 11722 711 14130 856
rect 14298 711 17350 856
rect 17518 711 19926 856
rect 20094 711 23146 856
rect 23314 711 25722 856
rect 25890 711 28942 856
rect 29110 711 31518 856
rect 31686 711 34738 856
rect 34906 711 37314 856
rect 37482 711 40534 856
rect 40702 711 43754 856
rect 43922 711 46330 856
rect 46498 711 49550 856
rect 49718 711 52126 856
rect 52294 711 55346 856
rect 55514 711 57922 856
rect 58090 711 61142 856
rect 61310 711 63718 856
rect 63886 711 66938 856
rect 67106 711 69514 856
rect 69682 711 72734 856
rect 72902 711 75310 856
rect 75478 711 78530 856
rect 78698 711 81106 856
rect 81274 711 84326 856
rect 84494 711 87546 856
rect 87714 711 90122 856
rect 90290 711 93342 856
rect 93510 711 95918 856
rect 96086 711 99138 856
rect 99306 711 101714 856
rect 101882 711 104934 856
rect 105102 711 107510 856
rect 107678 711 110730 856
rect 110898 711 113306 856
rect 113474 711 116526 856
rect 116694 711 119102 856
rect 119270 711 122322 856
rect 122490 711 125542 856
rect 125710 711 128118 856
rect 128286 711 131338 856
rect 131506 711 133914 856
rect 134082 711 137134 856
rect 137302 711 139710 856
rect 139878 711 142930 856
rect 143098 711 145506 856
rect 145674 711 148726 856
rect 148894 711 151302 856
rect 151470 711 154522 856
rect 154690 711 157098 856
rect 157266 711 160318 856
rect 160486 711 162894 856
rect 163062 711 166114 856
rect 166282 711 169334 856
rect 169502 711 171910 856
rect 172078 711 175130 856
rect 175298 711 177706 856
rect 177874 711 180926 856
rect 181094 711 183502 856
rect 183670 711 186722 856
rect 186890 711 189298 856
rect 189466 711 192518 856
rect 192686 711 195094 856
rect 195262 711 198314 856
rect 198482 711 200890 856
rect 201058 711 204110 856
rect 204278 711 206686 856
rect 206854 711 209906 856
rect 210074 711 213126 856
rect 213294 711 215702 856
rect 215870 711 218922 856
rect 219090 711 221498 856
rect 221666 711 224718 856
rect 224886 711 227294 856
rect 227462 711 230514 856
rect 230682 711 233090 856
rect 233258 711 236310 856
rect 236478 711 238886 856
rect 239054 711 242106 856
rect 242274 711 244682 856
rect 244850 711 247902 856
rect 248070 711 251122 856
rect 251290 711 253698 856
rect 253866 711 256918 856
rect 257086 711 259494 856
rect 259662 711 262714 856
rect 262882 711 265290 856
rect 265458 711 268510 856
rect 268678 711 271086 856
rect 271254 711 274306 856
rect 274474 711 276882 856
rect 277050 711 280102 856
rect 280270 711 282678 856
rect 282846 711 285898 856
rect 286066 711 288474 856
rect 288642 711 291694 856
rect 291862 711 294914 856
rect 295082 711 297490 856
rect 297658 711 299532 856
<< metal3 >>
rect 200 298528 800 298648
rect 299200 296488 299800 296608
rect 200 295808 800 295928
rect 299200 293088 299800 293208
rect 200 292408 800 292528
rect 299200 290368 299800 290488
rect 200 289688 800 289808
rect 299200 286968 299800 287088
rect 200 286288 800 286408
rect 299200 284248 299800 284368
rect 200 283568 800 283688
rect 299200 280848 299800 280968
rect 200 280168 800 280288
rect 299200 278128 299800 278248
rect 200 277448 800 277568
rect 299200 274728 299800 274848
rect 200 274048 800 274168
rect 299200 272008 299800 272128
rect 200 271328 800 271448
rect 299200 268608 299800 268728
rect 200 267928 800 268048
rect 299200 265888 299800 266008
rect 200 265208 800 265328
rect 299200 262488 299800 262608
rect 200 261808 800 261928
rect 299200 259768 299800 259888
rect 200 258408 800 258528
rect 299200 256368 299800 256488
rect 200 255688 800 255808
rect 299200 252968 299800 253088
rect 200 252288 800 252408
rect 299200 250248 299800 250368
rect 200 249568 800 249688
rect 299200 246848 299800 246968
rect 200 246168 800 246288
rect 299200 244128 299800 244248
rect 200 243448 800 243568
rect 299200 240728 299800 240848
rect 200 240048 800 240168
rect 299200 238008 299800 238128
rect 200 237328 800 237448
rect 299200 234608 299800 234728
rect 200 233928 800 234048
rect 299200 231888 299800 232008
rect 200 231208 800 231328
rect 299200 228488 299800 228608
rect 200 227808 800 227928
rect 299200 225768 299800 225888
rect 200 225088 800 225208
rect 299200 222368 299800 222488
rect 200 221688 800 221808
rect 299200 219648 299800 219768
rect 200 218288 800 218408
rect 299200 216248 299800 216368
rect 200 215568 800 215688
rect 299200 213528 299800 213648
rect 200 212168 800 212288
rect 299200 210128 299800 210248
rect 200 209448 800 209568
rect 299200 206728 299800 206848
rect 200 206048 800 206168
rect 299200 204008 299800 204128
rect 200 203328 800 203448
rect 299200 200608 299800 200728
rect 200 199928 800 200048
rect 299200 197888 299800 198008
rect 200 197208 800 197328
rect 299200 194488 299800 194608
rect 200 193808 800 193928
rect 299200 191768 299800 191888
rect 200 191088 800 191208
rect 299200 188368 299800 188488
rect 200 187688 800 187808
rect 299200 185648 299800 185768
rect 200 184968 800 185088
rect 299200 182248 299800 182368
rect 200 181568 800 181688
rect 299200 179528 299800 179648
rect 200 178848 800 178968
rect 299200 176128 299800 176248
rect 200 175448 800 175568
rect 299200 173408 299800 173528
rect 200 172048 800 172168
rect 299200 170008 299800 170128
rect 200 169328 800 169448
rect 299200 166608 299800 166728
rect 200 165928 800 166048
rect 299200 163888 299800 164008
rect 200 163208 800 163328
rect 299200 160488 299800 160608
rect 200 159808 800 159928
rect 299200 157768 299800 157888
rect 200 157088 800 157208
rect 299200 154368 299800 154488
rect 200 153688 800 153808
rect 299200 151648 299800 151768
rect 200 150968 800 151088
rect 299200 148248 299800 148368
rect 200 147568 800 147688
rect 299200 145528 299800 145648
rect 200 144848 800 144968
rect 299200 142128 299800 142248
rect 200 141448 800 141568
rect 299200 139408 299800 139528
rect 200 138728 800 138848
rect 299200 136008 299800 136128
rect 200 135328 800 135448
rect 299200 133288 299800 133408
rect 200 132608 800 132728
rect 299200 129888 299800 130008
rect 200 129208 800 129328
rect 299200 127168 299800 127288
rect 200 125808 800 125928
rect 299200 123768 299800 123888
rect 200 123088 800 123208
rect 299200 120368 299800 120488
rect 200 119688 800 119808
rect 299200 117648 299800 117768
rect 200 116968 800 117088
rect 299200 114248 299800 114368
rect 200 113568 800 113688
rect 299200 111528 299800 111648
rect 200 110848 800 110968
rect 299200 108128 299800 108248
rect 200 107448 800 107568
rect 299200 105408 299800 105528
rect 200 104728 800 104848
rect 299200 102008 299800 102128
rect 200 101328 800 101448
rect 299200 99288 299800 99408
rect 200 98608 800 98728
rect 299200 95888 299800 96008
rect 200 95208 800 95328
rect 299200 93168 299800 93288
rect 200 92488 800 92608
rect 299200 89768 299800 89888
rect 200 89088 800 89208
rect 299200 87048 299800 87168
rect 200 85688 800 85808
rect 299200 83648 299800 83768
rect 200 82968 800 83088
rect 299200 80928 299800 81048
rect 200 79568 800 79688
rect 299200 77528 299800 77648
rect 200 76848 800 76968
rect 299200 74128 299800 74248
rect 200 73448 800 73568
rect 299200 71408 299800 71528
rect 200 70728 800 70848
rect 299200 68008 299800 68128
rect 200 67328 800 67448
rect 299200 65288 299800 65408
rect 200 64608 800 64728
rect 299200 61888 299800 62008
rect 200 61208 800 61328
rect 299200 59168 299800 59288
rect 200 58488 800 58608
rect 299200 55768 299800 55888
rect 200 55088 800 55208
rect 299200 53048 299800 53168
rect 200 52368 800 52488
rect 299200 49648 299800 49768
rect 200 48968 800 49088
rect 299200 46928 299800 47048
rect 200 46248 800 46368
rect 299200 43528 299800 43648
rect 200 42848 800 42968
rect 299200 40808 299800 40928
rect 200 39448 800 39568
rect 299200 37408 299800 37528
rect 200 36728 800 36848
rect 299200 34008 299800 34128
rect 200 33328 800 33448
rect 299200 31288 299800 31408
rect 200 30608 800 30728
rect 299200 27888 299800 28008
rect 200 27208 800 27328
rect 299200 25168 299800 25288
rect 200 24488 800 24608
rect 299200 21768 299800 21888
rect 200 21088 800 21208
rect 299200 19048 299800 19168
rect 200 18368 800 18488
rect 299200 15648 299800 15768
rect 200 14968 800 15088
rect 299200 12928 299800 13048
rect 200 12248 800 12368
rect 299200 9528 299800 9648
rect 200 8848 800 8968
rect 299200 6808 299800 6928
rect 200 6128 800 6248
rect 299200 3408 299800 3528
rect 200 2728 800 2848
rect 299200 688 299800 808
<< obsm3 >>
rect 880 298448 299200 298621
rect 800 296688 299200 298448
rect 800 296408 299120 296688
rect 800 296008 299200 296408
rect 880 295728 299200 296008
rect 800 293288 299200 295728
rect 800 293008 299120 293288
rect 800 292608 299200 293008
rect 880 292328 299200 292608
rect 800 290568 299200 292328
rect 800 290288 299120 290568
rect 800 289888 299200 290288
rect 880 289608 299200 289888
rect 800 287168 299200 289608
rect 800 286888 299120 287168
rect 800 286488 299200 286888
rect 880 286208 299200 286488
rect 800 284448 299200 286208
rect 800 284168 299120 284448
rect 800 283768 299200 284168
rect 880 283488 299200 283768
rect 800 281048 299200 283488
rect 800 280768 299120 281048
rect 800 280368 299200 280768
rect 880 280088 299200 280368
rect 800 278328 299200 280088
rect 800 278048 299120 278328
rect 800 277648 299200 278048
rect 880 277368 299200 277648
rect 800 274928 299200 277368
rect 800 274648 299120 274928
rect 800 274248 299200 274648
rect 880 273968 299200 274248
rect 800 272208 299200 273968
rect 800 271928 299120 272208
rect 800 271528 299200 271928
rect 880 271248 299200 271528
rect 800 268808 299200 271248
rect 800 268528 299120 268808
rect 800 268128 299200 268528
rect 880 267848 299200 268128
rect 800 266088 299200 267848
rect 800 265808 299120 266088
rect 800 265408 299200 265808
rect 880 265128 299200 265408
rect 800 262688 299200 265128
rect 800 262408 299120 262688
rect 800 262008 299200 262408
rect 880 261728 299200 262008
rect 800 259968 299200 261728
rect 800 259688 299120 259968
rect 800 258608 299200 259688
rect 880 258328 299200 258608
rect 800 256568 299200 258328
rect 800 256288 299120 256568
rect 800 255888 299200 256288
rect 880 255608 299200 255888
rect 800 253168 299200 255608
rect 800 252888 299120 253168
rect 800 252488 299200 252888
rect 880 252208 299200 252488
rect 800 250448 299200 252208
rect 800 250168 299120 250448
rect 800 249768 299200 250168
rect 880 249488 299200 249768
rect 800 247048 299200 249488
rect 800 246768 299120 247048
rect 800 246368 299200 246768
rect 880 246088 299200 246368
rect 800 244328 299200 246088
rect 800 244048 299120 244328
rect 800 243648 299200 244048
rect 880 243368 299200 243648
rect 800 240928 299200 243368
rect 800 240648 299120 240928
rect 800 240248 299200 240648
rect 880 239968 299200 240248
rect 800 238208 299200 239968
rect 800 237928 299120 238208
rect 800 237528 299200 237928
rect 880 237248 299200 237528
rect 800 234808 299200 237248
rect 800 234528 299120 234808
rect 800 234128 299200 234528
rect 880 233848 299200 234128
rect 800 232088 299200 233848
rect 800 231808 299120 232088
rect 800 231408 299200 231808
rect 880 231128 299200 231408
rect 800 228688 299200 231128
rect 800 228408 299120 228688
rect 800 228008 299200 228408
rect 880 227728 299200 228008
rect 800 225968 299200 227728
rect 800 225688 299120 225968
rect 800 225288 299200 225688
rect 880 225008 299200 225288
rect 800 222568 299200 225008
rect 800 222288 299120 222568
rect 800 221888 299200 222288
rect 880 221608 299200 221888
rect 800 219848 299200 221608
rect 800 219568 299120 219848
rect 800 218488 299200 219568
rect 880 218208 299200 218488
rect 800 216448 299200 218208
rect 800 216168 299120 216448
rect 800 215768 299200 216168
rect 880 215488 299200 215768
rect 800 213728 299200 215488
rect 800 213448 299120 213728
rect 800 212368 299200 213448
rect 880 212088 299200 212368
rect 800 210328 299200 212088
rect 800 210048 299120 210328
rect 800 209648 299200 210048
rect 880 209368 299200 209648
rect 800 206928 299200 209368
rect 800 206648 299120 206928
rect 800 206248 299200 206648
rect 880 205968 299200 206248
rect 800 204208 299200 205968
rect 800 203928 299120 204208
rect 800 203528 299200 203928
rect 880 203248 299200 203528
rect 800 200808 299200 203248
rect 800 200528 299120 200808
rect 800 200128 299200 200528
rect 880 199848 299200 200128
rect 800 198088 299200 199848
rect 800 197808 299120 198088
rect 800 197408 299200 197808
rect 880 197128 299200 197408
rect 800 194688 299200 197128
rect 800 194408 299120 194688
rect 800 194008 299200 194408
rect 880 193728 299200 194008
rect 800 191968 299200 193728
rect 800 191688 299120 191968
rect 800 191288 299200 191688
rect 880 191008 299200 191288
rect 800 188568 299200 191008
rect 800 188288 299120 188568
rect 800 187888 299200 188288
rect 880 187608 299200 187888
rect 800 185848 299200 187608
rect 800 185568 299120 185848
rect 800 185168 299200 185568
rect 880 184888 299200 185168
rect 800 182448 299200 184888
rect 800 182168 299120 182448
rect 800 181768 299200 182168
rect 880 181488 299200 181768
rect 800 179728 299200 181488
rect 800 179448 299120 179728
rect 800 179048 299200 179448
rect 880 178768 299200 179048
rect 800 176328 299200 178768
rect 800 176048 299120 176328
rect 800 175648 299200 176048
rect 880 175368 299200 175648
rect 800 173608 299200 175368
rect 800 173328 299120 173608
rect 800 172248 299200 173328
rect 880 171968 299200 172248
rect 800 170208 299200 171968
rect 800 169928 299120 170208
rect 800 169528 299200 169928
rect 880 169248 299200 169528
rect 800 166808 299200 169248
rect 800 166528 299120 166808
rect 800 166128 299200 166528
rect 880 165848 299200 166128
rect 800 164088 299200 165848
rect 800 163808 299120 164088
rect 800 163408 299200 163808
rect 880 163128 299200 163408
rect 800 160688 299200 163128
rect 800 160408 299120 160688
rect 800 160008 299200 160408
rect 880 159728 299200 160008
rect 800 157968 299200 159728
rect 800 157688 299120 157968
rect 800 157288 299200 157688
rect 880 157008 299200 157288
rect 800 154568 299200 157008
rect 800 154288 299120 154568
rect 800 153888 299200 154288
rect 880 153608 299200 153888
rect 800 151848 299200 153608
rect 800 151568 299120 151848
rect 800 151168 299200 151568
rect 880 150888 299200 151168
rect 800 148448 299200 150888
rect 800 148168 299120 148448
rect 800 147768 299200 148168
rect 880 147488 299200 147768
rect 800 145728 299200 147488
rect 800 145448 299120 145728
rect 800 145048 299200 145448
rect 880 144768 299200 145048
rect 800 142328 299200 144768
rect 800 142048 299120 142328
rect 800 141648 299200 142048
rect 880 141368 299200 141648
rect 800 139608 299200 141368
rect 800 139328 299120 139608
rect 800 138928 299200 139328
rect 880 138648 299200 138928
rect 800 136208 299200 138648
rect 800 135928 299120 136208
rect 800 135528 299200 135928
rect 880 135248 299200 135528
rect 800 133488 299200 135248
rect 800 133208 299120 133488
rect 800 132808 299200 133208
rect 880 132528 299200 132808
rect 800 130088 299200 132528
rect 800 129808 299120 130088
rect 800 129408 299200 129808
rect 880 129128 299200 129408
rect 800 127368 299200 129128
rect 800 127088 299120 127368
rect 800 126008 299200 127088
rect 880 125728 299200 126008
rect 800 123968 299200 125728
rect 800 123688 299120 123968
rect 800 123288 299200 123688
rect 880 123008 299200 123288
rect 800 120568 299200 123008
rect 800 120288 299120 120568
rect 800 119888 299200 120288
rect 880 119608 299200 119888
rect 800 117848 299200 119608
rect 800 117568 299120 117848
rect 800 117168 299200 117568
rect 880 116888 299200 117168
rect 800 114448 299200 116888
rect 800 114168 299120 114448
rect 800 113768 299200 114168
rect 880 113488 299200 113768
rect 800 111728 299200 113488
rect 800 111448 299120 111728
rect 800 111048 299200 111448
rect 880 110768 299200 111048
rect 800 108328 299200 110768
rect 800 108048 299120 108328
rect 800 107648 299200 108048
rect 880 107368 299200 107648
rect 800 105608 299200 107368
rect 800 105328 299120 105608
rect 800 104928 299200 105328
rect 880 104648 299200 104928
rect 800 102208 299200 104648
rect 800 101928 299120 102208
rect 800 101528 299200 101928
rect 880 101248 299200 101528
rect 800 99488 299200 101248
rect 800 99208 299120 99488
rect 800 98808 299200 99208
rect 880 98528 299200 98808
rect 800 96088 299200 98528
rect 800 95808 299120 96088
rect 800 95408 299200 95808
rect 880 95128 299200 95408
rect 800 93368 299200 95128
rect 800 93088 299120 93368
rect 800 92688 299200 93088
rect 880 92408 299200 92688
rect 800 89968 299200 92408
rect 800 89688 299120 89968
rect 800 89288 299200 89688
rect 880 89008 299200 89288
rect 800 87248 299200 89008
rect 800 86968 299120 87248
rect 800 85888 299200 86968
rect 880 85608 299200 85888
rect 800 83848 299200 85608
rect 800 83568 299120 83848
rect 800 83168 299200 83568
rect 880 82888 299200 83168
rect 800 81128 299200 82888
rect 800 80848 299120 81128
rect 800 79768 299200 80848
rect 880 79488 299200 79768
rect 800 77728 299200 79488
rect 800 77448 299120 77728
rect 800 77048 299200 77448
rect 880 76768 299200 77048
rect 800 74328 299200 76768
rect 800 74048 299120 74328
rect 800 73648 299200 74048
rect 880 73368 299200 73648
rect 800 71608 299200 73368
rect 800 71328 299120 71608
rect 800 70928 299200 71328
rect 880 70648 299200 70928
rect 800 68208 299200 70648
rect 800 67928 299120 68208
rect 800 67528 299200 67928
rect 880 67248 299200 67528
rect 800 65488 299200 67248
rect 800 65208 299120 65488
rect 800 64808 299200 65208
rect 880 64528 299200 64808
rect 800 62088 299200 64528
rect 800 61808 299120 62088
rect 800 61408 299200 61808
rect 880 61128 299200 61408
rect 800 59368 299200 61128
rect 800 59088 299120 59368
rect 800 58688 299200 59088
rect 880 58408 299200 58688
rect 800 55968 299200 58408
rect 800 55688 299120 55968
rect 800 55288 299200 55688
rect 880 55008 299200 55288
rect 800 53248 299200 55008
rect 800 52968 299120 53248
rect 800 52568 299200 52968
rect 880 52288 299200 52568
rect 800 49848 299200 52288
rect 800 49568 299120 49848
rect 800 49168 299200 49568
rect 880 48888 299200 49168
rect 800 47128 299200 48888
rect 800 46848 299120 47128
rect 800 46448 299200 46848
rect 880 46168 299200 46448
rect 800 43728 299200 46168
rect 800 43448 299120 43728
rect 800 43048 299200 43448
rect 880 42768 299200 43048
rect 800 41008 299200 42768
rect 800 40728 299120 41008
rect 800 39648 299200 40728
rect 880 39368 299200 39648
rect 800 37608 299200 39368
rect 800 37328 299120 37608
rect 800 36928 299200 37328
rect 880 36648 299200 36928
rect 800 34208 299200 36648
rect 800 33928 299120 34208
rect 800 33528 299200 33928
rect 880 33248 299200 33528
rect 800 31488 299200 33248
rect 800 31208 299120 31488
rect 800 30808 299200 31208
rect 880 30528 299200 30808
rect 800 28088 299200 30528
rect 800 27808 299120 28088
rect 800 27408 299200 27808
rect 880 27128 299200 27408
rect 800 25368 299200 27128
rect 800 25088 299120 25368
rect 800 24688 299200 25088
rect 880 24408 299200 24688
rect 800 21968 299200 24408
rect 800 21688 299120 21968
rect 800 21288 299200 21688
rect 880 21008 299200 21288
rect 800 19248 299200 21008
rect 800 18968 299120 19248
rect 800 18568 299200 18968
rect 880 18288 299200 18568
rect 800 15848 299200 18288
rect 800 15568 299120 15848
rect 800 15168 299200 15568
rect 880 14888 299200 15168
rect 800 13128 299200 14888
rect 800 12848 299120 13128
rect 800 12448 299200 12848
rect 880 12168 299200 12448
rect 800 9728 299200 12168
rect 800 9448 299120 9728
rect 800 9048 299200 9448
rect 880 8768 299200 9048
rect 800 7008 299200 8768
rect 800 6728 299120 7008
rect 800 6328 299200 6728
rect 880 6048 299200 6328
rect 800 3608 299200 6048
rect 800 3328 299120 3608
rect 800 2928 299200 3328
rect 880 2648 299200 2928
rect 800 888 299200 2648
rect 800 715 299120 888
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 28211 297696 288453 298077
rect 28211 2048 34848 297696
rect 35328 2048 50208 297696
rect 50688 2048 65568 297696
rect 66048 2048 80928 297696
rect 81408 2048 96288 297696
rect 96768 2048 111648 297696
rect 112128 2048 127008 297696
rect 127488 2048 142368 297696
rect 142848 2048 157728 297696
rect 158208 2048 173088 297696
rect 173568 2048 188448 297696
rect 188928 2048 203808 297696
rect 204288 2048 219168 297696
rect 219648 2048 234528 297696
rect 235008 2048 249888 297696
rect 250368 2048 265248 297696
rect 265728 2048 280608 297696
rect 281088 2048 288453 297696
rect 28211 1395 288453 2048
<< labels >>
rlabel metal3 s 299200 49648 299800 49768 6 ALU_Output[0]
port 1 nsew signal output
rlabel metal3 s 299200 278128 299800 278248 6 ALU_Output[100]
port 2 nsew signal output
rlabel metal2 s 101770 200 101826 800 6 ALU_Output[101]
port 3 nsew signal output
rlabel metal2 s 165526 299200 165582 299800 6 ALU_Output[102]
port 4 nsew signal output
rlabel metal2 s 31574 200 31630 800 6 ALU_Output[103]
port 5 nsew signal output
rlabel metal3 s 200 181568 800 181688 6 ALU_Output[104]
port 6 nsew signal output
rlabel metal2 s 110142 299200 110198 299800 6 ALU_Output[105]
port 7 nsew signal output
rlabel metal3 s 299200 108128 299800 108248 6 ALU_Output[106]
port 8 nsew signal output
rlabel metal2 s 206742 200 206798 800 6 ALU_Output[107]
port 9 nsew signal output
rlabel metal3 s 200 159808 800 159928 6 ALU_Output[108]
port 10 nsew signal output
rlabel metal2 s 121734 299200 121790 299800 6 ALU_Output[109]
port 11 nsew signal output
rlabel metal3 s 200 21088 800 21208 6 ALU_Output[10]
port 12 nsew signal output
rlabel metal3 s 200 295808 800 295928 6 ALU_Output[110]
port 13 nsew signal output
rlabel metal2 s 182914 299200 182970 299800 6 ALU_Output[111]
port 14 nsew signal output
rlabel metal2 s 213182 200 213238 800 6 ALU_Output[112]
port 15 nsew signal output
rlabel metal2 s 45742 299200 45798 299800 6 ALU_Output[113]
port 16 nsew signal output
rlabel metal2 s 7746 299200 7802 299800 6 ALU_Output[114]
port 17 nsew signal output
rlabel metal3 s 299200 27888 299800 28008 6 ALU_Output[115]
port 18 nsew signal output
rlabel metal3 s 200 18368 800 18488 6 ALU_Output[116]
port 19 nsew signal output
rlabel metal3 s 299200 182248 299800 182368 6 ALU_Output[117]
port 20 nsew signal output
rlabel metal3 s 200 147568 800 147688 6 ALU_Output[118]
port 21 nsew signal output
rlabel metal3 s 299200 290368 299800 290488 6 ALU_Output[119]
port 22 nsew signal output
rlabel metal3 s 200 36728 800 36848 6 ALU_Output[11]
port 23 nsew signal output
rlabel metal2 s 69570 200 69626 800 6 ALU_Output[120]
port 24 nsew signal output
rlabel metal3 s 200 119688 800 119808 6 ALU_Output[121]
port 25 nsew signal output
rlabel metal3 s 299200 240728 299800 240848 6 ALU_Output[122]
port 26 nsew signal output
rlabel metal3 s 299200 268608 299800 268728 6 ALU_Output[123]
port 27 nsew signal output
rlabel metal3 s 200 165928 800 166048 6 ALU_Output[124]
port 28 nsew signal output
rlabel metal2 s 194506 299200 194562 299800 6 ALU_Output[125]
port 29 nsew signal output
rlabel metal3 s 200 33328 800 33448 6 ALU_Output[126]
port 30 nsew signal output
rlabel metal3 s 200 292408 800 292528 6 ALU_Output[127]
port 31 nsew signal output
rlabel metal3 s 299200 200608 299800 200728 6 ALU_Output[12]
port 32 nsew signal output
rlabel metal3 s 200 289688 800 289808 6 ALU_Output[13]
port 33 nsew signal output
rlabel metal2 s 215114 299200 215170 299800 6 ALU_Output[14]
port 34 nsew signal output
rlabel metal2 s 30930 299200 30986 299800 6 ALU_Output[15]
port 35 nsew signal output
rlabel metal3 s 200 123088 800 123208 6 ALU_Output[16]
port 36 nsew signal output
rlabel metal2 s 206098 299200 206154 299800 6 ALU_Output[17]
port 37 nsew signal output
rlabel metal2 s 63130 299200 63186 299800 6 ALU_Output[18]
port 38 nsew signal output
rlabel metal3 s 299200 163888 299800 164008 6 ALU_Output[19]
port 39 nsew signal output
rlabel metal2 s 276938 200 276994 800 6 ALU_Output[1]
port 40 nsew signal output
rlabel metal2 s 78586 200 78642 800 6 ALU_Output[20]
port 41 nsew signal output
rlabel metal2 s 273718 299200 273774 299800 6 ALU_Output[21]
port 42 nsew signal output
rlabel metal3 s 299200 284248 299800 284368 6 ALU_Output[22]
port 43 nsew signal output
rlabel metal2 s 268566 200 268622 800 6 ALU_Output[23]
port 44 nsew signal output
rlabel metal3 s 299200 145528 299800 145648 6 ALU_Output[24]
port 45 nsew signal output
rlabel metal2 s 49606 200 49662 800 6 ALU_Output[25]
port 46 nsew signal output
rlabel metal3 s 299200 129888 299800 130008 6 ALU_Output[26]
port 47 nsew signal output
rlabel metal3 s 299200 222368 299800 222488 6 ALU_Output[27]
port 48 nsew signal output
rlabel metal2 s 159730 299200 159786 299800 6 ALU_Output[28]
port 49 nsew signal output
rlabel metal2 s 22558 299200 22614 299800 6 ALU_Output[29]
port 50 nsew signal output
rlabel metal3 s 200 61208 800 61328 6 ALU_Output[2]
port 51 nsew signal output
rlabel metal2 s 95974 200 96030 800 6 ALU_Output[30]
port 52 nsew signal output
rlabel metal3 s 299200 206728 299800 206848 6 ALU_Output[31]
port 53 nsew signal output
rlabel metal3 s 200 163208 800 163328 6 ALU_Output[32]
port 54 nsew signal output
rlabel metal2 s 226706 299200 226762 299800 6 ALU_Output[33]
port 55 nsew signal output
rlabel metal2 s 294970 200 295026 800 6 ALU_Output[34]
port 56 nsew signal output
rlabel metal3 s 200 6128 800 6248 6 ALU_Output[35]
port 57 nsew signal output
rlabel metal3 s 299200 204008 299800 204128 6 ALU_Output[36]
port 58 nsew signal output
rlabel metal3 s 200 274048 800 274168 6 ALU_Output[37]
port 59 nsew signal output
rlabel metal2 s 127530 299200 127586 299800 6 ALU_Output[38]
port 60 nsew signal output
rlabel metal2 s 242162 200 242218 800 6 ALU_Output[39]
port 61 nsew signal output
rlabel metal3 s 200 107448 800 107568 6 ALU_Output[3]
port 62 nsew signal output
rlabel metal2 s 270498 299200 270554 299800 6 ALU_Output[40]
port 63 nsew signal output
rlabel metal3 s 200 110848 800 110968 6 ALU_Output[41]
port 64 nsew signal output
rlabel metal3 s 299200 61888 299800 62008 6 ALU_Output[42]
port 65 nsew signal output
rlabel metal2 s 57334 299200 57390 299800 6 ALU_Output[43]
port 66 nsew signal output
rlabel metal3 s 200 215568 800 215688 6 ALU_Output[44]
port 67 nsew signal output
rlabel metal2 s 293682 299200 293738 299800 6 ALU_Output[45]
port 68 nsew signal output
rlabel metal3 s 200 261808 800 261928 6 ALU_Output[46]
port 69 nsew signal output
rlabel metal3 s 299200 111528 299800 111648 6 ALU_Output[47]
port 70 nsew signal output
rlabel metal3 s 200 209448 800 209568 6 ALU_Output[48]
port 71 nsew signal output
rlabel metal3 s 299200 296488 299800 296608 6 ALU_Output[49]
port 72 nsew signal output
rlabel metal3 s 299200 262488 299800 262608 6 ALU_Output[4]
port 73 nsew signal output
rlabel metal3 s 200 249568 800 249688 6 ALU_Output[50]
port 74 nsew signal output
rlabel metal3 s 200 218288 800 218408 6 ALU_Output[51]
port 75 nsew signal output
rlabel metal2 s 139766 200 139822 800 6 ALU_Output[52]
port 76 nsew signal output
rlabel metal2 s 16762 299200 16818 299800 6 ALU_Output[53]
port 77 nsew signal output
rlabel metal3 s 299200 225768 299800 225888 6 ALU_Output[54]
port 78 nsew signal output
rlabel metal2 s 253110 299200 253166 299800 6 ALU_Output[55]
port 79 nsew signal output
rlabel metal3 s 299200 210128 299800 210248 6 ALU_Output[56]
port 80 nsew signal output
rlabel metal2 s 247958 200 248014 800 6 ALU_Output[57]
port 81 nsew signal output
rlabel metal3 s 200 157088 800 157208 6 ALU_Output[58]
port 82 nsew signal output
rlabel metal2 s 57978 200 58034 800 6 ALU_Output[59]
port 83 nsew signal output
rlabel metal2 s 177118 299200 177174 299800 6 ALU_Output[5]
port 84 nsew signal output
rlabel metal3 s 200 101328 800 101448 6 ALU_Output[60]
port 85 nsew signal output
rlabel metal3 s 299200 12928 299800 13048 6 ALU_Output[61]
port 86 nsew signal output
rlabel metal3 s 200 76848 800 76968 6 ALU_Output[62]
port 87 nsew signal output
rlabel metal2 s 171966 200 172022 800 6 ALU_Output[63]
port 88 nsew signal output
rlabel metal3 s 200 178848 800 178968 6 ALU_Output[64]
port 89 nsew signal output
rlabel metal2 s 296902 299200 296958 299800 6 ALU_Output[65]
port 90 nsew signal output
rlabel metal3 s 299200 102008 299800 102128 6 ALU_Output[66]
port 91 nsew signal output
rlabel metal3 s 200 225088 800 225208 6 ALU_Output[67]
port 92 nsew signal output
rlabel metal2 s 80518 299200 80574 299800 6 ALU_Output[68]
port 93 nsew signal output
rlabel metal2 s 133970 200 134026 800 6 ALU_Output[69]
port 94 nsew signal output
rlabel metal3 s 299200 87048 299800 87168 6 ALU_Output[6]
port 95 nsew signal output
rlabel metal2 s 37370 200 37426 800 6 ALU_Output[70]
port 96 nsew signal output
rlabel metal3 s 299200 74128 299800 74248 6 ALU_Output[71]
port 97 nsew signal output
rlabel metal3 s 299200 120368 299800 120488 6 ALU_Output[72]
port 98 nsew signal output
rlabel metal2 s 180982 200 181038 800 6 ALU_Output[73]
port 99 nsew signal output
rlabel metal2 s 262770 200 262826 800 6 ALU_Output[74]
port 100 nsew signal output
rlabel metal3 s 299200 31288 299800 31408 6 ALU_Output[75]
port 101 nsew signal output
rlabel metal3 s 200 48968 800 49088 6 ALU_Output[76]
port 102 nsew signal output
rlabel metal2 s 142342 299200 142398 299800 6 ALU_Output[77]
port 103 nsew signal output
rlabel metal2 s 188710 299200 188766 299800 6 ALU_Output[78]
port 104 nsew signal output
rlabel metal3 s 200 206048 800 206168 6 ALU_Output[79]
port 105 nsew signal output
rlabel metal2 s 154578 200 154634 800 6 ALU_Output[7]
port 106 nsew signal output
rlabel metal3 s 200 237328 800 237448 6 ALU_Output[80]
port 107 nsew signal output
rlabel metal2 s 189354 200 189410 800 6 ALU_Output[81]
port 108 nsew signal output
rlabel metal3 s 299200 43528 299800 43648 6 ALU_Output[82]
port 109 nsew signal output
rlabel metal2 s 118514 299200 118570 299800 6 ALU_Output[83]
port 110 nsew signal output
rlabel metal2 s 124310 299200 124366 299800 6 ALU_Output[84]
port 111 nsew signal output
rlabel metal3 s 200 231208 800 231328 6 ALU_Output[85]
port 112 nsew signal output
rlabel metal3 s 299200 197888 299800 198008 6 ALU_Output[86]
port 113 nsew signal output
rlabel metal3 s 200 197208 800 197328 6 ALU_Output[87]
port 114 nsew signal output
rlabel metal2 s 25134 299200 25190 299800 6 ALU_Output[88]
port 115 nsew signal output
rlabel metal3 s 200 193808 800 193928 6 ALU_Output[89]
port 116 nsew signal output
rlabel metal2 s 236366 200 236422 800 6 ALU_Output[8]
port 117 nsew signal output
rlabel metal3 s 200 172048 800 172168 6 ALU_Output[90]
port 118 nsew signal output
rlabel metal2 s 84382 200 84438 800 6 ALU_Output[91]
port 119 nsew signal output
rlabel metal3 s 299200 37408 299800 37528 6 ALU_Output[92]
port 120 nsew signal output
rlabel metal3 s 299200 105408 299800 105528 6 ALU_Output[93]
port 121 nsew signal output
rlabel metal3 s 299200 46928 299800 47048 6 ALU_Output[94]
port 122 nsew signal output
rlabel metal3 s 200 64608 800 64728 6 ALU_Output[95]
port 123 nsew signal output
rlabel metal2 s 19338 299200 19394 299800 6 ALU_Output[96]
port 124 nsew signal output
rlabel metal2 s 247314 299200 247370 299800 6 ALU_Output[97]
port 125 nsew signal output
rlabel metal3 s 200 280168 800 280288 6 ALU_Output[98]
port 126 nsew signal output
rlabel metal2 s 204166 200 204222 800 6 ALU_Output[99]
port 127 nsew signal output
rlabel metal2 s 192574 200 192630 800 6 ALU_Output[9]
port 128 nsew signal output
rlabel metal3 s 200 141448 800 141568 6 Exception[0]
port 129 nsew signal output
rlabel metal3 s 299200 246848 299800 246968 6 Exception[1]
port 130 nsew signal output
rlabel metal2 s 287886 299200 287942 299800 6 Exception[2]
port 131 nsew signal output
rlabel metal2 s 232502 299200 232558 299800 6 Exception[3]
port 132 nsew signal output
rlabel metal2 s 93398 200 93454 800 6 Operation[0]
port 133 nsew signal input
rlabel metal2 s 131394 200 131450 800 6 Operation[1]
port 134 nsew signal input
rlabel metal3 s 200 92488 800 92608 6 Operation[2]
port 135 nsew signal input
rlabel metal3 s 299200 154368 299800 154488 6 Operation[3]
port 136 nsew signal input
rlabel metal2 s 42522 299200 42578 299800 6 Overflow[0]
port 137 nsew signal output
rlabel metal3 s 299200 191768 299800 191888 6 Overflow[1]
port 138 nsew signal output
rlabel metal3 s 200 95208 800 95328 6 Overflow[2]
port 139 nsew signal output
rlabel metal2 s 169390 200 169446 800 6 Overflow[3]
port 140 nsew signal output
rlabel metal2 s 136546 299200 136602 299800 6 Underflow[0]
port 141 nsew signal output
rlabel metal2 s 209318 299200 209374 299800 6 Underflow[1]
port 142 nsew signal output
rlabel metal2 s 66994 200 67050 800 6 Underflow[2]
port 143 nsew signal output
rlabel metal2 s 139122 299200 139178 299800 6 Underflow[3]
port 144 nsew signal output
rlabel metal2 s 128174 200 128230 800 6 a_operand[0]
port 145 nsew signal input
rlabel metal2 s 235722 299200 235778 299800 6 a_operand[100]
port 146 nsew signal input
rlabel metal2 s 156510 299200 156566 299800 6 a_operand[101]
port 147 nsew signal input
rlabel metal3 s 299200 55768 299800 55888 6 a_operand[102]
port 148 nsew signal input
rlabel metal3 s 200 85688 800 85808 6 a_operand[103]
port 149 nsew signal input
rlabel metal2 s 186778 200 186834 800 6 a_operand[104]
port 150 nsew signal input
rlabel metal2 s 86314 299200 86370 299800 6 a_operand[105]
port 151 nsew signal input
rlabel metal2 s 99194 200 99250 800 6 a_operand[106]
port 152 nsew signal input
rlabel metal2 s 119158 200 119214 800 6 a_operand[107]
port 153 nsew signal input
rlabel metal3 s 200 135328 800 135448 6 a_operand[108]
port 154 nsew signal input
rlabel metal3 s 299200 216248 299800 216368 6 a_operand[109]
port 155 nsew signal input
rlabel metal3 s 200 132608 800 132728 6 a_operand[10]
port 156 nsew signal input
rlabel metal2 s 4526 299200 4582 299800 6 a_operand[110]
port 157 nsew signal input
rlabel metal3 s 200 243448 800 243568 6 a_operand[111]
port 158 nsew signal input
rlabel metal2 s 60554 299200 60610 299800 6 a_operand[112]
port 159 nsew signal input
rlabel metal3 s 200 144848 800 144968 6 a_operand[113]
port 160 nsew signal input
rlabel metal3 s 299200 234608 299800 234728 6 a_operand[114]
port 161 nsew signal input
rlabel metal2 s 173898 299200 173954 299800 6 a_operand[115]
port 162 nsew signal input
rlabel metal3 s 200 129208 800 129328 6 a_operand[116]
port 163 nsew signal input
rlabel metal2 s 98550 299200 98606 299800 6 a_operand[117]
port 164 nsew signal input
rlabel metal2 s 198370 200 198426 800 6 a_operand[118]
port 165 nsew signal input
rlabel metal2 s 87602 200 87658 800 6 a_operand[119]
port 166 nsew signal input
rlabel metal2 s 104990 200 105046 800 6 a_operand[11]
port 167 nsew signal input
rlabel metal3 s 299200 99288 299800 99408 6 a_operand[120]
port 168 nsew signal input
rlabel metal3 s 299200 259768 299800 259888 6 a_operand[121]
port 169 nsew signal input
rlabel metal2 s 66350 299200 66406 299800 6 a_operand[122]
port 170 nsew signal input
rlabel metal2 s 168102 299200 168158 299800 6 a_operand[123]
port 171 nsew signal input
rlabel metal3 s 299200 238008 299800 238128 6 a_operand[124]
port 172 nsew signal input
rlabel metal2 s 133326 299200 133382 299800 6 a_operand[125]
port 173 nsew signal input
rlabel metal3 s 299200 252968 299800 253088 6 a_operand[126]
port 174 nsew signal input
rlabel metal3 s 200 252288 800 252408 6 a_operand[127]
port 175 nsew signal input
rlabel metal2 s 10966 299200 11022 299800 6 a_operand[12]
port 176 nsew signal input
rlabel metal2 s 258906 299200 258962 299800 6 a_operand[13]
port 177 nsew signal input
rlabel metal2 s 180338 299200 180394 299800 6 a_operand[14]
port 178 nsew signal input
rlabel metal3 s 299200 65288 299800 65408 6 a_operand[15]
port 179 nsew signal input
rlabel metal2 s 151358 200 151414 800 6 a_operand[16]
port 180 nsew signal input
rlabel metal2 s 186134 299200 186190 299800 6 a_operand[17]
port 181 nsew signal input
rlabel metal3 s 200 283568 800 283688 6 a_operand[18]
port 182 nsew signal input
rlabel metal2 s 1950 299200 2006 299800 6 a_operand[19]
port 183 nsew signal input
rlabel metal2 s 122378 200 122434 800 6 a_operand[1]
port 184 nsew signal input
rlabel metal3 s 200 14968 800 15088 6 a_operand[20]
port 185 nsew signal input
rlabel metal3 s 299200 114248 299800 114368 6 a_operand[21]
port 186 nsew signal input
rlabel metal2 s 291750 200 291806 800 6 a_operand[22]
port 187 nsew signal input
rlabel metal3 s 200 240048 800 240168 6 a_operand[23]
port 188 nsew signal input
rlabel metal3 s 299200 34008 299800 34128 6 a_operand[24]
port 189 nsew signal input
rlabel metal2 s 137190 200 137246 800 6 a_operand[25]
port 190 nsew signal input
rlabel metal3 s 200 212168 800 212288 6 a_operand[26]
port 191 nsew signal input
rlabel metal2 s 34150 299200 34206 299800 6 a_operand[27]
port 192 nsew signal input
rlabel metal2 s 171322 299200 171378 299800 6 a_operand[28]
port 193 nsew signal input
rlabel metal2 s 285954 200 286010 800 6 a_operand[29]
port 194 nsew signal input
rlabel metal3 s 299200 19048 299800 19168 6 a_operand[2]
port 195 nsew signal input
rlabel metal3 s 200 70728 800 70848 6 a_operand[30]
port 196 nsew signal input
rlabel metal2 s 271142 200 271198 800 6 a_operand[31]
port 197 nsew signal input
rlabel metal3 s 200 221688 800 221808 6 a_operand[32]
port 198 nsew signal input
rlabel metal2 s 153934 299200 153990 299800 6 a_operand[33]
port 199 nsew signal input
rlabel metal2 s 17406 200 17462 800 6 a_operand[34]
port 200 nsew signal input
rlabel metal2 s 116582 200 116638 800 6 a_operand[35]
port 201 nsew signal input
rlabel metal3 s 200 199928 800 200048 6 a_operand[36]
port 202 nsew signal input
rlabel metal2 s 259550 200 259606 800 6 a_operand[37]
port 203 nsew signal input
rlabel metal3 s 200 227808 800 227928 6 a_operand[38]
port 204 nsew signal input
rlabel metal3 s 200 24488 800 24608 6 a_operand[39]
port 205 nsew signal input
rlabel metal2 s 256974 200 257030 800 6 a_operand[3]
port 206 nsew signal input
rlabel metal3 s 299200 136008 299800 136128 6 a_operand[40]
port 207 nsew signal input
rlabel metal2 s 68926 299200 68982 299800 6 a_operand[41]
port 208 nsew signal input
rlabel metal3 s 200 116968 800 117088 6 a_operand[42]
port 209 nsew signal input
rlabel metal3 s 299200 688 299800 808 6 a_operand[43]
port 210 nsew signal input
rlabel metal3 s 200 265208 800 265328 6 a_operand[44]
port 211 nsew signal input
rlabel metal2 s 48318 299200 48374 299800 6 a_operand[45]
port 212 nsew signal input
rlabel metal2 s 148138 299200 148194 299800 6 a_operand[46]
port 213 nsew signal input
rlabel metal3 s 299200 53048 299800 53168 6 a_operand[47]
port 214 nsew signal input
rlabel metal2 s 249890 299200 249946 299800 6 a_operand[48]
port 215 nsew signal input
rlabel metal3 s 200 58488 800 58608 6 a_operand[49]
port 216 nsew signal input
rlabel metal3 s 299200 250248 299800 250368 6 a_operand[4]
port 217 nsew signal input
rlabel metal3 s 299200 160488 299800 160608 6 a_operand[50]
port 218 nsew signal input
rlabel metal2 s 264702 299200 264758 299800 6 a_operand[51]
port 219 nsew signal input
rlabel metal2 s 75366 200 75422 800 6 a_operand[52]
port 220 nsew signal input
rlabel metal2 s 244738 200 244794 800 6 a_operand[53]
port 221 nsew signal input
rlabel metal3 s 200 138728 800 138848 6 a_operand[54]
port 222 nsew signal input
rlabel metal3 s 299200 68008 299800 68128 6 a_operand[55]
port 223 nsew signal input
rlabel metal3 s 299200 293088 299800 293208 6 a_operand[56]
port 224 nsew signal input
rlabel metal3 s 200 27208 800 27328 6 a_operand[57]
port 225 nsew signal input
rlabel metal3 s 299200 127168 299800 127288 6 a_operand[58]
port 226 nsew signal input
rlabel metal3 s 299200 95888 299800 96008 6 a_operand[59]
port 227 nsew signal input
rlabel metal3 s 200 298528 800 298648 6 a_operand[5]
port 228 nsew signal input
rlabel metal3 s 299200 151648 299800 151768 6 a_operand[60]
port 229 nsew signal input
rlabel metal2 s 101126 299200 101182 299800 6 a_operand[61]
port 230 nsew signal input
rlabel metal3 s 299200 157768 299800 157888 6 a_operand[62]
port 231 nsew signal input
rlabel metal3 s 200 12248 800 12368 6 a_operand[63]
port 232 nsew signal input
rlabel metal2 s 251178 200 251234 800 6 a_operand[64]
port 233 nsew signal input
rlabel metal2 s 40590 200 40646 800 6 a_operand[65]
port 234 nsew signal input
rlabel metal3 s 200 39448 800 39568 6 a_operand[66]
port 235 nsew signal input
rlabel metal2 s 227350 200 227406 800 6 a_operand[67]
port 236 nsew signal input
rlabel metal3 s 299200 9528 299800 9648 6 a_operand[68]
port 237 nsew signal input
rlabel metal2 s 54758 299200 54814 299800 6 a_operand[69]
port 238 nsew signal input
rlabel metal3 s 200 175448 800 175568 6 a_operand[6]
port 239 nsew signal input
rlabel metal2 s 144918 299200 144974 299800 6 a_operand[70]
port 240 nsew signal input
rlabel metal3 s 200 125808 800 125928 6 a_operand[71]
port 241 nsew signal input
rlabel metal2 s 81162 200 81218 800 6 a_operand[72]
port 242 nsew signal input
rlabel metal3 s 299200 170008 299800 170128 6 a_operand[73]
port 243 nsew signal input
rlabel metal2 s 253754 200 253810 800 6 a_operand[74]
port 244 nsew signal input
rlabel metal2 s 224130 299200 224186 299800 6 a_operand[75]
port 245 nsew signal input
rlabel metal2 s 52182 200 52238 800 6 a_operand[76]
port 246 nsew signal input
rlabel metal2 s 77942 299200 77998 299800 6 a_operand[77]
port 247 nsew signal input
rlabel metal3 s 299200 272008 299800 272128 6 a_operand[78]
port 248 nsew signal input
rlabel metal3 s 299200 286968 299800 287088 6 a_operand[79]
port 249 nsew signal input
rlabel metal3 s 299200 244128 299800 244248 6 a_operand[7]
port 250 nsew signal input
rlabel metal2 s 13542 299200 13598 299800 6 a_operand[80]
port 251 nsew signal input
rlabel metal3 s 299200 231888 299800 232008 6 a_operand[81]
port 252 nsew signal input
rlabel metal2 s 145562 200 145618 800 6 a_operand[82]
port 253 nsew signal input
rlabel metal2 s 279514 299200 279570 299800 6 a_operand[83]
port 254 nsew signal input
rlabel metal2 s 8390 200 8446 800 6 a_operand[84]
port 255 nsew signal input
rlabel metal2 s 2594 200 2650 800 6 a_operand[85]
port 256 nsew signal input
rlabel metal2 s 74722 299200 74778 299800 6 a_operand[86]
port 257 nsew signal input
rlabel metal2 s 148782 200 148838 800 6 a_operand[87]
port 258 nsew signal input
rlabel metal2 s 297546 200 297602 800 6 a_operand[88]
port 259 nsew signal input
rlabel metal2 s 299478 299200 299534 299800 6 a_operand[89]
port 260 nsew signal input
rlabel metal3 s 299200 21768 299800 21888 6 a_operand[8]
port 261 nsew signal input
rlabel metal2 s 130106 299200 130162 299800 6 a_operand[90]
port 262 nsew signal input
rlabel metal3 s 200 46248 800 46368 6 a_operand[91]
port 263 nsew signal input
rlabel metal2 s 55402 200 55458 800 6 a_operand[92]
port 264 nsew signal input
rlabel metal2 s 125598 200 125654 800 6 a_operand[93]
port 265 nsew signal input
rlabel metal2 s 262126 299200 262182 299800 6 a_operand[94]
port 266 nsew signal input
rlabel metal3 s 200 82968 800 83088 6 a_operand[95]
port 267 nsew signal input
rlabel metal2 s 107566 200 107622 800 6 a_operand[96]
port 268 nsew signal input
rlabel metal2 s 215758 200 215814 800 6 a_operand[97]
port 269 nsew signal input
rlabel metal3 s 299200 133288 299800 133408 6 a_operand[98]
port 270 nsew signal input
rlabel metal3 s 299200 188368 299800 188488 6 a_operand[99]
port 271 nsew signal input
rlabel metal2 s 221554 200 221610 800 6 a_operand[9]
port 272 nsew signal input
rlabel metal3 s 200 184968 800 185088 6 b_operand[0]
port 273 nsew signal input
rlabel metal2 s 282734 200 282790 800 6 b_operand[100]
port 274 nsew signal input
rlabel metal3 s 299200 179528 299800 179648 6 b_operand[101]
port 275 nsew signal input
rlabel metal2 s 218334 299200 218390 299800 6 b_operand[102]
port 276 nsew signal input
rlabel metal3 s 200 2728 800 2848 6 b_operand[103]
port 277 nsew signal input
rlabel metal3 s 200 233928 800 234048 6 b_operand[104]
port 278 nsew signal input
rlabel metal2 s 276294 299200 276350 299800 6 b_operand[105]
port 279 nsew signal input
rlabel metal3 s 299200 15648 299800 15768 6 b_operand[106]
port 280 nsew signal input
rlabel metal2 s 191930 299200 191986 299800 6 b_operand[107]
port 281 nsew signal input
rlabel metal2 s 265346 200 265402 800 6 b_operand[108]
port 282 nsew signal input
rlabel metal3 s 200 73448 800 73568 6 b_operand[109]
port 283 nsew signal input
rlabel metal2 s 34794 200 34850 800 6 b_operand[10]
port 284 nsew signal input
rlabel metal3 s 299200 139408 299800 139528 6 b_operand[110]
port 285 nsew signal input
rlabel metal3 s 200 277448 800 277568 6 b_operand[111]
port 286 nsew signal input
rlabel metal3 s 299200 185648 299800 185768 6 b_operand[112]
port 287 nsew signal input
rlabel metal2 s 72790 200 72846 800 6 b_operand[113]
port 288 nsew signal input
rlabel metal2 s 274362 200 274418 800 6 b_operand[114]
port 289 nsew signal input
rlabel metal2 s 104346 299200 104402 299800 6 b_operand[115]
port 290 nsew signal input
rlabel metal2 s 267922 299200 267978 299800 6 b_operand[116]
port 291 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 b_operand[117]
port 292 nsew signal input
rlabel metal2 s 92754 299200 92810 299800 6 b_operand[118]
port 293 nsew signal input
rlabel metal2 s 115938 299200 115994 299800 6 b_operand[119]
port 294 nsew signal input
rlabel metal3 s 299200 40808 299800 40928 6 b_operand[11]
port 295 nsew signal input
rlabel metal2 s 72146 299200 72202 299800 6 b_operand[120]
port 296 nsew signal input
rlabel metal3 s 299200 93168 299800 93288 6 b_operand[121]
port 297 nsew signal input
rlabel metal3 s 200 191088 800 191208 6 b_operand[122]
port 298 nsew signal input
rlabel metal2 s 150714 299200 150770 299800 6 b_operand[123]
port 299 nsew signal input
rlabel metal2 s 36726 299200 36782 299800 6 b_operand[124]
port 300 nsew signal input
rlabel metal2 s 25778 200 25834 800 6 b_operand[125]
port 301 nsew signal input
rlabel metal2 s 160374 200 160430 800 6 b_operand[126]
port 302 nsew signal input
rlabel metal3 s 299200 213528 299800 213648 6 b_operand[127]
port 303 nsew signal input
rlabel metal3 s 299200 194488 299800 194608 6 b_operand[12]
port 304 nsew signal input
rlabel metal2 s 183558 200 183614 800 6 b_operand[13]
port 305 nsew signal input
rlabel metal3 s 299200 173408 299800 173528 6 b_operand[14]
port 306 nsew signal input
rlabel metal3 s 299200 83648 299800 83768 6 b_operand[15]
port 307 nsew signal input
rlabel metal2 s 280158 200 280214 800 6 b_operand[16]
port 308 nsew signal input
rlabel metal2 s 203522 299200 203578 299800 6 b_operand[17]
port 309 nsew signal input
rlabel metal2 s 285310 299200 285366 299800 6 b_operand[18]
port 310 nsew signal input
rlabel metal2 s 162950 200 163006 800 6 b_operand[19]
port 311 nsew signal input
rlabel metal2 s 233146 200 233202 800 6 b_operand[1]
port 312 nsew signal input
rlabel metal3 s 299200 59168 299800 59288 6 b_operand[20]
port 313 nsew signal input
rlabel metal2 s 51538 299200 51594 299800 6 b_operand[21]
port 314 nsew signal input
rlabel metal3 s 200 55088 800 55208 6 b_operand[22]
port 315 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 b_operand[23]
port 316 nsew signal input
rlabel metal2 s 112718 299200 112774 299800 6 b_operand[24]
port 317 nsew signal input
rlabel metal3 s 200 113568 800 113688 6 b_operand[25]
port 318 nsew signal input
rlabel metal3 s 299200 280848 299800 280968 6 b_operand[26]
port 319 nsew signal input
rlabel metal2 s 113362 200 113418 800 6 b_operand[27]
port 320 nsew signal input
rlabel metal2 s 244094 299200 244150 299800 6 b_operand[28]
port 321 nsew signal input
rlabel metal3 s 299200 117648 299800 117768 6 b_operand[29]
port 322 nsew signal input
rlabel metal2 s 224774 200 224830 800 6 b_operand[2]
port 323 nsew signal input
rlabel metal2 s 238298 299200 238354 299800 6 b_operand[30]
port 324 nsew signal input
rlabel metal2 s 218978 200 219034 800 6 b_operand[31]
port 325 nsew signal input
rlabel metal3 s 200 153688 800 153808 6 b_operand[32]
port 326 nsew signal input
rlabel metal2 s 14186 200 14242 800 6 b_operand[33]
port 327 nsew signal input
rlabel metal2 s 288530 200 288586 800 6 b_operand[34]
port 328 nsew signal input
rlabel metal3 s 299200 71408 299800 71528 6 b_operand[35]
port 329 nsew signal input
rlabel metal2 s 106922 299200 106978 299800 6 b_operand[36]
port 330 nsew signal input
rlabel metal3 s 299200 256368 299800 256488 6 b_operand[37]
port 331 nsew signal input
rlabel metal3 s 200 246168 800 246288 6 b_operand[38]
port 332 nsew signal input
rlabel metal3 s 200 267928 800 268048 6 b_operand[39]
port 333 nsew signal input
rlabel metal3 s 200 258408 800 258528 6 b_operand[3]
port 334 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 b_operand[40]
port 335 nsew signal input
rlabel metal3 s 200 8848 800 8968 6 b_operand[41]
port 336 nsew signal input
rlabel metal3 s 299200 148248 299800 148368 6 b_operand[42]
port 337 nsew signal input
rlabel metal2 s 166170 200 166226 800 6 b_operand[43]
port 338 nsew signal input
rlabel metal3 s 200 52368 800 52488 6 b_operand[44]
port 339 nsew signal input
rlabel metal2 s 282090 299200 282146 299800 6 b_operand[45]
port 340 nsew signal input
rlabel metal2 s 28354 299200 28410 299800 6 b_operand[46]
port 341 nsew signal input
rlabel metal2 s 43810 200 43866 800 6 b_operand[47]
port 342 nsew signal input
rlabel metal3 s 200 79568 800 79688 6 b_operand[48]
port 343 nsew signal input
rlabel metal2 s 291106 299200 291162 299800 6 b_operand[49]
port 344 nsew signal input
rlabel metal3 s 200 187688 800 187808 6 b_operand[4]
port 345 nsew signal input
rlabel metal3 s 200 42848 800 42968 6 b_operand[50]
port 346 nsew signal input
rlabel metal3 s 299200 89768 299800 89888 6 b_operand[51]
port 347 nsew signal input
rlabel metal2 s 200946 200 201002 800 6 b_operand[52]
port 348 nsew signal input
rlabel metal2 s 255686 299200 255742 299800 6 b_operand[53]
port 349 nsew signal input
rlabel metal2 s 83738 299200 83794 299800 6 b_operand[54]
port 350 nsew signal input
rlabel metal2 s 90178 200 90234 800 6 b_operand[55]
port 351 nsew signal input
rlabel metal3 s 299200 176128 299800 176248 6 b_operand[56]
port 352 nsew signal input
rlabel metal2 s 238942 200 238998 800 6 b_operand[57]
port 353 nsew signal input
rlabel metal3 s 299200 80928 299800 81048 6 b_operand[58]
port 354 nsew signal input
rlabel metal3 s 200 169328 800 169448 6 b_operand[59]
port 355 nsew signal input
rlabel metal3 s 299200 3408 299800 3528 6 b_operand[5]
port 356 nsew signal input
rlabel metal2 s 46386 200 46442 800 6 b_operand[60]
port 357 nsew signal input
rlabel metal2 s 142986 200 143042 800 6 b_operand[61]
port 358 nsew signal input
rlabel metal3 s 299200 123768 299800 123888 6 b_operand[62]
port 359 nsew signal input
rlabel metal2 s 241518 299200 241574 299800 6 b_operand[63]
port 360 nsew signal input
rlabel metal3 s 299200 265888 299800 266008 6 b_operand[64]
port 361 nsew signal input
rlabel metal3 s 299200 6808 299800 6928 6 b_operand[65]
port 362 nsew signal input
rlabel metal2 s 23202 200 23258 800 6 b_operand[66]
port 363 nsew signal input
rlabel metal3 s 299200 166608 299800 166728 6 b_operand[67]
port 364 nsew signal input
rlabel metal2 s 5814 200 5870 800 6 b_operand[68]
port 365 nsew signal input
rlabel metal3 s 299200 274728 299800 274848 6 b_operand[69]
port 366 nsew signal input
rlabel metal2 s 229926 299200 229982 299800 6 b_operand[6]
port 367 nsew signal input
rlabel metal3 s 299200 25168 299800 25288 6 b_operand[70]
port 368 nsew signal input
rlabel metal2 s 220910 299200 220966 299800 6 b_operand[71]
port 369 nsew signal input
rlabel metal3 s 200 89088 800 89208 6 b_operand[72]
port 370 nsew signal input
rlabel metal3 s 200 98608 800 98728 6 b_operand[73]
port 371 nsew signal input
rlabel metal2 s 195150 200 195206 800 6 b_operand[74]
port 372 nsew signal input
rlabel metal2 s 18 200 74 800 6 b_operand[75]
port 373 nsew signal input
rlabel metal2 s 230570 200 230626 800 6 b_operand[76]
port 374 nsew signal input
rlabel metal3 s 200 150968 800 151088 6 b_operand[77]
port 375 nsew signal input
rlabel metal3 s 200 271328 800 271448 6 b_operand[78]
port 376 nsew signal input
rlabel metal2 s 89534 299200 89590 299800 6 b_operand[79]
port 377 nsew signal input
rlabel metal3 s 200 104728 800 104848 6 b_operand[7]
port 378 nsew signal input
rlabel metal2 s 61198 200 61254 800 6 b_operand[80]
port 379 nsew signal input
rlabel metal2 s 19982 200 20038 800 6 b_operand[81]
port 380 nsew signal input
rlabel metal2 s 162306 299200 162362 299800 6 b_operand[82]
port 381 nsew signal input
rlabel metal2 s 95330 299200 95386 299800 6 b_operand[83]
port 382 nsew signal input
rlabel metal2 s 157154 200 157210 800 6 b_operand[84]
port 383 nsew signal input
rlabel metal2 s 211894 299200 211950 299800 6 b_operand[85]
port 384 nsew signal input
rlabel metal3 s 299200 77528 299800 77648 6 b_operand[86]
port 385 nsew signal input
rlabel metal3 s 200 203328 800 203448 6 b_operand[87]
port 386 nsew signal input
rlabel metal3 s 299200 228488 299800 228608 6 b_operand[88]
port 387 nsew signal input
rlabel metal2 s 63774 200 63830 800 6 b_operand[89]
port 388 nsew signal input
rlabel metal2 s 110786 200 110842 800 6 b_operand[8]
port 389 nsew signal input
rlabel metal2 s 175186 200 175242 800 6 b_operand[90]
port 390 nsew signal input
rlabel metal3 s 299200 219648 299800 219768 6 b_operand[91]
port 391 nsew signal input
rlabel metal2 s 177762 200 177818 800 6 b_operand[92]
port 392 nsew signal input
rlabel metal2 s 200302 299200 200358 299800 6 b_operand[93]
port 393 nsew signal input
rlabel metal2 s 197726 299200 197782 299800 6 b_operand[94]
port 394 nsew signal input
rlabel metal3 s 200 286288 800 286408 6 b_operand[95]
port 395 nsew signal input
rlabel metal2 s 39946 299200 40002 299800 6 b_operand[96]
port 396 nsew signal input
rlabel metal2 s 209962 200 210018 800 6 b_operand[97]
port 397 nsew signal input
rlabel metal3 s 200 67328 800 67448 6 b_operand[98]
port 398 nsew signal input
rlabel metal3 s 200 255688 800 255808 6 b_operand[99]
port 399 nsew signal input
rlabel metal3 s 299200 142128 299800 142248 6 b_operand[9]
port 400 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 401 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 402 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 189269652
string GDS_FILE /home/urielcho/Proyectos_caravel/MPW8/gf180_vs_sky130/openlane/ALU/runs/22_12_22_14_19/results/signoff/Top_Module_4_ALU.magic.gds
string GDS_START 1760112
<< end >>

